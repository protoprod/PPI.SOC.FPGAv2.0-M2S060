-- Version: v11.8 11.8.0.26

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreAPB3 is

    port( m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR : in    std_logic_vector(15 downto 12);
          CoreAPB3_0_APBmslave0_PSELx            : out   std_logic;
          m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx : in    std_logic
        );

end CoreAPB3;

architecture DEF_ARCH of CoreAPB3 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \iPSELS_raw_1[0]_net_1\, GND_net_1, VCC_net_1
         : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \iPSELS_raw_1[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(15), B
         => m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(14), Y => 
        \iPSELS_raw_1[0]_net_1\);
    
    \iPSELS_raw[0]\ : CFG4
      generic map(INIT => x"0008")

      port map(A => m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx, B => 
        \iPSELS_raw_1[0]_net_1\, C => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(13), D => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(12), Y => 
        CoreAPB3_0_APBmslave0_PSELx);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_CommsFPGA_CCC_0_FCCC is

    port( m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC : in    std_logic;
          CommsFPGA_CCC_0_LOCK                      : out   std_logic;
          CommsFPGA_CCC_0_GL1                       : out   std_logic;
          CommsFPGA_CCC_0_GL0                       : out   std_logic
        );

end m2s010_som_CommsFPGA_CCC_0_FCCC;

architecture DEF_ARCH of m2s010_som_CommsFPGA_CCC_0_FCCC is 

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CCC

            generic (INIT:std_logic_vector(209 downto 0) := "00" & x"0000000000000000000000000000000000000000000000000000"; 
        VCOFREQUENCY:real := 0.0);

    port( Y0              : out   std_logic;
          Y1              : out   std_logic;
          Y2              : out   std_logic;
          Y3              : out   std_logic;
          PRDATA          : out   std_logic_vector(7 downto 0);
          LOCK            : out   std_logic;
          BUSY            : out   std_logic;
          CLK0            : in    std_logic := 'U';
          CLK1            : in    std_logic := 'U';
          CLK2            : in    std_logic := 'U';
          CLK3            : in    std_logic := 'U';
          NGMUX0_SEL      : in    std_logic := 'U';
          NGMUX1_SEL      : in    std_logic := 'U';
          NGMUX2_SEL      : in    std_logic := 'U';
          NGMUX3_SEL      : in    std_logic := 'U';
          NGMUX0_HOLD_N   : in    std_logic := 'U';
          NGMUX1_HOLD_N   : in    std_logic := 'U';
          NGMUX2_HOLD_N   : in    std_logic := 'U';
          NGMUX3_HOLD_N   : in    std_logic := 'U';
          NGMUX0_ARST_N   : in    std_logic := 'U';
          NGMUX1_ARST_N   : in    std_logic := 'U';
          NGMUX2_ARST_N   : in    std_logic := 'U';
          NGMUX3_ARST_N   : in    std_logic := 'U';
          PLL_BYPASS_N    : in    std_logic := 'U';
          PLL_ARST_N      : in    std_logic := 'U';
          PLL_POWERDOWN_N : in    std_logic := 'U';
          GPD0_ARST_N     : in    std_logic := 'U';
          GPD1_ARST_N     : in    std_logic := 'U';
          GPD2_ARST_N     : in    std_logic := 'U';
          GPD3_ARST_N     : in    std_logic := 'U';
          PRESET_N        : in    std_logic := 'U';
          PCLK            : in    std_logic := 'U';
          PSEL            : in    std_logic := 'U';
          PENABLE         : in    std_logic := 'U';
          PWRITE          : in    std_logic := 'U';
          PADDR           : in    std_logic_vector(7 downto 2) := (others => 'U');
          PWDATA          : in    std_logic_vector(7 downto 0) := (others => 'U');
          CLK0_PAD        : in    std_logic := 'U';
          CLK1_PAD        : in    std_logic := 'U';
          CLK2_PAD        : in    std_logic := 'U';
          CLK3_PAD        : in    std_logic := 'U';
          GL0             : out   std_logic;
          GL1             : out   std_logic;
          GL2             : out   std_logic;
          GL3             : out   std_logic;
          RCOSC_25_50MHZ  : in    std_logic := 'U';
          RCOSC_1MHZ      : in    std_logic := 'U';
          XTLOSC          : in    std_logic := 'U'
        );
  end component;

    signal GL0_net, GL1_net, VCC_net_1, GND_net_1 : std_logic;
    signal nc8, nc7, nc6, nc2, nc5, nc4, nc3, nc1 : std_logic;

begin 


    GL1_INST : CLKINT
      port map(A => GL1_net, Y => CommsFPGA_CCC_0_GL1);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    GL0_INST : CLKINT
      port map(A => GL0_net, Y => CommsFPGA_CCC_0_GL0);
    
    CCC_INST : CCC

              generic map(INIT => "00" & x"000007FB8000044164000F18C6309C231839DE40404C41803000",
         VCOFREQUENCY => 980.0)

      port map(Y0 => OPEN, Y1 => OPEN, Y2 => OPEN, Y3 => OPEN, 
        PRDATA(7) => nc8, PRDATA(6) => nc7, PRDATA(5) => nc6, 
        PRDATA(4) => nc2, PRDATA(3) => nc5, PRDATA(2) => nc4, 
        PRDATA(1) => nc3, PRDATA(0) => nc1, LOCK => 
        CommsFPGA_CCC_0_LOCK, BUSY => OPEN, CLK0 => VCC_net_1, 
        CLK1 => VCC_net_1, CLK2 => VCC_net_1, CLK3 => VCC_net_1, 
        NGMUX0_SEL => GND_net_1, NGMUX1_SEL => GND_net_1, 
        NGMUX2_SEL => GND_net_1, NGMUX3_SEL => GND_net_1, 
        NGMUX0_HOLD_N => VCC_net_1, NGMUX1_HOLD_N => VCC_net_1, 
        NGMUX2_HOLD_N => VCC_net_1, NGMUX3_HOLD_N => VCC_net_1, 
        NGMUX0_ARST_N => VCC_net_1, NGMUX1_ARST_N => VCC_net_1, 
        NGMUX2_ARST_N => VCC_net_1, NGMUX3_ARST_N => VCC_net_1, 
        PLL_BYPASS_N => VCC_net_1, PLL_ARST_N => VCC_net_1, 
        PLL_POWERDOWN_N => VCC_net_1, GPD0_ARST_N => VCC_net_1, 
        GPD1_ARST_N => VCC_net_1, GPD2_ARST_N => VCC_net_1, 
        GPD3_ARST_N => VCC_net_1, PRESET_N => GND_net_1, PCLK => 
        VCC_net_1, PSEL => VCC_net_1, PENABLE => VCC_net_1, 
        PWRITE => VCC_net_1, PADDR(7) => VCC_net_1, PADDR(6) => 
        VCC_net_1, PADDR(5) => VCC_net_1, PADDR(4) => VCC_net_1, 
        PADDR(3) => VCC_net_1, PADDR(2) => VCC_net_1, PWDATA(7)
         => VCC_net_1, PWDATA(6) => VCC_net_1, PWDATA(5) => 
        VCC_net_1, PWDATA(4) => VCC_net_1, PWDATA(3) => VCC_net_1, 
        PWDATA(2) => VCC_net_1, PWDATA(1) => VCC_net_1, PWDATA(0)
         => VCC_net_1, CLK0_PAD => GND_net_1, CLK1_PAD => 
        GND_net_1, CLK2_PAD => GND_net_1, CLK3_PAD => GND_net_1, 
        GL0 => GL0_net, GL1 => GL1_net, GL2 => OPEN, GL3 => OPEN, 
        RCOSC_25_50MHZ => GND_net_1, RCOSC_1MHZ => GND_net_1, 
        XTLOSC => m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_ID_RES_0_IO is

    port( ID_RES  : in    std_logic_vector(3 downto 0);
          Y_net_0 : out   std_logic_vector(3 downto 0)
        );

end m2s010_som_ID_RES_0_IO;

architecture DEF_ARCH of m2s010_som_ID_RES_0_IO is 

  component INBUF
    generic (IOSTD:string := "");

    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    U0_0 : INBUF
      port map(PAD => ID_RES(0), Y => Y_net_0(0));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    U0_3 : INBUF
      port map(PAD => ID_RES(3), Y => Y_net_0(3));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    U0_2 : INBUF
      port map(PAD => ID_RES(2), Y => Y_net_0(2));
    
    U0_1 : INBUF
      port map(PAD => ID_RES(1), Y => Y_net_0(1));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb_GPIO_1_IO is

    port( GPIO_1_BI_0                       : inout std_logic := 'Z';
          GPIO_1_in_0                       : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_1_M2F_OE : in    std_logic;
          GPIO_1_M2F                        : in    std_logic
        );

end m2s010_som_sb_GPIO_1_IO;

architecture DEF_ARCH of m2s010_som_sb_GPIO_1_IO is 

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    U0_0 : BIBUF
      generic map(IOSTD => "LVCMOS33")

      port map(PAD => GPIO_1_BI_0, D => GPIO_1_M2F, E => 
        m2s010_som_sb_MSS_0_GPIO_1_M2F_OE, Y => GPIO_1_in_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb_CAM_SPI_1_CLK_IO is

    port( CAM_SPI_1_CLK_Y_0                    : out   std_logic;
          SPI_1_CLK_0                          : inout std_logic := 'Z';
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE : in    std_logic;
          m2s010_som_sb_MSS_0_SPI_1_CLK_M2F    : in    std_logic
        );

end m2s010_som_sb_CAM_SPI_1_CLK_IO;

architecture DEF_ARCH of m2s010_som_sb_CAM_SPI_1_CLK_IO is 

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    U0_0 : BIBUF
      port map(PAD => SPI_1_CLK_0, D => 
        m2s010_som_sb_MSS_0_SPI_1_CLK_M2F, E => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE, Y => 
        CAM_SPI_1_CLK_Y_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb_GPIO_7_IO is

    port( GPIO_7_PADI_0                     : inout std_logic := 'Z';
          GPIO_7_Y_0                        : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_7_M2F_OE : in    std_logic;
          m2s010_som_sb_MSS_0_GPIO_7_M2F    : in    std_logic
        );

end m2s010_som_sb_GPIO_7_IO;

architecture DEF_ARCH of m2s010_som_sb_GPIO_7_IO is 

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    U0_0 : BIBUF
      port map(PAD => GPIO_7_PADI_0, D => 
        m2s010_som_sb_MSS_0_GPIO_7_M2F, E => 
        m2s010_som_sb_MSS_0_GPIO_7_M2F_OE, Y => GPIO_7_Y_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb_CAM_SPI_1_SS0_IO is

    port( SPI_1_SS0_CAM_0                      : inout std_logic := 'Z';
          CAM_SPI_1_SS0_Y_0                    : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE : in    std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F    : in    std_logic
        );

end m2s010_som_sb_CAM_SPI_1_SS0_IO;

architecture DEF_ARCH of m2s010_som_sb_CAM_SPI_1_SS0_IO is 

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    U0_0 : BIBUF
      port map(PAD => SPI_1_SS0_CAM_0, D => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F, E => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE, Y => 
        CAM_SPI_1_SS0_Y_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb_MSS is

    port( CORECONFIGP_0_MDDR_APBmslave_PWDATA              : in    std_logic_vector(15 downto 0);
          CORECONFIGP_0_MDDR_APBmslave_PADDR               : in    std_logic_vector(10 downto 2);
          MAC_MII_RXD_c                                    : in    std_logic_vector(3 downto 0);
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA  : in    std_logic_vector(17 downto 0);
          Y_net_0                                          : in    std_logic_vector(3 downto 0);
          CoreAPB3_0_APBmslave0_PRDATA_m                   : in    std_logic_vector(7 downto 0);
          CORECONFIGP_0_MDDR_APBmslave_PRDATA              : out   std_logic_vector(15 downto 1);
          MAC_MII_TXD_c                                    : out   std_logic_vector(3 downto 0);
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA  : out   std_logic_vector(16 downto 0);
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR   : out   std_logic_vector(15 downto 2);
          CoreAPB3_0_APBmslave0_PWDATA                     : out   std_logic_vector(7 downto 0);
          m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR           : out   std_logic_vector(15 downto 12);
          CoreAPB3_0_APBmslave0_PADDR                      : out   std_logic_vector(7 downto 0);
          MDDR_ADDR                                        : out   std_logic_vector(15 downto 0);
          MDDR_BA                                          : out   std_logic_vector(2 downto 0);
          MDDR_DM_RDQS                                     : inout std_logic_vector(1 downto 0) := (others => 'Z');
          MDDR_DQ                                          : inout std_logic_vector(15 downto 0) := (others => 'Z');
          MDDR_DQS                                         : inout std_logic_vector(1 downto 0) := (others => 'Z');
          CAM_SPI_1_CLK_Y_0                                : in    std_logic;
          GPIO_7_Y_0                                       : in    std_logic;
          GPIO_6_Y_0                                       : in    std_logic;
          DEBOUNCE_OUT_net_0_0                             : in    std_logic;
          GPIO_1_in_0                                      : in    std_logic;
          state_0                                          : in    std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PRDATA_reto_0       : out   std_logic;
          MDDR_CLK                                         : out   std_logic;
          MDDR_CLK_N                                       : out   std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PWRITE              : in    std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PSELx               : in    std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PENABLE             : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz                        : in    std_logic;
          MAC_MII_TX_CLK_c                                 : in    std_logic;
          SPI_1_SS0_MX_Y                                   : in    std_logic;
          SPI_1_DI                                         : in    std_logic;
          MAC_MII_RX_ER_c                                  : in    std_logic;
          MAC_MII_RX_DV_c                                  : in    std_logic;
          MAC_MII_RX_CLK_c                                 : in    std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR : in    std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY  : in    std_logic;
          MMUART_0_RXD_F2M_c                               : in    std_logic;
          DEBOUNCE_OUT_2_c                                 : in    std_logic;
          DEBOUNCE_OUT_1_c                                 : in    std_logic;
          BIBUF_0_Y                                        : in    std_logic;
          FAB_CCC_LOCK                                     : in    std_logic;
          CoreAPB3_0_APBmslave0_PREADY_i_m_i               : in    std_logic;
          CommsFPGA_top_0_INT                              : in    std_logic;
          MAC_MII_CRS_c                                    : in    std_logic;
          MAC_MII_COL_c                                    : in    std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PSLVERR             : out   std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PREADY              : out   std_logic;
          MAC_MII_TX_EN_c                                  : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE             : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F                : out   std_logic;
          SPI_1_DO_CAM_c                                   : out   std_logic;
          GPIO_11_M2F_c                                    : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_CLK_M2F                : out   std_logic;
          GPIO_8_M2F_c                                     : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_7_M2F                   : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_7_M2F_OE                : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_6_M2F                   : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_6_M2F_OE                : out   std_logic;
          GPIO_5_M2F_c                                     : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE  : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx   : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE : out   std_logic;
          GPIO_24_M2F_c                                    : out   std_logic;
          MMUART_0_TXD_M2F_c                               : out   std_logic;
          m2s010_som_sb_0_GPIO_28_SW_RESET                 : out   std_logic;
          GPIO_21_M2F_c                                    : out   std_logic;
          GPIO_22_M2F_c                                    : out   std_logic;
          m2s010_som_sb_MSS_0_MAC_MII_MDO                  : out   std_logic;
          m2s010_som_sb_MSS_0_MAC_MII_MDO_EN               : out   std_logic;
          MAC_MII_MDC_c                                    : out   std_logic;
          GPIO_1_M2F                                       : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_1_M2F_OE                : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F          : out   std_logic;
          CoreAPB3_0_APBmslave0_PWRITE                     : out   std_logic;
          m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx           : out   std_logic;
          CoreAPB3_0_APBmslave0_PENABLE                    : out   std_logic;
          GPIO_0_BI                                        : inout std_logic := 'Z';
          GPIO_3_BI                                        : inout std_logic := 'Z';
          GPIO_4_BI                                        : inout std_logic := 'Z';
          GPIO_12_BI                                       : inout std_logic := 'Z';
          GPIO_14_BI                                       : inout std_logic := 'Z';
          GPIO_15_BI                                       : inout std_logic := 'Z';
          GPIO_16_BI                                       : inout std_logic := 'Z';
          GPIO_17_BI                                       : inout std_logic := 'Z';
          GPIO_18_BI                                       : inout std_logic := 'Z';
          GPIO_20_OUT                                      : out   std_logic;
          GPIO_25_BI                                       : inout std_logic := 'Z';
          GPIO_26_BI                                       : inout std_logic := 'Z';
          GPIO_31_BI                                       : inout std_logic := 'Z';
          I2C_1_SCL                                        : inout std_logic := 'Z';
          I2C_1_SDA                                        : inout std_logic := 'Z';
          MDDR_CAS_N                                       : out   std_logic;
          MDDR_CKE                                         : out   std_logic;
          MDDR_CS_N                                        : out   std_logic;
          MDDR_DQS_TMATCH_0_IN                             : in    std_logic;
          MDDR_DQS_TMATCH_0_OUT                            : out   std_logic;
          MDDR_ODT                                         : out   std_logic;
          MDDR_RAS_N                                       : out   std_logic;
          MDDR_RESET_N                                     : out   std_logic;
          MDDR_WE_N                                        : out   std_logic;
          MMUART_1_RXD                                     : in    std_logic;
          MMUART_1_TXD                                     : out   std_logic;
          SPI_0_CLK                                        : inout std_logic := 'Z';
          SPI_0_DI                                         : in    std_logic;
          SPI_0_DO                                         : out   std_logic;
          SPI_0_SS0                                        : inout std_logic := 'Z';
          SPI_0_SS1                                        : out   std_logic;
          CORECONFIGP_0_APB_S_PCLK_i                       : out   std_logic;
          CORECONFIGP_0_APB_S_PRESET_N                     : out   std_logic;
          CORECONFIGP_0_APB_S_PCLK                         : out   std_logic
        );

end m2s010_som_sb_MSS;

architecture DEF_ARCH of m2s010_som_sb_MSS is 

  component OUTBUF
    generic (IOSTD:string := "");

    port( D   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component TRIBUFF
    generic (IOSTD:string := "");

    port( D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component INBUF
    generic (IOSTD:string := "");

    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component MSS_060

            generic (INIT:std_logic_vector(1437 downto 0) := "00" & x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"; 
        ACT_UBITS:std_logic_vector(55 downto 0) := x"FFFFFFFFFFFFFF"; 
        MEMORYFILE:string := ""; RTC_MAIN_XTL_FREQ:real := 0.0; 
        RTC_MAIN_XTL_MODE:string := "1"; DDR_CLK_FREQ:real := 0.0
        );

    port( CAN_RXBUS_MGPIO3A_H2F_A                 : out   std_logic;
          CAN_RXBUS_MGPIO3A_H2F_B                 : out   std_logic;
          CAN_TX_EBL_MGPIO4A_H2F_A                : out   std_logic;
          CAN_TX_EBL_MGPIO4A_H2F_B                : out   std_logic;
          CAN_TXBUS_MGPIO2A_H2F_A                 : out   std_logic;
          CAN_TXBUS_MGPIO2A_H2F_B                 : out   std_logic;
          CLK_CONFIG_APB                          : out   std_logic;
          COMMS_INT                               : out   std_logic;
          CONFIG_PRESET_N                         : out   std_logic;
          EDAC_ERROR                              : out   std_logic_vector(7 downto 0);
          F_FM0_RDATA                             : out   std_logic_vector(31 downto 0);
          F_FM0_READYOUT                          : out   std_logic;
          F_FM0_RESP                              : out   std_logic;
          F_HM0_ADDR                              : out   std_logic_vector(31 downto 0);
          F_HM0_ENABLE                            : out   std_logic;
          F_HM0_SEL                               : out   std_logic;
          F_HM0_SIZE                              : out   std_logic_vector(1 downto 0);
          F_HM0_TRANS1                            : out   std_logic;
          F_HM0_WDATA                             : out   std_logic_vector(31 downto 0);
          F_HM0_WRITE                             : out   std_logic;
          FAB_CHRGVBUS                            : out   std_logic;
          FAB_DISCHRGVBUS                         : out   std_logic;
          FAB_DMPULLDOWN                          : out   std_logic;
          FAB_DPPULLDOWN                          : out   std_logic;
          FAB_DRVVBUS                             : out   std_logic;
          FAB_IDPULLUP                            : out   std_logic;
          FAB_OPMODE                              : out   std_logic_vector(1 downto 0);
          FAB_SUSPENDM                            : out   std_logic;
          FAB_TERMSEL                             : out   std_logic;
          FAB_TXVALID                             : out   std_logic;
          FAB_VCONTROL                            : out   std_logic_vector(3 downto 0);
          FAB_VCONTROLLOADM                       : out   std_logic;
          FAB_XCVRSEL                             : out   std_logic_vector(1 downto 0);
          FAB_XDATAOUT                            : out   std_logic_vector(7 downto 0);
          FACC_GLMUX_SEL                          : out   std_logic;
          FIC32_0_MASTER                          : out   std_logic_vector(1 downto 0);
          FIC32_1_MASTER                          : out   std_logic_vector(1 downto 0);
          FPGA_RESET_N                            : out   std_logic;
          GTX_CLK                                 : out   std_logic;
          H2F_INTERRUPT                           : out   std_logic_vector(15 downto 0);
          H2F_NMI                                 : out   std_logic;
          H2FCALIB                                : out   std_logic;
          I2C0_SCL_MGPIO31B_H2F_A                 : out   std_logic;
          I2C0_SCL_MGPIO31B_H2F_B                 : out   std_logic;
          I2C0_SDA_MGPIO30B_H2F_A                 : out   std_logic;
          I2C0_SDA_MGPIO30B_H2F_B                 : out   std_logic;
          I2C1_SCL_MGPIO1A_H2F_A                  : out   std_logic;
          I2C1_SCL_MGPIO1A_H2F_B                  : out   std_logic;
          I2C1_SDA_MGPIO0A_H2F_A                  : out   std_logic;
          I2C1_SDA_MGPIO0A_H2F_B                  : out   std_logic;
          MDCF                                    : out   std_logic;
          MDOENF                                  : out   std_logic;
          MDOF                                    : out   std_logic;
          MMUART0_CTS_MGPIO19B_H2F_A              : out   std_logic;
          MMUART0_CTS_MGPIO19B_H2F_B              : out   std_logic;
          MMUART0_DCD_MGPIO22B_H2F_A              : out   std_logic;
          MMUART0_DCD_MGPIO22B_H2F_B              : out   std_logic;
          MMUART0_DSR_MGPIO20B_H2F_A              : out   std_logic;
          MMUART0_DSR_MGPIO20B_H2F_B              : out   std_logic;
          MMUART0_DTR_MGPIO18B_H2F_A              : out   std_logic;
          MMUART0_DTR_MGPIO18B_H2F_B              : out   std_logic;
          MMUART0_RI_MGPIO21B_H2F_A               : out   std_logic;
          MMUART0_RI_MGPIO21B_H2F_B               : out   std_logic;
          MMUART0_RTS_MGPIO17B_H2F_A              : out   std_logic;
          MMUART0_RTS_MGPIO17B_H2F_B              : out   std_logic;
          MMUART0_RXD_MGPIO28B_H2F_A              : out   std_logic;
          MMUART0_RXD_MGPIO28B_H2F_B              : out   std_logic;
          MMUART0_SCK_MGPIO29B_H2F_A              : out   std_logic;
          MMUART0_SCK_MGPIO29B_H2F_B              : out   std_logic;
          MMUART0_TXD_MGPIO27B_H2F_A              : out   std_logic;
          MMUART0_TXD_MGPIO27B_H2F_B              : out   std_logic;
          MMUART1_DTR_MGPIO12B_H2F_A              : out   std_logic;
          MMUART1_RTS_MGPIO11B_H2F_A              : out   std_logic;
          MMUART1_RTS_MGPIO11B_H2F_B              : out   std_logic;
          MMUART1_RXD_MGPIO26B_H2F_A              : out   std_logic;
          MMUART1_RXD_MGPIO26B_H2F_B              : out   std_logic;
          MMUART1_SCK_MGPIO25B_H2F_A              : out   std_logic;
          MMUART1_SCK_MGPIO25B_H2F_B              : out   std_logic;
          MMUART1_TXD_MGPIO24B_H2F_A              : out   std_logic;
          MMUART1_TXD_MGPIO24B_H2F_B              : out   std_logic;
          MPLL_LOCK                               : out   std_logic;
          PER2_FABRIC_PADDR                       : out   std_logic_vector(15 downto 2);
          PER2_FABRIC_PENABLE                     : out   std_logic;
          PER2_FABRIC_PSEL                        : out   std_logic;
          PER2_FABRIC_PWDATA                      : out   std_logic_vector(31 downto 0);
          PER2_FABRIC_PWRITE                      : out   std_logic;
          RTC_MATCH                               : out   std_logic;
          SLEEPDEEP                               : out   std_logic;
          SLEEPHOLDACK                            : out   std_logic;
          SLEEPING                                : out   std_logic;
          SMBALERT_NO0                            : out   std_logic;
          SMBALERT_NO1                            : out   std_logic;
          SMBSUS_NO0                              : out   std_logic;
          SMBSUS_NO1                              : out   std_logic;
          SPI0_CLK_OUT                            : out   std_logic;
          SPI0_SDI_MGPIO5A_H2F_A                  : out   std_logic;
          SPI0_SDI_MGPIO5A_H2F_B                  : out   std_logic;
          SPI0_SDO_MGPIO6A_H2F_A                  : out   std_logic;
          SPI0_SDO_MGPIO6A_H2F_B                  : out   std_logic;
          SPI0_SS0_MGPIO7A_H2F_A                  : out   std_logic;
          SPI0_SS0_MGPIO7A_H2F_B                  : out   std_logic;
          SPI0_SS1_MGPIO8A_H2F_A                  : out   std_logic;
          SPI0_SS1_MGPIO8A_H2F_B                  : out   std_logic;
          SPI0_SS2_MGPIO9A_H2F_A                  : out   std_logic;
          SPI0_SS2_MGPIO9A_H2F_B                  : out   std_logic;
          SPI0_SS3_MGPIO10A_H2F_A                 : out   std_logic;
          SPI0_SS3_MGPIO10A_H2F_B                 : out   std_logic;
          SPI0_SS4_MGPIO19A_H2F_A                 : out   std_logic;
          SPI0_SS5_MGPIO20A_H2F_A                 : out   std_logic;
          SPI0_SS6_MGPIO21A_H2F_A                 : out   std_logic;
          SPI0_SS7_MGPIO22A_H2F_A                 : out   std_logic;
          SPI1_CLK_OUT                            : out   std_logic;
          SPI1_SDI_MGPIO11A_H2F_A                 : out   std_logic;
          SPI1_SDI_MGPIO11A_H2F_B                 : out   std_logic;
          SPI1_SDO_MGPIO12A_H2F_A                 : out   std_logic;
          SPI1_SDO_MGPIO12A_H2F_B                 : out   std_logic;
          SPI1_SS0_MGPIO13A_H2F_A                 : out   std_logic;
          SPI1_SS0_MGPIO13A_H2F_B                 : out   std_logic;
          SPI1_SS1_MGPIO14A_H2F_A                 : out   std_logic;
          SPI1_SS1_MGPIO14A_H2F_B                 : out   std_logic;
          SPI1_SS2_MGPIO15A_H2F_A                 : out   std_logic;
          SPI1_SS2_MGPIO15A_H2F_B                 : out   std_logic;
          SPI1_SS3_MGPIO16A_H2F_A                 : out   std_logic;
          SPI1_SS3_MGPIO16A_H2F_B                 : out   std_logic;
          SPI1_SS4_MGPIO17A_H2F_A                 : out   std_logic;
          SPI1_SS5_MGPIO18A_H2F_A                 : out   std_logic;
          SPI1_SS6_MGPIO23A_H2F_A                 : out   std_logic;
          SPI1_SS7_MGPIO24A_H2F_A                 : out   std_logic;
          TCGF                                    : out   std_logic_vector(9 downto 0);
          TRACECLK                                : out   std_logic;
          TRACEDATA                               : out   std_logic_vector(3 downto 0);
          TX_CLK                                  : out   std_logic;
          TX_ENF                                  : out   std_logic;
          TX_ERRF                                 : out   std_logic;
          TXCTL_EN_RIF                            : out   std_logic;
          TXD_RIF                                 : out   std_logic_vector(3 downto 0);
          TXDF                                    : out   std_logic_vector(7 downto 0);
          TXEV                                    : out   std_logic;
          WDOGTIMEOUT                             : out   std_logic;
          F_ARREADY_HREADYOUT1                    : out   std_logic;
          F_AWREADY_HREADYOUT0                    : out   std_logic;
          F_BID                                   : out   std_logic_vector(3 downto 0);
          F_BRESP_HRESP0                          : out   std_logic_vector(1 downto 0);
          F_BVALID                                : out   std_logic;
          F_RDATA_HRDATA01                        : out   std_logic_vector(63 downto 0);
          F_RID                                   : out   std_logic_vector(3 downto 0);
          F_RLAST                                 : out   std_logic;
          F_RRESP_HRESP1                          : out   std_logic_vector(1 downto 0);
          F_RVALID                                : out   std_logic;
          F_WREADY                                : out   std_logic;
          MDDR_FABRIC_PRDATA                      : out   std_logic_vector(15 downto 0);
          MDDR_FABRIC_PREADY                      : out   std_logic;
          MDDR_FABRIC_PSLVERR                     : out   std_logic;
          CAN_RXBUS_F2H_SCP                       : in    std_logic := 'U';
          CAN_TX_EBL_F2H_SCP                      : in    std_logic := 'U';
          CAN_TXBUS_F2H_SCP                       : in    std_logic := 'U';
          COLF                                    : in    std_logic := 'U';
          CRSF                                    : in    std_logic := 'U';
          F2_DMAREADY                             : in    std_logic_vector(1 downto 0) := (others => 'U');
          F2H_INTERRUPT                           : in    std_logic_vector(15 downto 0) := (others => 'U');
          F2HCALIB                                : in    std_logic := 'U';
          F_DMAREADY                              : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_FM0_ADDR                              : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_FM0_ENABLE                            : in    std_logic := 'U';
          F_FM0_MASTLOCK                          : in    std_logic := 'U';
          F_FM0_READY                             : in    std_logic := 'U';
          F_FM0_SEL                               : in    std_logic := 'U';
          F_FM0_SIZE                              : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_FM0_TRANS1                            : in    std_logic := 'U';
          F_FM0_WDATA                             : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_FM0_WRITE                             : in    std_logic := 'U';
          F_HM0_RDATA                             : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_HM0_READY                             : in    std_logic := 'U';
          F_HM0_RESP                              : in    std_logic := 'U';
          FAB_AVALID                              : in    std_logic := 'U';
          FAB_HOSTDISCON                          : in    std_logic := 'U';
          FAB_IDDIG                               : in    std_logic := 'U';
          FAB_LINESTATE                           : in    std_logic_vector(1 downto 0) := (others => 'U');
          FAB_M3_RESET_N                          : in    std_logic := 'U';
          FAB_PLL_LOCK                            : in    std_logic := 'U';
          FAB_RXACTIVE                            : in    std_logic := 'U';
          FAB_RXERROR                             : in    std_logic := 'U';
          FAB_RXVALID                             : in    std_logic := 'U';
          FAB_RXVALIDH                            : in    std_logic := 'U';
          FAB_SESSEND                             : in    std_logic := 'U';
          FAB_TXREADY                             : in    std_logic := 'U';
          FAB_VBUSVALID                           : in    std_logic := 'U';
          FAB_VSTATUS                             : in    std_logic_vector(7 downto 0) := (others => 'U');
          FAB_XDATAIN                             : in    std_logic_vector(7 downto 0) := (others => 'U');
          GTX_CLKPF                               : in    std_logic := 'U';
          I2C0_BCLK                               : in    std_logic := 'U';
          I2C0_SCL_F2H_SCP                        : in    std_logic := 'U';
          I2C0_SDA_F2H_SCP                        : in    std_logic := 'U';
          I2C1_BCLK                               : in    std_logic := 'U';
          I2C1_SCL_F2H_SCP                        : in    std_logic := 'U';
          I2C1_SDA_F2H_SCP                        : in    std_logic := 'U';
          MDIF                                    : in    std_logic := 'U';
          MGPIO0A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO10A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO11A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO11B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO12A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO13A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO14A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO15A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO16A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO17B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO18B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO19B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO1A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO20B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO21B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO22B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO24B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO25B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO26B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO27B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO28B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO29B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO2A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO30B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO31B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO3A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO4A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO5A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO6A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO7A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO8A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO9A_F2H_GPIN                        : in    std_logic := 'U';
          MMUART0_CTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DCD_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DSR_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DTR_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_RI_F2H_SCP                      : in    std_logic := 'U';
          MMUART0_RTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_RXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_SCK_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_TXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_CTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_DCD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_DSR_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_RI_F2H_SCP                      : in    std_logic := 'U';
          MMUART1_RTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_RXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_SCK_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_TXD_F2H_SCP                     : in    std_logic := 'U';
          PER2_FABRIC_PRDATA                      : in    std_logic_vector(31 downto 0) := (others => 'U');
          PER2_FABRIC_PREADY                      : in    std_logic := 'U';
          PER2_FABRIC_PSLVERR                     : in    std_logic := 'U';
          RCGF                                    : in    std_logic_vector(9 downto 0) := (others => 'U');
          RX_CLKPF                                : in    std_logic := 'U';
          RX_DVF                                  : in    std_logic := 'U';
          RX_ERRF                                 : in    std_logic := 'U';
          RX_EV                                   : in    std_logic := 'U';
          RXDF                                    : in    std_logic_vector(7 downto 0) := (others => 'U');
          SLEEPHOLDREQ                            : in    std_logic := 'U';
          SMBALERT_NI0                            : in    std_logic := 'U';
          SMBALERT_NI1                            : in    std_logic := 'U';
          SMBSUS_NI0                              : in    std_logic := 'U';
          SMBSUS_NI1                              : in    std_logic := 'U';
          SPI0_CLK_IN                             : in    std_logic := 'U';
          SPI0_SDI_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SDO_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS0_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS1_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS2_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS3_F2H_SCP                        : in    std_logic := 'U';
          SPI1_CLK_IN                             : in    std_logic := 'U';
          SPI1_SDI_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SDO_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS0_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS1_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS2_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS3_F2H_SCP                        : in    std_logic := 'U';
          TX_CLKPF                                : in    std_logic := 'U';
          USER_MSS_GPIO_RESET_N                   : in    std_logic := 'U';
          USER_MSS_RESET_N                        : in    std_logic := 'U';
          XCLK_FAB                                : in    std_logic := 'U';
          CLK_BASE                                : in    std_logic := 'U';
          CLK_MDDR_APB                            : in    std_logic := 'U';
          F_ARADDR_HADDR1                         : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_ARBURST_HTRANS1                       : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARID_HSEL1                            : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_ARLEN_HBURST1                         : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_ARLOCK_HMASTLOCK1                     : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARSIZE_HSIZE1                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARVALID_HWRITE1                       : in    std_logic := 'U';
          F_AWADDR_HADDR0                         : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_AWBURST_HTRANS0                       : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWID_HSEL0                            : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_AWLEN_HBURST0                         : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_AWLOCK_HMASTLOCK0                     : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWSIZE_HSIZE0                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWVALID_HWRITE0                       : in    std_logic := 'U';
          F_BREADY                                : in    std_logic := 'U';
          F_RMW_AXI                               : in    std_logic := 'U';
          F_RREADY                                : in    std_logic := 'U';
          F_WDATA_HWDATA01                        : in    std_logic_vector(63 downto 0) := (others => 'U');
          F_WID_HREADY01                          : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_WLAST                                 : in    std_logic := 'U';
          F_WSTRB                                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          F_WVALID                                : in    std_logic := 'U';
          FPGA_MDDR_ARESET_N                      : in    std_logic := 'U';
          MDDR_FABRIC_PADDR                       : in    std_logic_vector(10 downto 2) := (others => 'U');
          MDDR_FABRIC_PENABLE                     : in    std_logic := 'U';
          MDDR_FABRIC_PSEL                        : in    std_logic := 'U';
          MDDR_FABRIC_PWDATA                      : in    std_logic_vector(15 downto 0) := (others => 'U');
          MDDR_FABRIC_PWRITE                      : in    std_logic := 'U';
          PRESET_N                                : in    std_logic := 'U';
          CAN_RXBUS_USBA_DATA1_MGPIO3A_IN         : in    std_logic := 'U';
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN        : in    std_logic := 'U';
          CAN_TXBUS_USBA_DATA0_MGPIO2A_IN         : in    std_logic := 'U';
          DM_IN                                   : in    std_logic_vector(2 downto 0) := (others => 'U');
          DRAM_DQ_IN                              : in    std_logic_vector(17 downto 0) := (others => 'U');
          DRAM_DQS_IN                             : in    std_logic_vector(2 downto 0) := (others => 'U');
          DRAM_FIFO_WE_IN                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          I2C0_SCL_USBC_DATA1_MGPIO31B_IN         : in    std_logic := 'U';
          I2C0_SDA_USBC_DATA0_MGPIO30B_IN         : in    std_logic := 'U';
          I2C1_SCL_USBA_DATA4_MGPIO1A_IN          : in    std_logic := 'U';
          I2C1_SDA_USBA_DATA3_MGPIO0A_IN          : in    std_logic := 'U';
          MGPIO0B_IN                              : in    std_logic := 'U';
          MGPIO10B_IN                             : in    std_logic := 'U';
          MGPIO1B_IN                              : in    std_logic := 'U';
          MGPIO25A_IN                             : in    std_logic := 'U';
          MGPIO26A_IN                             : in    std_logic := 'U';
          MGPIO27A_IN                             : in    std_logic := 'U';
          MGPIO28A_IN                             : in    std_logic := 'U';
          MGPIO29A_IN                             : in    std_logic := 'U';
          MGPIO2B_IN                              : in    std_logic := 'U';
          MGPIO30A_IN                             : in    std_logic := 'U';
          MGPIO31A_IN                             : in    std_logic := 'U';
          MGPIO3B_IN                              : in    std_logic := 'U';
          MGPIO4B_IN                              : in    std_logic := 'U';
          MGPIO5B_IN                              : in    std_logic := 'U';
          MGPIO6B_IN                              : in    std_logic := 'U';
          MGPIO7B_IN                              : in    std_logic := 'U';
          MGPIO8B_IN                              : in    std_logic := 'U';
          MGPIO9B_IN                              : in    std_logic := 'U';
          MMUART0_CTS_USBC_DATA7_MGPIO19B_IN      : in    std_logic := 'U';
          MMUART0_DCD_MGPIO22B_IN                 : in    std_logic := 'U';
          MMUART0_DSR_MGPIO20B_IN                 : in    std_logic := 'U';
          MMUART0_DTR_USBC_DATA6_MGPIO18B_IN      : in    std_logic := 'U';
          MMUART0_RI_MGPIO21B_IN                  : in    std_logic := 'U';
          MMUART0_RTS_USBC_DATA5_MGPIO17B_IN      : in    std_logic := 'U';
          MMUART0_RXD_USBC_STP_MGPIO28B_IN        : in    std_logic := 'U';
          MMUART0_SCK_USBC_NXT_MGPIO29B_IN        : in    std_logic := 'U';
          MMUART0_TXD_USBC_DIR_MGPIO27B_IN        : in    std_logic := 'U';
          MMUART1_CTS_MGPIO13B_IN                 : in    std_logic := 'U';
          MMUART1_DCD_MGPIO16B_IN                 : in    std_logic := 'U';
          MMUART1_DSR_MGPIO14B_IN                 : in    std_logic := 'U';
          MMUART1_DTR_MGPIO12B_IN                 : in    std_logic := 'U';
          MMUART1_RI_MGPIO15B_IN                  : in    std_logic := 'U';
          MMUART1_RTS_MGPIO11B_IN                 : in    std_logic := 'U';
          MMUART1_RXD_USBC_DATA3_MGPIO26B_IN      : in    std_logic := 'U';
          MMUART1_SCK_USBC_DATA4_MGPIO25B_IN      : in    std_logic := 'U';
          MMUART1_TXD_USBC_DATA2_MGPIO24B_IN      : in    std_logic := 'U';
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN     : in    std_logic := 'U';
          RGMII_MDC_RMII_MDC_IN                   : in    std_logic := 'U';
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN      : in    std_logic := 'U';
          RGMII_RX_CLK_IN                         : in    std_logic := 'U';
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN  : in    std_logic := 'U';
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN      : in    std_logic := 'U';
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN      : in    std_logic := 'U';
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN     : in    std_logic := 'U';
          RGMII_RXD3_USBB_DATA4_IN                : in    std_logic := 'U';
          RGMII_TX_CLK_IN                         : in    std_logic := 'U';
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN     : in    std_logic := 'U';
          RGMII_TXD0_RMII_TXD0_USBB_DIR_IN        : in    std_logic := 'U';
          RGMII_TXD1_RMII_TXD1_USBB_STP_IN        : in    std_logic := 'U';
          RGMII_TXD2_USBB_DATA5_IN                : in    std_logic := 'U';
          RGMII_TXD3_USBB_DATA6_IN                : in    std_logic := 'U';
          SPI0_SCK_USBA_XCLK_IN                   : in    std_logic := 'U';
          SPI0_SDI_USBA_DIR_MGPIO5A_IN            : in    std_logic := 'U';
          SPI0_SDO_USBA_STP_MGPIO6A_IN            : in    std_logic := 'U';
          SPI0_SS0_USBA_NXT_MGPIO7A_IN            : in    std_logic := 'U';
          SPI0_SS1_USBA_DATA5_MGPIO8A_IN          : in    std_logic := 'U';
          SPI0_SS2_USBA_DATA6_MGPIO9A_IN          : in    std_logic := 'U';
          SPI0_SS3_USBA_DATA7_MGPIO10A_IN         : in    std_logic := 'U';
          SPI0_SS4_MGPIO19A_IN                    : in    std_logic := 'U';
          SPI0_SS5_MGPIO20A_IN                    : in    std_logic := 'U';
          SPI0_SS6_MGPIO21A_IN                    : in    std_logic := 'U';
          SPI0_SS7_MGPIO22A_IN                    : in    std_logic := 'U';
          SPI1_SCK_IN                             : in    std_logic := 'U';
          SPI1_SDI_MGPIO11A_IN                    : in    std_logic := 'U';
          SPI1_SDO_MGPIO12A_IN                    : in    std_logic := 'U';
          SPI1_SS0_MGPIO13A_IN                    : in    std_logic := 'U';
          SPI1_SS1_MGPIO14A_IN                    : in    std_logic := 'U';
          SPI1_SS2_MGPIO15A_IN                    : in    std_logic := 'U';
          SPI1_SS3_MGPIO16A_IN                    : in    std_logic := 'U';
          SPI1_SS4_MGPIO17A_IN                    : in    std_logic := 'U';
          SPI1_SS5_MGPIO18A_IN                    : in    std_logic := 'U';
          SPI1_SS6_MGPIO23A_IN                    : in    std_logic := 'U';
          SPI1_SS7_MGPIO24A_IN                    : in    std_logic := 'U';
          USBC_XCLK_IN                            : in    std_logic := 'U';
          USBD_DATA0_IN                           : in    std_logic := 'U';
          USBD_DATA1_IN                           : in    std_logic := 'U';
          USBD_DATA2_IN                           : in    std_logic := 'U';
          USBD_DATA3_IN                           : in    std_logic := 'U';
          USBD_DATA4_IN                           : in    std_logic := 'U';
          USBD_DATA5_IN                           : in    std_logic := 'U';
          USBD_DATA6_IN                           : in    std_logic := 'U';
          USBD_DATA7_MGPIO23B_IN                  : in    std_logic := 'U';
          USBD_DIR_IN                             : in    std_logic := 'U';
          USBD_NXT_IN                             : in    std_logic := 'U';
          USBD_STP_IN                             : in    std_logic := 'U';
          USBD_XCLK_IN                            : in    std_logic := 'U';
          CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT        : out   std_logic;
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT       : out   std_logic;
          CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT        : out   std_logic;
          DRAM_ADDR                               : out   std_logic_vector(15 downto 0);
          DRAM_BA                                 : out   std_logic_vector(2 downto 0);
          DRAM_CASN                               : out   std_logic;
          DRAM_CKE                                : out   std_logic;
          DRAM_CLK                                : out   std_logic;
          DRAM_CSN                                : out   std_logic;
          DRAM_DM_RDQS_OUT                        : out   std_logic_vector(2 downto 0);
          DRAM_DQ_OUT                             : out   std_logic_vector(17 downto 0);
          DRAM_DQS_OUT                            : out   std_logic_vector(2 downto 0);
          DRAM_FIFO_WE_OUT                        : out   std_logic_vector(1 downto 0);
          DRAM_ODT                                : out   std_logic;
          DRAM_RASN                               : out   std_logic;
          DRAM_RSTN                               : out   std_logic;
          DRAM_WEN                                : out   std_logic;
          I2C0_SCL_USBC_DATA1_MGPIO31B_OUT        : out   std_logic;
          I2C0_SDA_USBC_DATA0_MGPIO30B_OUT        : out   std_logic;
          I2C1_SCL_USBA_DATA4_MGPIO1A_OUT         : out   std_logic;
          I2C1_SDA_USBA_DATA3_MGPIO0A_OUT         : out   std_logic;
          MGPIO0B_OUT                             : out   std_logic;
          MGPIO10B_OUT                            : out   std_logic;
          MGPIO1B_OUT                             : out   std_logic;
          MGPIO25A_OUT                            : out   std_logic;
          MGPIO26A_OUT                            : out   std_logic;
          MGPIO27A_OUT                            : out   std_logic;
          MGPIO28A_OUT                            : out   std_logic;
          MGPIO29A_OUT                            : out   std_logic;
          MGPIO2B_OUT                             : out   std_logic;
          MGPIO30A_OUT                            : out   std_logic;
          MGPIO31A_OUT                            : out   std_logic;
          MGPIO3B_OUT                             : out   std_logic;
          MGPIO4B_OUT                             : out   std_logic;
          MGPIO5B_OUT                             : out   std_logic;
          MGPIO6B_OUT                             : out   std_logic;
          MGPIO7B_OUT                             : out   std_logic;
          MGPIO8B_OUT                             : out   std_logic;
          MGPIO9B_OUT                             : out   std_logic;
          MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT     : out   std_logic;
          MMUART0_DCD_MGPIO22B_OUT                : out   std_logic;
          MMUART0_DSR_MGPIO20B_OUT                : out   std_logic;
          MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT     : out   std_logic;
          MMUART0_RI_MGPIO21B_OUT                 : out   std_logic;
          MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT     : out   std_logic;
          MMUART0_RXD_USBC_STP_MGPIO28B_OUT       : out   std_logic;
          MMUART0_SCK_USBC_NXT_MGPIO29B_OUT       : out   std_logic;
          MMUART0_TXD_USBC_DIR_MGPIO27B_OUT       : out   std_logic;
          MMUART1_CTS_MGPIO13B_OUT                : out   std_logic;
          MMUART1_DCD_MGPIO16B_OUT                : out   std_logic;
          MMUART1_DSR_MGPIO14B_OUT                : out   std_logic;
          MMUART1_DTR_MGPIO12B_OUT                : out   std_logic;
          MMUART1_RI_MGPIO15B_OUT                 : out   std_logic;
          MMUART1_RTS_MGPIO11B_OUT                : out   std_logic;
          MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT     : out   std_logic;
          MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT     : out   std_logic;
          MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT     : out   std_logic;
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT    : out   std_logic;
          RGMII_MDC_RMII_MDC_OUT                  : out   std_logic;
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT     : out   std_logic;
          RGMII_RX_CLK_OUT                        : out   std_logic;
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT : out   std_logic;
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT     : out   std_logic;
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT     : out   std_logic;
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT    : out   std_logic;
          RGMII_RXD3_USBB_DATA4_OUT               : out   std_logic;
          RGMII_TX_CLK_OUT                        : out   std_logic;
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT    : out   std_logic;
          RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT       : out   std_logic;
          RGMII_TXD1_RMII_TXD1_USBB_STP_OUT       : out   std_logic;
          RGMII_TXD2_USBB_DATA5_OUT               : out   std_logic;
          RGMII_TXD3_USBB_DATA6_OUT               : out   std_logic;
          SPI0_SCK_USBA_XCLK_OUT                  : out   std_logic;
          SPI0_SDI_USBA_DIR_MGPIO5A_OUT           : out   std_logic;
          SPI0_SDO_USBA_STP_MGPIO6A_OUT           : out   std_logic;
          SPI0_SS0_USBA_NXT_MGPIO7A_OUT           : out   std_logic;
          SPI0_SS1_USBA_DATA5_MGPIO8A_OUT         : out   std_logic;
          SPI0_SS2_USBA_DATA6_MGPIO9A_OUT         : out   std_logic;
          SPI0_SS3_USBA_DATA7_MGPIO10A_OUT        : out   std_logic;
          SPI0_SS4_MGPIO19A_OUT                   : out   std_logic;
          SPI0_SS5_MGPIO20A_OUT                   : out   std_logic;
          SPI0_SS6_MGPIO21A_OUT                   : out   std_logic;
          SPI0_SS7_MGPIO22A_OUT                   : out   std_logic;
          SPI1_SCK_OUT                            : out   std_logic;
          SPI1_SDI_MGPIO11A_OUT                   : out   std_logic;
          SPI1_SDO_MGPIO12A_OUT                   : out   std_logic;
          SPI1_SS0_MGPIO13A_OUT                   : out   std_logic;
          SPI1_SS1_MGPIO14A_OUT                   : out   std_logic;
          SPI1_SS2_MGPIO15A_OUT                   : out   std_logic;
          SPI1_SS3_MGPIO16A_OUT                   : out   std_logic;
          SPI1_SS4_MGPIO17A_OUT                   : out   std_logic;
          SPI1_SS5_MGPIO18A_OUT                   : out   std_logic;
          SPI1_SS6_MGPIO23A_OUT                   : out   std_logic;
          SPI1_SS7_MGPIO24A_OUT                   : out   std_logic;
          USBC_XCLK_OUT                           : out   std_logic;
          USBD_DATA0_OUT                          : out   std_logic;
          USBD_DATA1_OUT                          : out   std_logic;
          USBD_DATA2_OUT                          : out   std_logic;
          USBD_DATA3_OUT                          : out   std_logic;
          USBD_DATA4_OUT                          : out   std_logic;
          USBD_DATA5_OUT                          : out   std_logic;
          USBD_DATA6_OUT                          : out   std_logic;
          USBD_DATA7_MGPIO23B_OUT                 : out   std_logic;
          USBD_DIR_OUT                            : out   std_logic;
          USBD_NXT_OUT                            : out   std_logic;
          USBD_STP_OUT                            : out   std_logic;
          USBD_XCLK_OUT                           : out   std_logic;
          CAN_RXBUS_USBA_DATA1_MGPIO3A_OE         : out   std_logic;
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE        : out   std_logic;
          CAN_TXBUS_USBA_DATA0_MGPIO2A_OE         : out   std_logic;
          DM_OE                                   : out   std_logic_vector(2 downto 0);
          DRAM_DQ_OE                              : out   std_logic_vector(17 downto 0);
          DRAM_DQS_OE                             : out   std_logic_vector(2 downto 0);
          I2C0_SCL_USBC_DATA1_MGPIO31B_OE         : out   std_logic;
          I2C0_SDA_USBC_DATA0_MGPIO30B_OE         : out   std_logic;
          I2C1_SCL_USBA_DATA4_MGPIO1A_OE          : out   std_logic;
          I2C1_SDA_USBA_DATA3_MGPIO0A_OE          : out   std_logic;
          MGPIO0B_OE                              : out   std_logic;
          MGPIO10B_OE                             : out   std_logic;
          MGPIO1B_OE                              : out   std_logic;
          MGPIO25A_OE                             : out   std_logic;
          MGPIO26A_OE                             : out   std_logic;
          MGPIO27A_OE                             : out   std_logic;
          MGPIO28A_OE                             : out   std_logic;
          MGPIO29A_OE                             : out   std_logic;
          MGPIO2B_OE                              : out   std_logic;
          MGPIO30A_OE                             : out   std_logic;
          MGPIO31A_OE                             : out   std_logic;
          MGPIO3B_OE                              : out   std_logic;
          MGPIO4B_OE                              : out   std_logic;
          MGPIO5B_OE                              : out   std_logic;
          MGPIO6B_OE                              : out   std_logic;
          MGPIO7B_OE                              : out   std_logic;
          MGPIO8B_OE                              : out   std_logic;
          MGPIO9B_OE                              : out   std_logic;
          MMUART0_CTS_USBC_DATA7_MGPIO19B_OE      : out   std_logic;
          MMUART0_DCD_MGPIO22B_OE                 : out   std_logic;
          MMUART0_DSR_MGPIO20B_OE                 : out   std_logic;
          MMUART0_DTR_USBC_DATA6_MGPIO18B_OE      : out   std_logic;
          MMUART0_RI_MGPIO21B_OE                  : out   std_logic;
          MMUART0_RTS_USBC_DATA5_MGPIO17B_OE      : out   std_logic;
          MMUART0_RXD_USBC_STP_MGPIO28B_OE        : out   std_logic;
          MMUART0_SCK_USBC_NXT_MGPIO29B_OE        : out   std_logic;
          MMUART0_TXD_USBC_DIR_MGPIO27B_OE        : out   std_logic;
          MMUART1_CTS_MGPIO13B_OE                 : out   std_logic;
          MMUART1_DCD_MGPIO16B_OE                 : out   std_logic;
          MMUART1_DSR_MGPIO14B_OE                 : out   std_logic;
          MMUART1_DTR_MGPIO12B_OE                 : out   std_logic;
          MMUART1_RI_MGPIO15B_OE                  : out   std_logic;
          MMUART1_RTS_MGPIO11B_OE                 : out   std_logic;
          MMUART1_RXD_USBC_DATA3_MGPIO26B_OE      : out   std_logic;
          MMUART1_SCK_USBC_DATA4_MGPIO25B_OE      : out   std_logic;
          MMUART1_TXD_USBC_DATA2_MGPIO24B_OE      : out   std_logic;
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE     : out   std_logic;
          RGMII_MDC_RMII_MDC_OE                   : out   std_logic;
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE      : out   std_logic;
          RGMII_RX_CLK_OE                         : out   std_logic;
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE  : out   std_logic;
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE      : out   std_logic;
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE      : out   std_logic;
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE     : out   std_logic;
          RGMII_RXD3_USBB_DATA4_OE                : out   std_logic;
          RGMII_TX_CLK_OE                         : out   std_logic;
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE     : out   std_logic;
          RGMII_TXD0_RMII_TXD0_USBB_DIR_OE        : out   std_logic;
          RGMII_TXD1_RMII_TXD1_USBB_STP_OE        : out   std_logic;
          RGMII_TXD2_USBB_DATA5_OE                : out   std_logic;
          RGMII_TXD3_USBB_DATA6_OE                : out   std_logic;
          SPI0_SCK_USBA_XCLK_OE                   : out   std_logic;
          SPI0_SDI_USBA_DIR_MGPIO5A_OE            : out   std_logic;
          SPI0_SDO_USBA_STP_MGPIO6A_OE            : out   std_logic;
          SPI0_SS0_USBA_NXT_MGPIO7A_OE            : out   std_logic;
          SPI0_SS1_USBA_DATA5_MGPIO8A_OE          : out   std_logic;
          SPI0_SS2_USBA_DATA6_MGPIO9A_OE          : out   std_logic;
          SPI0_SS3_USBA_DATA7_MGPIO10A_OE         : out   std_logic;
          SPI0_SS4_MGPIO19A_OE                    : out   std_logic;
          SPI0_SS5_MGPIO20A_OE                    : out   std_logic;
          SPI0_SS6_MGPIO21A_OE                    : out   std_logic;
          SPI0_SS7_MGPIO22A_OE                    : out   std_logic;
          SPI1_SCK_OE                             : out   std_logic;
          SPI1_SDI_MGPIO11A_OE                    : out   std_logic;
          SPI1_SDO_MGPIO12A_OE                    : out   std_logic;
          SPI1_SS0_MGPIO13A_OE                    : out   std_logic;
          SPI1_SS1_MGPIO14A_OE                    : out   std_logic;
          SPI1_SS2_MGPIO15A_OE                    : out   std_logic;
          SPI1_SS3_MGPIO16A_OE                    : out   std_logic;
          SPI1_SS4_MGPIO17A_OE                    : out   std_logic;
          SPI1_SS5_MGPIO18A_OE                    : out   std_logic;
          SPI1_SS6_MGPIO23A_OE                    : out   std_logic;
          SPI1_SS7_MGPIO24A_OE                    : out   std_logic;
          USBC_XCLK_OE                            : out   std_logic;
          USBD_DATA0_OE                           : out   std_logic;
          USBD_DATA1_OE                           : out   std_logic;
          USBD_DATA2_OE                           : out   std_logic;
          USBD_DATA3_OE                           : out   std_logic;
          USBD_DATA4_OE                           : out   std_logic;
          USBD_DATA5_OE                           : out   std_logic;
          USBD_DATA6_OE                           : out   std_logic;
          USBD_DATA7_MGPIO23B_OE                  : out   std_logic;
          USBD_DIR_OE                             : out   std_logic;
          USBD_NXT_OE                             : out   std_logic;
          USBD_STP_OE                             : out   std_logic;
          USBD_XCLK_OE                            : out   std_logic
        );
  end component;

  component OUTBUF_DIFF
    generic (IOSTD:string := "");

    port( D    : in    std_logic := 'U';
          PADP : out   std_logic;
          PADN : out   std_logic
        );
  end component;

    signal \CORECONFIGP_0_APB_S_PCLK\, FIC_2_APB_M_PCLK, 
        \CORECONFIGP_0_APB_S_PRESET_N\, CONFIG_PRESET_N, 
        VCC_net_1, \CORECONFIGP_0_MDDR_APBmslave_PRDATA[0]\, 
        GND_net_1, MSS_ADLIB_INST_SPI0_SS1_USBA_DATA5_MGPIO8A_OUT, 
        MSS_ADLIB_INST_SPI0_SS1_USBA_DATA5_MGPIO8A_OE, 
        SPI_0_SS0_PAD_Y, 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT, 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE, 
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT, 
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE, 
        SPI_0_DI_PAD_Y, SPI_0_CLK_PAD_Y, 
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT, 
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE, 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT, 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE, 
        MMUART_1_RXD_PAD_Y, MSS_ADLIB_INST_DRAM_WEN, 
        MSS_ADLIB_INST_DRAM_RSTN, MSS_ADLIB_INST_DRAM_RASN, 
        MSS_ADLIB_INST_DRAM_ODT, \DRAM_FIFO_WE_OUT_net_0[0]\, 
        MDDR_DQS_TMATCH_0_IN_PAD_Y, MDDR_DQS_1_PAD_Y, 
        \DRAM_DQS_OUT_net_0[1]\, \DRAM_DQS_OE_net_0[1]\, 
        MDDR_DQS_0_PAD_Y, \DRAM_DQS_OUT_net_0[0]\, 
        \DRAM_DQS_OE_net_0[0]\, MDDR_DQ_15_PAD_Y, 
        \DRAM_DQ_OUT_net_0[15]\, \DRAM_DQ_OE_net_0[15]\, 
        MDDR_DQ_14_PAD_Y, \DRAM_DQ_OUT_net_0[14]\, 
        \DRAM_DQ_OE_net_0[14]\, MDDR_DQ_13_PAD_Y, 
        \DRAM_DQ_OUT_net_0[13]\, \DRAM_DQ_OE_net_0[13]\, 
        MDDR_DQ_12_PAD_Y, \DRAM_DQ_OUT_net_0[12]\, 
        \DRAM_DQ_OE_net_0[12]\, MDDR_DQ_11_PAD_Y, 
        \DRAM_DQ_OUT_net_0[11]\, \DRAM_DQ_OE_net_0[11]\, 
        MDDR_DQ_10_PAD_Y, \DRAM_DQ_OUT_net_0[10]\, 
        \DRAM_DQ_OE_net_0[10]\, MDDR_DQ_9_PAD_Y, 
        \DRAM_DQ_OUT_net_0[9]\, \DRAM_DQ_OE_net_0[9]\, 
        MDDR_DQ_8_PAD_Y, \DRAM_DQ_OUT_net_0[8]\, 
        \DRAM_DQ_OE_net_0[8]\, MDDR_DQ_7_PAD_Y, 
        \DRAM_DQ_OUT_net_0[7]\, \DRAM_DQ_OE_net_0[7]\, 
        MDDR_DQ_6_PAD_Y, \DRAM_DQ_OUT_net_0[6]\, 
        \DRAM_DQ_OE_net_0[6]\, MDDR_DQ_5_PAD_Y, 
        \DRAM_DQ_OUT_net_0[5]\, \DRAM_DQ_OE_net_0[5]\, 
        MDDR_DQ_4_PAD_Y, \DRAM_DQ_OUT_net_0[4]\, 
        \DRAM_DQ_OE_net_0[4]\, MDDR_DQ_3_PAD_Y, 
        \DRAM_DQ_OUT_net_0[3]\, \DRAM_DQ_OE_net_0[3]\, 
        MDDR_DQ_2_PAD_Y, \DRAM_DQ_OUT_net_0[2]\, 
        \DRAM_DQ_OE_net_0[2]\, MDDR_DQ_1_PAD_Y, 
        \DRAM_DQ_OUT_net_0[1]\, \DRAM_DQ_OE_net_0[1]\, 
        MDDR_DQ_0_PAD_Y, \DRAM_DQ_OUT_net_0[0]\, 
        \DRAM_DQ_OE_net_0[0]\, MDDR_DM_RDQS_1_PAD_Y, 
        \DRAM_DM_RDQS_OUT_net_0[1]\, \DM_OE_net_0[1]\, 
        MDDR_DM_RDQS_0_PAD_Y, \DRAM_DM_RDQS_OUT_net_0[0]\, 
        \DM_OE_net_0[0]\, MSS_ADLIB_INST_DRAM_CSN, 
        MSS_ADLIB_INST_DRAM_CKE, MSS_ADLIB_INST_DRAM_CASN, 
        \DRAM_BA_net_0[2]\, \DRAM_BA_net_0[1]\, 
        \DRAM_BA_net_0[0]\, \DRAM_ADDR_net_0[15]\, 
        \DRAM_ADDR_net_0[14]\, \DRAM_ADDR_net_0[13]\, 
        \DRAM_ADDR_net_0[12]\, \DRAM_ADDR_net_0[11]\, 
        \DRAM_ADDR_net_0[10]\, \DRAM_ADDR_net_0[9]\, 
        \DRAM_ADDR_net_0[8]\, \DRAM_ADDR_net_0[7]\, 
        \DRAM_ADDR_net_0[6]\, \DRAM_ADDR_net_0[5]\, 
        \DRAM_ADDR_net_0[4]\, \DRAM_ADDR_net_0[3]\, 
        \DRAM_ADDR_net_0[2]\, \DRAM_ADDR_net_0[1]\, 
        \DRAM_ADDR_net_0[0]\, I2C_1_SDA_PAD_Y, 
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OUT, 
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OE, 
        I2C_1_SCL_PAD_Y, 
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OUT, 
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OE, 
        GPIO_GPIO_31_BI_PAD_Y, MSS_ADLIB_INST_MGPIO31A_OUT, 
        MSS_ADLIB_INST_MGPIO31A_OE, GPIO_GPIO_26_BI_PAD_Y, 
        MSS_ADLIB_INST_MGPIO26A_OUT, MSS_ADLIB_INST_MGPIO26A_OE, 
        GPIO_GPIO_25_BI_PAD_Y, MSS_ADLIB_INST_MGPIO25A_OUT, 
        MSS_ADLIB_INST_MGPIO25A_OE, 
        MSS_ADLIB_INST_SPI0_SS5_MGPIO20A_OUT, 
        GPIO_GPIO_18_BI_PAD_Y, 
        MSS_ADLIB_INST_SPI1_SS5_MGPIO18A_OUT, 
        MSS_ADLIB_INST_SPI1_SS5_MGPIO18A_OE, 
        GPIO_GPIO_17_BI_PAD_Y, 
        MSS_ADLIB_INST_SPI1_SS4_MGPIO17A_OUT, 
        MSS_ADLIB_INST_SPI1_SS4_MGPIO17A_OE, 
        GPIO_GPIO_16_BI_PAD_Y, 
        MSS_ADLIB_INST_MMUART1_DCD_MGPIO16B_OUT, 
        MSS_ADLIB_INST_MMUART1_DCD_MGPIO16B_OE, 
        GPIO_GPIO_15_BI_PAD_Y, 
        MSS_ADLIB_INST_MMUART1_RI_MGPIO15B_OUT, 
        MSS_ADLIB_INST_MMUART1_RI_MGPIO15B_OE, 
        GPIO_GPIO_14_BI_PAD_Y, 
        MSS_ADLIB_INST_MMUART1_DSR_MGPIO14B_OUT, 
        MSS_ADLIB_INST_MMUART1_DSR_MGPIO14B_OE, 
        GPIO_GPIO_12_BI_PAD_Y, 
        MSS_ADLIB_INST_MMUART1_DTR_MGPIO12B_OUT, 
        MSS_ADLIB_INST_MMUART1_DTR_MGPIO12B_OE, 
        GPIO_GPIO_4_BI_PAD_Y, 
        MSS_ADLIB_INST_CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT, 
        MSS_ADLIB_INST_CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE, 
        GPIO_GPIO_3_BI_PAD_Y, 
        MSS_ADLIB_INST_CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT, 
        MSS_ADLIB_INST_CAN_RXBUS_USBA_DATA1_MGPIO3A_OE, 
        GPIO_GPIO_0_BI_PAD_Y, MSS_ADLIB_INST_MGPIO0B_OUT, 
        MSS_ADLIB_INST_MGPIO0B_OE, MSS_ADLIB_INST_DRAM_CLK
         : std_logic;
    signal nc228, nc203, nc216, nc194, nc151, nc23, nc175, nc58, 
        nc116, nc74, nc133, nc238, nc167, nc84, nc39, nc72, nc212, 
        nc205, nc82, nc145, nc181, nc160, nc57, nc156, nc125, 
        nc211, nc73, nc107, nc66, nc83, nc9, nc171, nc54, nc135, 
        nc41, nc100, nc52, nc186, nc29, nc118, nc60, nc141, nc193, 
        nc214, nc240, nc45, nc53, nc121, nc176, nc220, nc158, 
        nc209, nc246, nc162, nc11, nc131, nc96, nc79, nc226, 
        nc146, nc230, nc89, nc119, nc48, nc213, nc126, nc195, 
        nc188, nc242, nc15, nc236, nc102, nc3, nc207, nc47, nc90, 
        nc222, nc159, nc136, nc241, nc178, nc215, nc59, nc221, 
        nc232, nc18, nc44, nc117, nc189, nc164, nc148, nc42, 
        nc231, nc191, nc17, nc2, nc110, nc128, nc244, nc43, nc179, 
        nc157, nc36, nc224, nc61, nc104, nc138, nc14, nc150, 
        nc196, nc234, nc149, nc12, nc219, nc30, nc243, nc187, 
        nc65, nc7, nc129, nc8, nc223, nc13, nc180, nc26, nc177, 
        nc139, nc245, nc233, nc163, nc112, nc68, nc49, nc217, 
        nc170, nc91, nc225, nc5, nc20, nc198, nc147, nc67, nc152, 
        nc127, nc103, nc235, nc76, nc208, nc140, nc86, nc95, 
        nc120, nc165, nc137, nc64, nc19, nc70, nc182, nc62, nc199, 
        nc80, nc130, nc98, nc114, nc56, nc105, nc63, nc172, nc229, 
        nc97, nc161, nc31, nc154, nc50, nc239, nc142, nc94, nc197, 
        nc122, nc35, nc4, nc227, nc92, nc101, nc184, nc200, nc190, 
        nc166, nc132, nc21, nc237, nc93, nc69, nc206, nc174, nc38, 
        nc113, nc218, nc106, nc25, nc1, nc37, nc202, nc144, nc153, 
        nc46, nc71, nc124, nc81, nc201, nc168, nc34, nc28, nc115, 
        nc192, nc134, nc32, nc40, nc99, nc75, nc183, nc85, nc27, 
        nc108, nc16, nc155, nc51, nc33, nc204, nc173, nc169, nc78, 
        nc24, nc88, nc111, nc55, nc10, nc22, nc210, nc185, nc143, 
        nc77, nc6, nc109, nc87, nc123 : std_logic;

begin 

    CORECONFIGP_0_APB_S_PRESET_N <= 
        \CORECONFIGP_0_APB_S_PRESET_N\;
    CORECONFIGP_0_APB_S_PCLK <= \CORECONFIGP_0_APB_S_PCLK\;

    MDDR_ADDR_6_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[6]\, PAD => MDDR_ADDR(6));
    
    MDDR_CAS_N_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => MSS_ADLIB_INST_DRAM_CASN, PAD => MDDR_CAS_N);
    
    MDDR_RESET_N_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => MSS_ADLIB_INST_DRAM_RSTN, PAD => MDDR_RESET_N);
    
    MDDR_ODT_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => MSS_ADLIB_INST_DRAM_ODT, PAD => MDDR_ODT);
    
    GPIO_GPIO_31_BI_PAD : BIBUF
      port map(PAD => GPIO_31_BI, D => 
        MSS_ADLIB_INST_MGPIO31A_OUT, E => 
        MSS_ADLIB_INST_MGPIO31A_OE, Y => GPIO_GPIO_31_BI_PAD_Y);
    
    MDDR_ADDR_11_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[11]\, PAD => MDDR_ADDR(11));
    
    MMUART_1_TXD_PAD : TRIBUFF
      port map(D => 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT, E => 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE, PAD
         => MMUART_1_TXD);
    
    MDDR_DQ_10_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(10), D => \DRAM_DQ_OUT_net_0[10]\, 
        E => \DRAM_DQ_OE_net_0[10]\, Y => MDDR_DQ_10_PAD_Y);
    
    FIC_2_APB_M_PRDATA_0_ret : SLE
      port map(D => \CORECONFIGP_0_MDDR_APBmslave_PRDATA[0]\, CLK
         => \CORECONFIGP_0_APB_S_PCLK\, EN => state_0, ALn => 
        \CORECONFIGP_0_APB_S_PRESET_N\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA_reto_0);
    
    MDDR_DQ_1_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(1), D => \DRAM_DQ_OUT_net_0[1]\, E
         => \DRAM_DQ_OE_net_0[1]\, Y => MDDR_DQ_1_PAD_Y);
    
    MDDR_ADDR_7_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[7]\, PAD => MDDR_ADDR(7));
    
    MDDR_DQ_11_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(11), D => \DRAM_DQ_OUT_net_0[11]\, 
        E => \DRAM_DQ_OE_net_0[11]\, Y => MDDR_DQ_11_PAD_Y);
    
    MDDR_DQ_9_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(9), D => \DRAM_DQ_OUT_net_0[9]\, E
         => \DRAM_DQ_OE_net_0[9]\, Y => MDDR_DQ_9_PAD_Y);
    
    MSS_ADLIB_INST_RNI1CJ7 : CLKINT
      port map(A => CONFIG_PRESET_N, Y => 
        \CORECONFIGP_0_APB_S_PRESET_N\);
    
    MDDR_DQ_3_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(3), D => \DRAM_DQ_OUT_net_0[3]\, E
         => \DRAM_DQ_OE_net_0[3]\, Y => MDDR_DQ_3_PAD_Y);
    
    GPIO_GPIO_25_BI_PAD : BIBUF
      port map(PAD => GPIO_25_BI, D => 
        MSS_ADLIB_INST_MGPIO25A_OUT, E => 
        MSS_ADLIB_INST_MGPIO25A_OE, Y => GPIO_GPIO_25_BI_PAD_Y);
    
    MDDR_DQ_0_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(0), D => \DRAM_DQ_OUT_net_0[0]\, E
         => \DRAM_DQ_OE_net_0[0]\, Y => MDDR_DQ_0_PAD_Y);
    
    MDDR_ADDR_12_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[12]\, PAD => MDDR_ADDR(12));
    
    GPIO_GPIO_17_BI_PAD : BIBUF
      port map(PAD => GPIO_17_BI, D => 
        MSS_ADLIB_INST_SPI1_SS4_MGPIO17A_OUT, E => 
        MSS_ADLIB_INST_SPI1_SS4_MGPIO17A_OE, Y => 
        GPIO_GPIO_17_BI_PAD_Y);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    MDDR_DQ_2_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(2), D => \DRAM_DQ_OUT_net_0[2]\, E
         => \DRAM_DQ_OE_net_0[2]\, Y => MDDR_DQ_2_PAD_Y);
    
    MDDR_DQ_12_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(12), D => \DRAM_DQ_OUT_net_0[12]\, 
        E => \DRAM_DQ_OE_net_0[12]\, Y => MDDR_DQ_12_PAD_Y);
    
    MDDR_CKE_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => MSS_ADLIB_INST_DRAM_CKE, PAD => MDDR_CKE);
    
    MDDR_ADDR_2_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[2]\, PAD => MDDR_ADDR(2));
    
    GPIO_GPIO_0_BI_PAD : BIBUF
      port map(PAD => GPIO_0_BI, D => MSS_ADLIB_INST_MGPIO0B_OUT, 
        E => MSS_ADLIB_INST_MGPIO0B_OE, Y => GPIO_GPIO_0_BI_PAD_Y);
    
    FIC_2_APB_M_PCLK_inferred_clock_RNIPG5_0 : CFG1
      generic map(INIT => "01")

      port map(A => \CORECONFIGP_0_APB_S_PCLK\, Y => 
        CORECONFIGP_0_APB_S_PCLK_i);
    
    MDDR_ADDR_13_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[13]\, PAD => MDDR_ADDR(13));
    
    I2C_1_SDA_PAD : BIBUF
      port map(PAD => I2C_1_SDA, D => 
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OUT, E => 
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OE, Y => 
        I2C_1_SDA_PAD_Y);
    
    I2C_1_SCL_PAD : BIBUF
      port map(PAD => I2C_1_SCL, D => 
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OUT, E => 
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OE, Y => 
        I2C_1_SCL_PAD_Y);
    
    MDDR_ADDR_5_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[5]\, PAD => MDDR_ADDR(5));
    
    MDDR_DM_RDQS_1_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DM_RDQS(1), D => 
        \DRAM_DM_RDQS_OUT_net_0[1]\, E => \DM_OE_net_0[1]\, Y => 
        MDDR_DM_RDQS_1_PAD_Y);
    
    GPIO_GPIO_12_BI_PAD : BIBUF
      port map(PAD => GPIO_12_BI, D => 
        MSS_ADLIB_INST_MMUART1_DTR_MGPIO12B_OUT, E => 
        MSS_ADLIB_INST_MMUART1_DTR_MGPIO12B_OE, Y => 
        GPIO_GPIO_12_BI_PAD_Y);
    
    SPI_0_DO_PAD : TRIBUFF
      port map(D => MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT, 
        E => MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE, PAD => 
        SPI_0_DO);
    
    MDDR_DQS_0_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQS(0), D => \DRAM_DQS_OUT_net_0[0]\, 
        E => \DRAM_DQS_OE_net_0[0]\, Y => MDDR_DQS_0_PAD_Y);
    
    MDDR_DQS_1_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQS(1), D => \DRAM_DQS_OUT_net_0[1]\, 
        E => \DRAM_DQS_OE_net_0[1]\, Y => MDDR_DQS_1_PAD_Y);
    
    MDDR_DQ_15_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(15), D => \DRAM_DQ_OUT_net_0[15]\, 
        E => \DRAM_DQ_OE_net_0[15]\, Y => MDDR_DQ_15_PAD_Y);
    
    MDDR_DM_RDQS_0_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DM_RDQS(0), D => 
        \DRAM_DM_RDQS_OUT_net_0[0]\, E => \DM_OE_net_0[0]\, Y => 
        MDDR_DM_RDQS_0_PAD_Y);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    SPI_0_DI_PAD : INBUF
      port map(PAD => SPI_0_DI, Y => SPI_0_DI_PAD_Y);
    
    MDDR_DQ_8_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(8), D => \DRAM_DQ_OUT_net_0[8]\, E
         => \DRAM_DQ_OE_net_0[8]\, Y => MDDR_DQ_8_PAD_Y);
    
    GPIO_GPIO_14_BI_PAD : BIBUF
      port map(PAD => GPIO_14_BI, D => 
        MSS_ADLIB_INST_MMUART1_DSR_MGPIO14B_OUT, E => 
        MSS_ADLIB_INST_MMUART1_DSR_MGPIO14B_OE, Y => 
        GPIO_GPIO_14_BI_PAD_Y);
    
    GPIO_GPIO_4_BI_PAD : BIBUF
      port map(PAD => GPIO_4_BI, D => 
        MSS_ADLIB_INST_CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT, E => 
        MSS_ADLIB_INST_CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE, Y => 
        GPIO_GPIO_4_BI_PAD_Y);
    
    MDDR_ADDR_9_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[9]\, PAD => MDDR_ADDR(9));
    
    MDDR_BA_2_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_BA_net_0[2]\, PAD => MDDR_BA(2));
    
    MDDR_ADDR_14_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[14]\, PAD => MDDR_ADDR(14));
    
    MSS_ADLIB_INST : MSS_060

              generic map(INIT => "00" & x"000000000000030000000000000003610008090A4290800908000000090A42000000000C03000000009000000000200012036190A4200001004000000000000000000000000000000000000F000000000000000000000000000000007FFFFFFFB000001007C35C804248006090801041A3FFFFE400000000000846809D001F0F41C000000025A00010842108421000001FE34001FF8000000400000000020CD1007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
         ACT_UBITS => x"FFFFFFFFFFFFFF",
         MEMORYFILE => "ENVM_init.mem", RTC_MAIN_XTL_FREQ => 0.0,
         DDR_CLK_FREQ => 142.0)

      port map(CAN_RXBUS_MGPIO3A_H2F_A => OPEN, 
        CAN_RXBUS_MGPIO3A_H2F_B => OPEN, CAN_TX_EBL_MGPIO4A_H2F_A
         => OPEN, CAN_TX_EBL_MGPIO4A_H2F_B => OPEN, 
        CAN_TXBUS_MGPIO2A_H2F_A => OPEN, CAN_TXBUS_MGPIO2A_H2F_B
         => OPEN, CLK_CONFIG_APB => FIC_2_APB_M_PCLK, COMMS_INT
         => OPEN, CONFIG_PRESET_N => CONFIG_PRESET_N, 
        EDAC_ERROR(7) => nc228, EDAC_ERROR(6) => nc203, 
        EDAC_ERROR(5) => nc216, EDAC_ERROR(4) => nc194, 
        EDAC_ERROR(3) => nc151, EDAC_ERROR(2) => nc23, 
        EDAC_ERROR(1) => nc175, EDAC_ERROR(0) => nc58, 
        F_FM0_RDATA(31) => nc116, F_FM0_RDATA(30) => nc74, 
        F_FM0_RDATA(29) => nc133, F_FM0_RDATA(28) => nc238, 
        F_FM0_RDATA(27) => nc167, F_FM0_RDATA(26) => nc84, 
        F_FM0_RDATA(25) => nc39, F_FM0_RDATA(24) => nc72, 
        F_FM0_RDATA(23) => nc212, F_FM0_RDATA(22) => nc205, 
        F_FM0_RDATA(21) => nc82, F_FM0_RDATA(20) => nc145, 
        F_FM0_RDATA(19) => nc181, F_FM0_RDATA(18) => nc160, 
        F_FM0_RDATA(17) => nc57, F_FM0_RDATA(16) => nc156, 
        F_FM0_RDATA(15) => nc125, F_FM0_RDATA(14) => nc211, 
        F_FM0_RDATA(13) => nc73, F_FM0_RDATA(12) => nc107, 
        F_FM0_RDATA(11) => nc66, F_FM0_RDATA(10) => nc83, 
        F_FM0_RDATA(9) => nc9, F_FM0_RDATA(8) => nc171, 
        F_FM0_RDATA(7) => nc54, F_FM0_RDATA(6) => nc135, 
        F_FM0_RDATA(5) => nc41, F_FM0_RDATA(4) => nc100, 
        F_FM0_RDATA(3) => nc52, F_FM0_RDATA(2) => nc186, 
        F_FM0_RDATA(1) => nc29, F_FM0_RDATA(0) => nc118, 
        F_FM0_READYOUT => OPEN, F_FM0_RESP => OPEN, 
        F_HM0_ADDR(31) => nc60, F_HM0_ADDR(30) => nc141, 
        F_HM0_ADDR(29) => nc193, F_HM0_ADDR(28) => nc214, 
        F_HM0_ADDR(27) => nc240, F_HM0_ADDR(26) => nc45, 
        F_HM0_ADDR(25) => nc53, F_HM0_ADDR(24) => nc121, 
        F_HM0_ADDR(23) => nc176, F_HM0_ADDR(22) => nc220, 
        F_HM0_ADDR(21) => nc158, F_HM0_ADDR(20) => nc209, 
        F_HM0_ADDR(19) => nc246, F_HM0_ADDR(18) => nc162, 
        F_HM0_ADDR(17) => nc11, F_HM0_ADDR(16) => nc131, 
        F_HM0_ADDR(15) => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(15), 
        F_HM0_ADDR(14) => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(14), 
        F_HM0_ADDR(13) => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(13), 
        F_HM0_ADDR(12) => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(12), 
        F_HM0_ADDR(11) => nc96, F_HM0_ADDR(10) => nc79, 
        F_HM0_ADDR(9) => nc226, F_HM0_ADDR(8) => nc146, 
        F_HM0_ADDR(7) => CoreAPB3_0_APBmslave0_PADDR(7), 
        F_HM0_ADDR(6) => CoreAPB3_0_APBmslave0_PADDR(6), 
        F_HM0_ADDR(5) => CoreAPB3_0_APBmslave0_PADDR(5), 
        F_HM0_ADDR(4) => CoreAPB3_0_APBmslave0_PADDR(4), 
        F_HM0_ADDR(3) => CoreAPB3_0_APBmslave0_PADDR(3), 
        F_HM0_ADDR(2) => CoreAPB3_0_APBmslave0_PADDR(2), 
        F_HM0_ADDR(1) => CoreAPB3_0_APBmslave0_PADDR(1), 
        F_HM0_ADDR(0) => CoreAPB3_0_APBmslave0_PADDR(0), 
        F_HM0_ENABLE => CoreAPB3_0_APBmslave0_PENABLE, F_HM0_SEL
         => m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx, F_HM0_SIZE(1)
         => nc230, F_HM0_SIZE(0) => nc89, F_HM0_TRANS1 => OPEN, 
        F_HM0_WDATA(31) => nc119, F_HM0_WDATA(30) => nc48, 
        F_HM0_WDATA(29) => nc213, F_HM0_WDATA(28) => nc126, 
        F_HM0_WDATA(27) => nc195, F_HM0_WDATA(26) => nc188, 
        F_HM0_WDATA(25) => nc242, F_HM0_WDATA(24) => nc15, 
        F_HM0_WDATA(23) => nc236, F_HM0_WDATA(22) => nc102, 
        F_HM0_WDATA(21) => nc3, F_HM0_WDATA(20) => nc207, 
        F_HM0_WDATA(19) => nc47, F_HM0_WDATA(18) => nc90, 
        F_HM0_WDATA(17) => nc222, F_HM0_WDATA(16) => nc159, 
        F_HM0_WDATA(15) => nc136, F_HM0_WDATA(14) => nc241, 
        F_HM0_WDATA(13) => nc178, F_HM0_WDATA(12) => nc215, 
        F_HM0_WDATA(11) => nc59, F_HM0_WDATA(10) => nc221, 
        F_HM0_WDATA(9) => nc232, F_HM0_WDATA(8) => nc18, 
        F_HM0_WDATA(7) => CoreAPB3_0_APBmslave0_PWDATA(7), 
        F_HM0_WDATA(6) => CoreAPB3_0_APBmslave0_PWDATA(6), 
        F_HM0_WDATA(5) => CoreAPB3_0_APBmslave0_PWDATA(5), 
        F_HM0_WDATA(4) => CoreAPB3_0_APBmslave0_PWDATA(4), 
        F_HM0_WDATA(3) => CoreAPB3_0_APBmslave0_PWDATA(3), 
        F_HM0_WDATA(2) => CoreAPB3_0_APBmslave0_PWDATA(2), 
        F_HM0_WDATA(1) => CoreAPB3_0_APBmslave0_PWDATA(1), 
        F_HM0_WDATA(0) => CoreAPB3_0_APBmslave0_PWDATA(0), 
        F_HM0_WRITE => CoreAPB3_0_APBmslave0_PWRITE, FAB_CHRGVBUS
         => OPEN, FAB_DISCHRGVBUS => OPEN, FAB_DMPULLDOWN => OPEN, 
        FAB_DPPULLDOWN => OPEN, FAB_DRVVBUS => OPEN, FAB_IDPULLUP
         => OPEN, FAB_OPMODE(1) => nc44, FAB_OPMODE(0) => nc117, 
        FAB_SUSPENDM => OPEN, FAB_TERMSEL => OPEN, FAB_TXVALID
         => OPEN, FAB_VCONTROL(3) => nc189, FAB_VCONTROL(2) => 
        nc164, FAB_VCONTROL(1) => nc148, FAB_VCONTROL(0) => nc42, 
        FAB_VCONTROLLOADM => OPEN, FAB_XCVRSEL(1) => nc231, 
        FAB_XCVRSEL(0) => nc191, FAB_XDATAOUT(7) => nc17, 
        FAB_XDATAOUT(6) => nc2, FAB_XDATAOUT(5) => nc110, 
        FAB_XDATAOUT(4) => nc128, FAB_XDATAOUT(3) => nc244, 
        FAB_XDATAOUT(2) => nc43, FAB_XDATAOUT(1) => nc179, 
        FAB_XDATAOUT(0) => nc157, FACC_GLMUX_SEL => OPEN, 
        FIC32_0_MASTER(1) => nc36, FIC32_0_MASTER(0) => nc224, 
        FIC32_1_MASTER(1) => nc61, FIC32_1_MASTER(0) => nc104, 
        FPGA_RESET_N => m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        GTX_CLK => OPEN, H2F_INTERRUPT(15) => nc138, 
        H2F_INTERRUPT(14) => nc14, H2F_INTERRUPT(13) => nc150, 
        H2F_INTERRUPT(12) => nc196, H2F_INTERRUPT(11) => nc234, 
        H2F_INTERRUPT(10) => nc149, H2F_INTERRUPT(9) => nc12, 
        H2F_INTERRUPT(8) => nc219, H2F_INTERRUPT(7) => nc30, 
        H2F_INTERRUPT(6) => nc243, H2F_INTERRUPT(5) => nc187, 
        H2F_INTERRUPT(4) => nc65, H2F_INTERRUPT(3) => nc7, 
        H2F_INTERRUPT(2) => nc129, H2F_INTERRUPT(1) => nc8, 
        H2F_INTERRUPT(0) => nc223, H2F_NMI => OPEN, H2FCALIB => 
        OPEN, I2C0_SCL_MGPIO31B_H2F_A => OPEN, 
        I2C0_SCL_MGPIO31B_H2F_B => OPEN, I2C0_SDA_MGPIO30B_H2F_A
         => OPEN, I2C0_SDA_MGPIO30B_H2F_B => OPEN, 
        I2C1_SCL_MGPIO1A_H2F_A => 
        m2s010_som_sb_MSS_0_GPIO_1_M2F_OE, I2C1_SCL_MGPIO1A_H2F_B
         => GPIO_1_M2F, I2C1_SDA_MGPIO0A_H2F_A => OPEN, 
        I2C1_SDA_MGPIO0A_H2F_B => OPEN, MDCF => MAC_MII_MDC_c, 
        MDOENF => m2s010_som_sb_MSS_0_MAC_MII_MDO_EN, MDOF => 
        m2s010_som_sb_MSS_0_MAC_MII_MDO, 
        MMUART0_CTS_MGPIO19B_H2F_A => OPEN, 
        MMUART0_CTS_MGPIO19B_H2F_B => OPEN, 
        MMUART0_DCD_MGPIO22B_H2F_A => OPEN, 
        MMUART0_DCD_MGPIO22B_H2F_B => GPIO_22_M2F_c, 
        MMUART0_DSR_MGPIO20B_H2F_A => OPEN, 
        MMUART0_DSR_MGPIO20B_H2F_B => OPEN, 
        MMUART0_DTR_MGPIO18B_H2F_A => OPEN, 
        MMUART0_DTR_MGPIO18B_H2F_B => OPEN, 
        MMUART0_RI_MGPIO21B_H2F_A => OPEN, 
        MMUART0_RI_MGPIO21B_H2F_B => GPIO_21_M2F_c, 
        MMUART0_RTS_MGPIO17B_H2F_A => OPEN, 
        MMUART0_RTS_MGPIO17B_H2F_B => OPEN, 
        MMUART0_RXD_MGPIO28B_H2F_A => OPEN, 
        MMUART0_RXD_MGPIO28B_H2F_B => 
        m2s010_som_sb_0_GPIO_28_SW_RESET, 
        MMUART0_SCK_MGPIO29B_H2F_A => OPEN, 
        MMUART0_SCK_MGPIO29B_H2F_B => OPEN, 
        MMUART0_TXD_MGPIO27B_H2F_A => MMUART_0_TXD_M2F_c, 
        MMUART0_TXD_MGPIO27B_H2F_B => OPEN, 
        MMUART1_DTR_MGPIO12B_H2F_A => OPEN, 
        MMUART1_RTS_MGPIO11B_H2F_A => OPEN, 
        MMUART1_RTS_MGPIO11B_H2F_B => OPEN, 
        MMUART1_RXD_MGPIO26B_H2F_A => OPEN, 
        MMUART1_RXD_MGPIO26B_H2F_B => OPEN, 
        MMUART1_SCK_MGPIO25B_H2F_A => OPEN, 
        MMUART1_SCK_MGPIO25B_H2F_B => OPEN, 
        MMUART1_TXD_MGPIO24B_H2F_A => OPEN, 
        MMUART1_TXD_MGPIO24B_H2F_B => GPIO_24_M2F_c, MPLL_LOCK
         => OPEN, PER2_FABRIC_PADDR(15) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(15), 
        PER2_FABRIC_PADDR(14) => nc13, PER2_FABRIC_PADDR(13) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(13), 
        PER2_FABRIC_PADDR(12) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(12), 
        PER2_FABRIC_PADDR(11) => nc180, PER2_FABRIC_PADDR(10) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(10), 
        PER2_FABRIC_PADDR(9) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(9), 
        PER2_FABRIC_PADDR(8) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(8), 
        PER2_FABRIC_PADDR(7) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(7), 
        PER2_FABRIC_PADDR(6) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(6), 
        PER2_FABRIC_PADDR(5) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(5), 
        PER2_FABRIC_PADDR(4) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), 
        PER2_FABRIC_PADDR(3) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), 
        PER2_FABRIC_PADDR(2) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), 
        PER2_FABRIC_PENABLE => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE, 
        PER2_FABRIC_PSEL => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx, 
        PER2_FABRIC_PWDATA(31) => nc26, PER2_FABRIC_PWDATA(30)
         => nc177, PER2_FABRIC_PWDATA(29) => nc139, 
        PER2_FABRIC_PWDATA(28) => nc245, PER2_FABRIC_PWDATA(27)
         => nc233, PER2_FABRIC_PWDATA(26) => nc163, 
        PER2_FABRIC_PWDATA(25) => nc112, PER2_FABRIC_PWDATA(24)
         => nc68, PER2_FABRIC_PWDATA(23) => nc49, 
        PER2_FABRIC_PWDATA(22) => nc217, PER2_FABRIC_PWDATA(21)
         => nc170, PER2_FABRIC_PWDATA(20) => nc91, 
        PER2_FABRIC_PWDATA(19) => nc225, PER2_FABRIC_PWDATA(18)
         => nc5, PER2_FABRIC_PWDATA(17) => nc20, 
        PER2_FABRIC_PWDATA(16) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(16), 
        PER2_FABRIC_PWDATA(15) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(15), 
        PER2_FABRIC_PWDATA(14) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(14), 
        PER2_FABRIC_PWDATA(13) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(13), 
        PER2_FABRIC_PWDATA(12) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(12), 
        PER2_FABRIC_PWDATA(11) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(11), 
        PER2_FABRIC_PWDATA(10) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(10), 
        PER2_FABRIC_PWDATA(9) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(9), 
        PER2_FABRIC_PWDATA(8) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(8), 
        PER2_FABRIC_PWDATA(7) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(7), 
        PER2_FABRIC_PWDATA(6) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(6), 
        PER2_FABRIC_PWDATA(5) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(5), 
        PER2_FABRIC_PWDATA(4) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(4), 
        PER2_FABRIC_PWDATA(3) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(3), 
        PER2_FABRIC_PWDATA(2) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(2), 
        PER2_FABRIC_PWDATA(1) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(1), 
        PER2_FABRIC_PWDATA(0) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(0), 
        PER2_FABRIC_PWRITE => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE, 
        RTC_MATCH => OPEN, SLEEPDEEP => OPEN, SLEEPHOLDACK => 
        OPEN, SLEEPING => OPEN, SMBALERT_NO0 => OPEN, 
        SMBALERT_NO1 => OPEN, SMBSUS_NO0 => OPEN, SMBSUS_NO1 => 
        OPEN, SPI0_CLK_OUT => OPEN, SPI0_SDI_MGPIO5A_H2F_A => 
        OPEN, SPI0_SDI_MGPIO5A_H2F_B => GPIO_5_M2F_c, 
        SPI0_SDO_MGPIO6A_H2F_A => 
        m2s010_som_sb_MSS_0_GPIO_6_M2F_OE, SPI0_SDO_MGPIO6A_H2F_B
         => m2s010_som_sb_MSS_0_GPIO_6_M2F, 
        SPI0_SS0_MGPIO7A_H2F_A => 
        m2s010_som_sb_MSS_0_GPIO_7_M2F_OE, SPI0_SS0_MGPIO7A_H2F_B
         => m2s010_som_sb_MSS_0_GPIO_7_M2F, 
        SPI0_SS1_MGPIO8A_H2F_A => OPEN, SPI0_SS1_MGPIO8A_H2F_B
         => GPIO_8_M2F_c, SPI0_SS2_MGPIO9A_H2F_A => OPEN, 
        SPI0_SS2_MGPIO9A_H2F_B => OPEN, SPI0_SS3_MGPIO10A_H2F_A
         => OPEN, SPI0_SS3_MGPIO10A_H2F_B => OPEN, 
        SPI0_SS4_MGPIO19A_H2F_A => OPEN, SPI0_SS5_MGPIO20A_H2F_A
         => OPEN, SPI0_SS6_MGPIO21A_H2F_A => OPEN, 
        SPI0_SS7_MGPIO22A_H2F_A => OPEN, SPI1_CLK_OUT => 
        m2s010_som_sb_MSS_0_SPI_1_CLK_M2F, 
        SPI1_SDI_MGPIO11A_H2F_A => OPEN, SPI1_SDI_MGPIO11A_H2F_B
         => GPIO_11_M2F_c, SPI1_SDO_MGPIO12A_H2F_A => 
        SPI_1_DO_CAM_c, SPI1_SDO_MGPIO12A_H2F_B => OPEN, 
        SPI1_SS0_MGPIO13A_H2F_A => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F, 
        SPI1_SS0_MGPIO13A_H2F_B => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE, 
        SPI1_SS1_MGPIO14A_H2F_A => OPEN, SPI1_SS1_MGPIO14A_H2F_B
         => OPEN, SPI1_SS2_MGPIO15A_H2F_A => OPEN, 
        SPI1_SS2_MGPIO15A_H2F_B => OPEN, SPI1_SS3_MGPIO16A_H2F_A
         => OPEN, SPI1_SS3_MGPIO16A_H2F_B => OPEN, 
        SPI1_SS4_MGPIO17A_H2F_A => OPEN, SPI1_SS5_MGPIO18A_H2F_A
         => OPEN, SPI1_SS6_MGPIO23A_H2F_A => OPEN, 
        SPI1_SS7_MGPIO24A_H2F_A => OPEN, TCGF(9) => nc198, 
        TCGF(8) => nc147, TCGF(7) => nc67, TCGF(6) => nc152, 
        TCGF(5) => nc127, TCGF(4) => nc103, TCGF(3) => nc235, 
        TCGF(2) => nc76, TCGF(1) => nc208, TCGF(0) => nc140, 
        TRACECLK => OPEN, TRACEDATA(3) => nc86, TRACEDATA(2) => 
        nc95, TRACEDATA(1) => nc120, TRACEDATA(0) => nc165, 
        TX_CLK => OPEN, TX_ENF => MAC_MII_TX_EN_c, TX_ERRF => 
        OPEN, TXCTL_EN_RIF => OPEN, TXD_RIF(3) => nc137, 
        TXD_RIF(2) => nc64, TXD_RIF(1) => nc19, TXD_RIF(0) => 
        nc70, TXDF(7) => nc182, TXDF(6) => nc62, TXDF(5) => nc199, 
        TXDF(4) => nc80, TXDF(3) => MAC_MII_TXD_c(3), TXDF(2) => 
        MAC_MII_TXD_c(2), TXDF(1) => MAC_MII_TXD_c(1), TXDF(0)
         => MAC_MII_TXD_c(0), TXEV => OPEN, WDOGTIMEOUT => OPEN, 
        F_ARREADY_HREADYOUT1 => OPEN, F_AWREADY_HREADYOUT0 => 
        OPEN, F_BID(3) => nc130, F_BID(2) => nc98, F_BID(1) => 
        nc114, F_BID(0) => nc56, F_BRESP_HRESP0(1) => nc105, 
        F_BRESP_HRESP0(0) => nc63, F_BVALID => OPEN, 
        F_RDATA_HRDATA01(63) => nc172, F_RDATA_HRDATA01(62) => 
        nc229, F_RDATA_HRDATA01(61) => nc97, F_RDATA_HRDATA01(60)
         => nc161, F_RDATA_HRDATA01(59) => nc31, 
        F_RDATA_HRDATA01(58) => nc154, F_RDATA_HRDATA01(57) => 
        nc50, F_RDATA_HRDATA01(56) => nc239, F_RDATA_HRDATA01(55)
         => nc142, F_RDATA_HRDATA01(54) => nc94, 
        F_RDATA_HRDATA01(53) => nc197, F_RDATA_HRDATA01(52) => 
        nc122, F_RDATA_HRDATA01(51) => nc35, F_RDATA_HRDATA01(50)
         => nc4, F_RDATA_HRDATA01(49) => nc227, 
        F_RDATA_HRDATA01(48) => nc92, F_RDATA_HRDATA01(47) => 
        nc101, F_RDATA_HRDATA01(46) => nc184, 
        F_RDATA_HRDATA01(45) => nc200, F_RDATA_HRDATA01(44) => 
        nc190, F_RDATA_HRDATA01(43) => nc166, 
        F_RDATA_HRDATA01(42) => nc132, F_RDATA_HRDATA01(41) => 
        nc21, F_RDATA_HRDATA01(40) => nc237, F_RDATA_HRDATA01(39)
         => nc93, F_RDATA_HRDATA01(38) => nc69, 
        F_RDATA_HRDATA01(37) => nc206, F_RDATA_HRDATA01(36) => 
        nc174, F_RDATA_HRDATA01(35) => nc38, F_RDATA_HRDATA01(34)
         => nc113, F_RDATA_HRDATA01(33) => nc218, 
        F_RDATA_HRDATA01(32) => nc106, F_RDATA_HRDATA01(31) => 
        nc25, F_RDATA_HRDATA01(30) => nc1, F_RDATA_HRDATA01(29)
         => nc37, F_RDATA_HRDATA01(28) => nc202, 
        F_RDATA_HRDATA01(27) => nc144, F_RDATA_HRDATA01(26) => 
        nc153, F_RDATA_HRDATA01(25) => nc46, F_RDATA_HRDATA01(24)
         => nc71, F_RDATA_HRDATA01(23) => nc124, 
        F_RDATA_HRDATA01(22) => nc81, F_RDATA_HRDATA01(21) => 
        nc201, F_RDATA_HRDATA01(20) => nc168, 
        F_RDATA_HRDATA01(19) => nc34, F_RDATA_HRDATA01(18) => 
        nc28, F_RDATA_HRDATA01(17) => nc115, F_RDATA_HRDATA01(16)
         => nc192, F_RDATA_HRDATA01(15) => nc134, 
        F_RDATA_HRDATA01(14) => nc32, F_RDATA_HRDATA01(13) => 
        nc40, F_RDATA_HRDATA01(12) => nc99, F_RDATA_HRDATA01(11)
         => nc75, F_RDATA_HRDATA01(10) => nc183, 
        F_RDATA_HRDATA01(9) => nc85, F_RDATA_HRDATA01(8) => nc27, 
        F_RDATA_HRDATA01(7) => nc108, F_RDATA_HRDATA01(6) => nc16, 
        F_RDATA_HRDATA01(5) => nc155, F_RDATA_HRDATA01(4) => nc51, 
        F_RDATA_HRDATA01(3) => nc33, F_RDATA_HRDATA01(2) => nc204, 
        F_RDATA_HRDATA01(1) => nc173, F_RDATA_HRDATA01(0) => 
        nc169, F_RID(3) => nc78, F_RID(2) => nc24, F_RID(1) => 
        nc88, F_RID(0) => nc111, F_RLAST => OPEN, 
        F_RRESP_HRESP1(1) => nc55, F_RRESP_HRESP1(0) => nc10, 
        F_RVALID => OPEN, F_WREADY => OPEN, 
        MDDR_FABRIC_PRDATA(15) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(15), 
        MDDR_FABRIC_PRDATA(14) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(14), 
        MDDR_FABRIC_PRDATA(13) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(13), 
        MDDR_FABRIC_PRDATA(12) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(12), 
        MDDR_FABRIC_PRDATA(11) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(11), 
        MDDR_FABRIC_PRDATA(10) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(10), 
        MDDR_FABRIC_PRDATA(9) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(9), 
        MDDR_FABRIC_PRDATA(8) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(8), 
        MDDR_FABRIC_PRDATA(7) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(7), 
        MDDR_FABRIC_PRDATA(6) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(6), 
        MDDR_FABRIC_PRDATA(5) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(5), 
        MDDR_FABRIC_PRDATA(4) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(4), 
        MDDR_FABRIC_PRDATA(3) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(3), 
        MDDR_FABRIC_PRDATA(2) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(2), 
        MDDR_FABRIC_PRDATA(1) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(1), 
        MDDR_FABRIC_PRDATA(0) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[0]\, 
        MDDR_FABRIC_PREADY => CORECONFIGP_0_MDDR_APBmslave_PREADY, 
        MDDR_FABRIC_PSLVERR => 
        CORECONFIGP_0_MDDR_APBmslave_PSLVERR, CAN_RXBUS_F2H_SCP
         => VCC_net_1, CAN_TX_EBL_F2H_SCP => VCC_net_1, 
        CAN_TXBUS_F2H_SCP => VCC_net_1, COLF => MAC_MII_COL_c, 
        CRSF => MAC_MII_CRS_c, F2_DMAREADY(1) => VCC_net_1, 
        F2_DMAREADY(0) => VCC_net_1, F2H_INTERRUPT(15) => 
        GND_net_1, F2H_INTERRUPT(14) => GND_net_1, 
        F2H_INTERRUPT(13) => GND_net_1, F2H_INTERRUPT(12) => 
        GND_net_1, F2H_INTERRUPT(11) => GND_net_1, 
        F2H_INTERRUPT(10) => GND_net_1, F2H_INTERRUPT(9) => 
        GND_net_1, F2H_INTERRUPT(8) => GND_net_1, 
        F2H_INTERRUPT(7) => GND_net_1, F2H_INTERRUPT(6) => 
        GND_net_1, F2H_INTERRUPT(5) => GND_net_1, 
        F2H_INTERRUPT(4) => GND_net_1, F2H_INTERRUPT(3) => 
        GND_net_1, F2H_INTERRUPT(2) => GND_net_1, 
        F2H_INTERRUPT(1) => GND_net_1, F2H_INTERRUPT(0) => 
        CommsFPGA_top_0_INT, F2HCALIB => VCC_net_1, F_DMAREADY(1)
         => VCC_net_1, F_DMAREADY(0) => VCC_net_1, F_FM0_ADDR(31)
         => GND_net_1, F_FM0_ADDR(30) => GND_net_1, 
        F_FM0_ADDR(29) => GND_net_1, F_FM0_ADDR(28) => GND_net_1, 
        F_FM0_ADDR(27) => GND_net_1, F_FM0_ADDR(26) => GND_net_1, 
        F_FM0_ADDR(25) => GND_net_1, F_FM0_ADDR(24) => GND_net_1, 
        F_FM0_ADDR(23) => GND_net_1, F_FM0_ADDR(22) => GND_net_1, 
        F_FM0_ADDR(21) => GND_net_1, F_FM0_ADDR(20) => GND_net_1, 
        F_FM0_ADDR(19) => GND_net_1, F_FM0_ADDR(18) => GND_net_1, 
        F_FM0_ADDR(17) => GND_net_1, F_FM0_ADDR(16) => GND_net_1, 
        F_FM0_ADDR(15) => GND_net_1, F_FM0_ADDR(14) => GND_net_1, 
        F_FM0_ADDR(13) => GND_net_1, F_FM0_ADDR(12) => GND_net_1, 
        F_FM0_ADDR(11) => GND_net_1, F_FM0_ADDR(10) => GND_net_1, 
        F_FM0_ADDR(9) => GND_net_1, F_FM0_ADDR(8) => GND_net_1, 
        F_FM0_ADDR(7) => GND_net_1, F_FM0_ADDR(6) => GND_net_1, 
        F_FM0_ADDR(5) => GND_net_1, F_FM0_ADDR(4) => GND_net_1, 
        F_FM0_ADDR(3) => GND_net_1, F_FM0_ADDR(2) => GND_net_1, 
        F_FM0_ADDR(1) => GND_net_1, F_FM0_ADDR(0) => GND_net_1, 
        F_FM0_ENABLE => GND_net_1, F_FM0_MASTLOCK => GND_net_1, 
        F_FM0_READY => VCC_net_1, F_FM0_SEL => GND_net_1, 
        F_FM0_SIZE(1) => GND_net_1, F_FM0_SIZE(0) => GND_net_1, 
        F_FM0_TRANS1 => GND_net_1, F_FM0_WDATA(31) => GND_net_1, 
        F_FM0_WDATA(30) => GND_net_1, F_FM0_WDATA(29) => 
        GND_net_1, F_FM0_WDATA(28) => GND_net_1, F_FM0_WDATA(27)
         => GND_net_1, F_FM0_WDATA(26) => GND_net_1, 
        F_FM0_WDATA(25) => GND_net_1, F_FM0_WDATA(24) => 
        GND_net_1, F_FM0_WDATA(23) => GND_net_1, F_FM0_WDATA(22)
         => GND_net_1, F_FM0_WDATA(21) => GND_net_1, 
        F_FM0_WDATA(20) => GND_net_1, F_FM0_WDATA(19) => 
        GND_net_1, F_FM0_WDATA(18) => GND_net_1, F_FM0_WDATA(17)
         => GND_net_1, F_FM0_WDATA(16) => GND_net_1, 
        F_FM0_WDATA(15) => GND_net_1, F_FM0_WDATA(14) => 
        GND_net_1, F_FM0_WDATA(13) => GND_net_1, F_FM0_WDATA(12)
         => GND_net_1, F_FM0_WDATA(11) => GND_net_1, 
        F_FM0_WDATA(10) => GND_net_1, F_FM0_WDATA(9) => GND_net_1, 
        F_FM0_WDATA(8) => GND_net_1, F_FM0_WDATA(7) => GND_net_1, 
        F_FM0_WDATA(6) => GND_net_1, F_FM0_WDATA(5) => GND_net_1, 
        F_FM0_WDATA(4) => GND_net_1, F_FM0_WDATA(3) => GND_net_1, 
        F_FM0_WDATA(2) => GND_net_1, F_FM0_WDATA(1) => GND_net_1, 
        F_FM0_WDATA(0) => GND_net_1, F_FM0_WRITE => GND_net_1, 
        F_HM0_RDATA(31) => GND_net_1, F_HM0_RDATA(30) => 
        GND_net_1, F_HM0_RDATA(29) => GND_net_1, F_HM0_RDATA(28)
         => GND_net_1, F_HM0_RDATA(27) => GND_net_1, 
        F_HM0_RDATA(26) => GND_net_1, F_HM0_RDATA(25) => 
        GND_net_1, F_HM0_RDATA(24) => GND_net_1, F_HM0_RDATA(23)
         => GND_net_1, F_HM0_RDATA(22) => GND_net_1, 
        F_HM0_RDATA(21) => GND_net_1, F_HM0_RDATA(20) => 
        GND_net_1, F_HM0_RDATA(19) => GND_net_1, F_HM0_RDATA(18)
         => GND_net_1, F_HM0_RDATA(17) => GND_net_1, 
        F_HM0_RDATA(16) => GND_net_1, F_HM0_RDATA(15) => 
        GND_net_1, F_HM0_RDATA(14) => GND_net_1, F_HM0_RDATA(13)
         => GND_net_1, F_HM0_RDATA(12) => GND_net_1, 
        F_HM0_RDATA(11) => GND_net_1, F_HM0_RDATA(10) => 
        GND_net_1, F_HM0_RDATA(9) => GND_net_1, F_HM0_RDATA(8)
         => GND_net_1, F_HM0_RDATA(7) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(7), F_HM0_RDATA(6) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(6), F_HM0_RDATA(5) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(5), F_HM0_RDATA(4) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(4), F_HM0_RDATA(3) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(3), F_HM0_RDATA(2) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(2), F_HM0_RDATA(1) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(1), F_HM0_RDATA(0) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(0), F_HM0_READY => 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i, F_HM0_RESP => 
        GND_net_1, FAB_AVALID => VCC_net_1, FAB_HOSTDISCON => 
        VCC_net_1, FAB_IDDIG => VCC_net_1, FAB_LINESTATE(1) => 
        VCC_net_1, FAB_LINESTATE(0) => VCC_net_1, FAB_M3_RESET_N
         => VCC_net_1, FAB_PLL_LOCK => FAB_CCC_LOCK, FAB_RXACTIVE
         => VCC_net_1, FAB_RXERROR => VCC_net_1, FAB_RXVALID => 
        VCC_net_1, FAB_RXVALIDH => GND_net_1, FAB_SESSEND => 
        VCC_net_1, FAB_TXREADY => VCC_net_1, FAB_VBUSVALID => 
        VCC_net_1, FAB_VSTATUS(7) => VCC_net_1, FAB_VSTATUS(6)
         => VCC_net_1, FAB_VSTATUS(5) => VCC_net_1, 
        FAB_VSTATUS(4) => VCC_net_1, FAB_VSTATUS(3) => VCC_net_1, 
        FAB_VSTATUS(2) => VCC_net_1, FAB_VSTATUS(1) => VCC_net_1, 
        FAB_VSTATUS(0) => VCC_net_1, FAB_XDATAIN(7) => VCC_net_1, 
        FAB_XDATAIN(6) => VCC_net_1, FAB_XDATAIN(5) => VCC_net_1, 
        FAB_XDATAIN(4) => VCC_net_1, FAB_XDATAIN(3) => VCC_net_1, 
        FAB_XDATAIN(2) => VCC_net_1, FAB_XDATAIN(1) => VCC_net_1, 
        FAB_XDATAIN(0) => VCC_net_1, GTX_CLKPF => VCC_net_1, 
        I2C0_BCLK => VCC_net_1, I2C0_SCL_F2H_SCP => VCC_net_1, 
        I2C0_SDA_F2H_SCP => VCC_net_1, I2C1_BCLK => VCC_net_1, 
        I2C1_SCL_F2H_SCP => VCC_net_1, I2C1_SDA_F2H_SCP => 
        VCC_net_1, MDIF => BIBUF_0_Y, MGPIO0A_F2H_GPIN => 
        VCC_net_1, MGPIO10A_F2H_GPIN => Y_net_0(3), 
        MGPIO11A_F2H_GPIN => VCC_net_1, MGPIO11B_F2H_GPIN => 
        VCC_net_1, MGPIO12A_F2H_GPIN => VCC_net_1, 
        MGPIO13A_F2H_GPIN => VCC_net_1, MGPIO14A_F2H_GPIN => 
        VCC_net_1, MGPIO15A_F2H_GPIN => VCC_net_1, 
        MGPIO16A_F2H_GPIN => VCC_net_1, MGPIO17B_F2H_GPIN => 
        VCC_net_1, MGPIO18B_F2H_GPIN => VCC_net_1, 
        MGPIO19B_F2H_GPIN => Y_net_0(1), MGPIO1A_F2H_GPIN => 
        GPIO_1_in_0, MGPIO20B_F2H_GPIN => VCC_net_1, 
        MGPIO21B_F2H_GPIN => VCC_net_1, MGPIO22B_F2H_GPIN => 
        VCC_net_1, MGPIO24B_F2H_GPIN => VCC_net_1, 
        MGPIO25B_F2H_GPIN => VCC_net_1, MGPIO26B_F2H_GPIN => 
        VCC_net_1, MGPIO27B_F2H_GPIN => DEBOUNCE_OUT_1_c, 
        MGPIO28B_F2H_GPIN => VCC_net_1, MGPIO29B_F2H_GPIN => 
        DEBOUNCE_OUT_2_c, MGPIO2A_F2H_GPIN => Y_net_0(2), 
        MGPIO30B_F2H_GPIN => DEBOUNCE_OUT_net_0_0, 
        MGPIO31B_F2H_GPIN => VCC_net_1, MGPIO3A_F2H_GPIN => 
        VCC_net_1, MGPIO4A_F2H_GPIN => VCC_net_1, 
        MGPIO5A_F2H_GPIN => VCC_net_1, MGPIO6A_F2H_GPIN => 
        GPIO_6_Y_0, MGPIO7A_F2H_GPIN => GPIO_7_Y_0, 
        MGPIO8A_F2H_GPIN => VCC_net_1, MGPIO9A_F2H_GPIN => 
        Y_net_0(0), MMUART0_CTS_F2H_SCP => VCC_net_1, 
        MMUART0_DCD_F2H_SCP => VCC_net_1, MMUART0_DSR_F2H_SCP => 
        VCC_net_1, MMUART0_DTR_F2H_SCP => VCC_net_1, 
        MMUART0_RI_F2H_SCP => VCC_net_1, MMUART0_RTS_F2H_SCP => 
        VCC_net_1, MMUART0_RXD_F2H_SCP => MMUART_0_RXD_F2M_c, 
        MMUART0_SCK_F2H_SCP => VCC_net_1, MMUART0_TXD_F2H_SCP => 
        VCC_net_1, MMUART1_CTS_F2H_SCP => VCC_net_1, 
        MMUART1_DCD_F2H_SCP => VCC_net_1, MMUART1_DSR_F2H_SCP => 
        VCC_net_1, MMUART1_RI_F2H_SCP => VCC_net_1, 
        MMUART1_RTS_F2H_SCP => VCC_net_1, MMUART1_RXD_F2H_SCP => 
        VCC_net_1, MMUART1_SCK_F2H_SCP => VCC_net_1, 
        MMUART1_TXD_F2H_SCP => VCC_net_1, PER2_FABRIC_PRDATA(31)
         => GND_net_1, PER2_FABRIC_PRDATA(30) => GND_net_1, 
        PER2_FABRIC_PRDATA(29) => GND_net_1, 
        PER2_FABRIC_PRDATA(28) => GND_net_1, 
        PER2_FABRIC_PRDATA(27) => GND_net_1, 
        PER2_FABRIC_PRDATA(26) => GND_net_1, 
        PER2_FABRIC_PRDATA(25) => GND_net_1, 
        PER2_FABRIC_PRDATA(24) => GND_net_1, 
        PER2_FABRIC_PRDATA(23) => GND_net_1, 
        PER2_FABRIC_PRDATA(22) => GND_net_1, 
        PER2_FABRIC_PRDATA(21) => GND_net_1, 
        PER2_FABRIC_PRDATA(20) => GND_net_1, 
        PER2_FABRIC_PRDATA(19) => GND_net_1, 
        PER2_FABRIC_PRDATA(18) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(17), 
        PER2_FABRIC_PRDATA(17) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(17), 
        PER2_FABRIC_PRDATA(16) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(16), 
        PER2_FABRIC_PRDATA(15) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(15), 
        PER2_FABRIC_PRDATA(14) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(14), 
        PER2_FABRIC_PRDATA(13) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(13), 
        PER2_FABRIC_PRDATA(12) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(12), 
        PER2_FABRIC_PRDATA(11) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(11), 
        PER2_FABRIC_PRDATA(10) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(10), 
        PER2_FABRIC_PRDATA(9) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(9), 
        PER2_FABRIC_PRDATA(8) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(8), 
        PER2_FABRIC_PRDATA(7) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(7), 
        PER2_FABRIC_PRDATA(6) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(6), 
        PER2_FABRIC_PRDATA(5) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(5), 
        PER2_FABRIC_PRDATA(4) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(4), 
        PER2_FABRIC_PRDATA(3) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(3), 
        PER2_FABRIC_PRDATA(2) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(2), 
        PER2_FABRIC_PRDATA(1) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(1), 
        PER2_FABRIC_PRDATA(0) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(0), 
        PER2_FABRIC_PREADY => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY, 
        PER2_FABRIC_PSLVERR => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR, RCGF(9)
         => VCC_net_1, RCGF(8) => VCC_net_1, RCGF(7) => VCC_net_1, 
        RCGF(6) => VCC_net_1, RCGF(5) => VCC_net_1, RCGF(4) => 
        VCC_net_1, RCGF(3) => VCC_net_1, RCGF(2) => VCC_net_1, 
        RCGF(1) => VCC_net_1, RCGF(0) => VCC_net_1, RX_CLKPF => 
        MAC_MII_RX_CLK_c, RX_DVF => MAC_MII_RX_DV_c, RX_ERRF => 
        MAC_MII_RX_ER_c, RX_EV => VCC_net_1, RXDF(7) => VCC_net_1, 
        RXDF(6) => VCC_net_1, RXDF(5) => VCC_net_1, RXDF(4) => 
        VCC_net_1, RXDF(3) => MAC_MII_RXD_c(3), RXDF(2) => 
        MAC_MII_RXD_c(2), RXDF(1) => MAC_MII_RXD_c(1), RXDF(0)
         => MAC_MII_RXD_c(0), SLEEPHOLDREQ => GND_net_1, 
        SMBALERT_NI0 => VCC_net_1, SMBALERT_NI1 => VCC_net_1, 
        SMBSUS_NI0 => VCC_net_1, SMBSUS_NI1 => VCC_net_1, 
        SPI0_CLK_IN => VCC_net_1, SPI0_SDI_F2H_SCP => VCC_net_1, 
        SPI0_SDO_F2H_SCP => VCC_net_1, SPI0_SS0_F2H_SCP => 
        VCC_net_1, SPI0_SS1_F2H_SCP => VCC_net_1, 
        SPI0_SS2_F2H_SCP => VCC_net_1, SPI0_SS3_F2H_SCP => 
        VCC_net_1, SPI1_CLK_IN => CAM_SPI_1_CLK_Y_0, 
        SPI1_SDI_F2H_SCP => SPI_1_DI, SPI1_SDO_F2H_SCP => 
        VCC_net_1, SPI1_SS0_F2H_SCP => SPI_1_SS0_MX_Y, 
        SPI1_SS1_F2H_SCP => VCC_net_1, SPI1_SS2_F2H_SCP => 
        VCC_net_1, SPI1_SS3_F2H_SCP => VCC_net_1, TX_CLKPF => 
        MAC_MII_TX_CLK_c, USER_MSS_GPIO_RESET_N => VCC_net_1, 
        USER_MSS_RESET_N => VCC_net_1, XCLK_FAB => VCC_net_1, 
        CLK_BASE => m2s010_som_sb_0_CCC_71MHz, CLK_MDDR_APB => 
        \CORECONFIGP_0_APB_S_PCLK\, F_ARADDR_HADDR1(31) => 
        VCC_net_1, F_ARADDR_HADDR1(30) => VCC_net_1, 
        F_ARADDR_HADDR1(29) => VCC_net_1, F_ARADDR_HADDR1(28) => 
        VCC_net_1, F_ARADDR_HADDR1(27) => VCC_net_1, 
        F_ARADDR_HADDR1(26) => VCC_net_1, F_ARADDR_HADDR1(25) => 
        VCC_net_1, F_ARADDR_HADDR1(24) => VCC_net_1, 
        F_ARADDR_HADDR1(23) => VCC_net_1, F_ARADDR_HADDR1(22) => 
        VCC_net_1, F_ARADDR_HADDR1(21) => VCC_net_1, 
        F_ARADDR_HADDR1(20) => VCC_net_1, F_ARADDR_HADDR1(19) => 
        VCC_net_1, F_ARADDR_HADDR1(18) => VCC_net_1, 
        F_ARADDR_HADDR1(17) => VCC_net_1, F_ARADDR_HADDR1(16) => 
        VCC_net_1, F_ARADDR_HADDR1(15) => VCC_net_1, 
        F_ARADDR_HADDR1(14) => VCC_net_1, F_ARADDR_HADDR1(13) => 
        VCC_net_1, F_ARADDR_HADDR1(12) => VCC_net_1, 
        F_ARADDR_HADDR1(11) => VCC_net_1, F_ARADDR_HADDR1(10) => 
        VCC_net_1, F_ARADDR_HADDR1(9) => VCC_net_1, 
        F_ARADDR_HADDR1(8) => VCC_net_1, F_ARADDR_HADDR1(7) => 
        VCC_net_1, F_ARADDR_HADDR1(6) => VCC_net_1, 
        F_ARADDR_HADDR1(5) => VCC_net_1, F_ARADDR_HADDR1(4) => 
        VCC_net_1, F_ARADDR_HADDR1(3) => VCC_net_1, 
        F_ARADDR_HADDR1(2) => VCC_net_1, F_ARADDR_HADDR1(1) => 
        VCC_net_1, F_ARADDR_HADDR1(0) => VCC_net_1, 
        F_ARBURST_HTRANS1(1) => GND_net_1, F_ARBURST_HTRANS1(0)
         => GND_net_1, F_ARID_HSEL1(3) => GND_net_1, 
        F_ARID_HSEL1(2) => GND_net_1, F_ARID_HSEL1(1) => 
        GND_net_1, F_ARID_HSEL1(0) => GND_net_1, 
        F_ARLEN_HBURST1(3) => GND_net_1, F_ARLEN_HBURST1(2) => 
        GND_net_1, F_ARLEN_HBURST1(1) => GND_net_1, 
        F_ARLEN_HBURST1(0) => GND_net_1, F_ARLOCK_HMASTLOCK1(1)
         => GND_net_1, F_ARLOCK_HMASTLOCK1(0) => GND_net_1, 
        F_ARSIZE_HSIZE1(1) => GND_net_1, F_ARSIZE_HSIZE1(0) => 
        GND_net_1, F_ARVALID_HWRITE1 => GND_net_1, 
        F_AWADDR_HADDR0(31) => VCC_net_1, F_AWADDR_HADDR0(30) => 
        VCC_net_1, F_AWADDR_HADDR0(29) => VCC_net_1, 
        F_AWADDR_HADDR0(28) => VCC_net_1, F_AWADDR_HADDR0(27) => 
        VCC_net_1, F_AWADDR_HADDR0(26) => VCC_net_1, 
        F_AWADDR_HADDR0(25) => VCC_net_1, F_AWADDR_HADDR0(24) => 
        VCC_net_1, F_AWADDR_HADDR0(23) => VCC_net_1, 
        F_AWADDR_HADDR0(22) => VCC_net_1, F_AWADDR_HADDR0(21) => 
        VCC_net_1, F_AWADDR_HADDR0(20) => VCC_net_1, 
        F_AWADDR_HADDR0(19) => VCC_net_1, F_AWADDR_HADDR0(18) => 
        VCC_net_1, F_AWADDR_HADDR0(17) => VCC_net_1, 
        F_AWADDR_HADDR0(16) => VCC_net_1, F_AWADDR_HADDR0(15) => 
        VCC_net_1, F_AWADDR_HADDR0(14) => VCC_net_1, 
        F_AWADDR_HADDR0(13) => VCC_net_1, F_AWADDR_HADDR0(12) => 
        VCC_net_1, F_AWADDR_HADDR0(11) => VCC_net_1, 
        F_AWADDR_HADDR0(10) => VCC_net_1, F_AWADDR_HADDR0(9) => 
        VCC_net_1, F_AWADDR_HADDR0(8) => VCC_net_1, 
        F_AWADDR_HADDR0(7) => VCC_net_1, F_AWADDR_HADDR0(6) => 
        VCC_net_1, F_AWADDR_HADDR0(5) => VCC_net_1, 
        F_AWADDR_HADDR0(4) => VCC_net_1, F_AWADDR_HADDR0(3) => 
        VCC_net_1, F_AWADDR_HADDR0(2) => VCC_net_1, 
        F_AWADDR_HADDR0(1) => VCC_net_1, F_AWADDR_HADDR0(0) => 
        VCC_net_1, F_AWBURST_HTRANS0(1) => GND_net_1, 
        F_AWBURST_HTRANS0(0) => GND_net_1, F_AWID_HSEL0(3) => 
        GND_net_1, F_AWID_HSEL0(2) => GND_net_1, F_AWID_HSEL0(1)
         => GND_net_1, F_AWID_HSEL0(0) => GND_net_1, 
        F_AWLEN_HBURST0(3) => GND_net_1, F_AWLEN_HBURST0(2) => 
        GND_net_1, F_AWLEN_HBURST0(1) => GND_net_1, 
        F_AWLEN_HBURST0(0) => GND_net_1, F_AWLOCK_HMASTLOCK0(1)
         => GND_net_1, F_AWLOCK_HMASTLOCK0(0) => GND_net_1, 
        F_AWSIZE_HSIZE0(1) => GND_net_1, F_AWSIZE_HSIZE0(0) => 
        GND_net_1, F_AWVALID_HWRITE0 => GND_net_1, F_BREADY => 
        GND_net_1, F_RMW_AXI => GND_net_1, F_RREADY => GND_net_1, 
        F_WDATA_HWDATA01(63) => VCC_net_1, F_WDATA_HWDATA01(62)
         => VCC_net_1, F_WDATA_HWDATA01(61) => VCC_net_1, 
        F_WDATA_HWDATA01(60) => VCC_net_1, F_WDATA_HWDATA01(59)
         => VCC_net_1, F_WDATA_HWDATA01(58) => VCC_net_1, 
        F_WDATA_HWDATA01(57) => VCC_net_1, F_WDATA_HWDATA01(56)
         => VCC_net_1, F_WDATA_HWDATA01(55) => VCC_net_1, 
        F_WDATA_HWDATA01(54) => VCC_net_1, F_WDATA_HWDATA01(53)
         => VCC_net_1, F_WDATA_HWDATA01(52) => VCC_net_1, 
        F_WDATA_HWDATA01(51) => VCC_net_1, F_WDATA_HWDATA01(50)
         => VCC_net_1, F_WDATA_HWDATA01(49) => VCC_net_1, 
        F_WDATA_HWDATA01(48) => VCC_net_1, F_WDATA_HWDATA01(47)
         => VCC_net_1, F_WDATA_HWDATA01(46) => VCC_net_1, 
        F_WDATA_HWDATA01(45) => VCC_net_1, F_WDATA_HWDATA01(44)
         => VCC_net_1, F_WDATA_HWDATA01(43) => VCC_net_1, 
        F_WDATA_HWDATA01(42) => VCC_net_1, F_WDATA_HWDATA01(41)
         => VCC_net_1, F_WDATA_HWDATA01(40) => VCC_net_1, 
        F_WDATA_HWDATA01(39) => VCC_net_1, F_WDATA_HWDATA01(38)
         => VCC_net_1, F_WDATA_HWDATA01(37) => VCC_net_1, 
        F_WDATA_HWDATA01(36) => VCC_net_1, F_WDATA_HWDATA01(35)
         => VCC_net_1, F_WDATA_HWDATA01(34) => VCC_net_1, 
        F_WDATA_HWDATA01(33) => VCC_net_1, F_WDATA_HWDATA01(32)
         => VCC_net_1, F_WDATA_HWDATA01(31) => VCC_net_1, 
        F_WDATA_HWDATA01(30) => VCC_net_1, F_WDATA_HWDATA01(29)
         => VCC_net_1, F_WDATA_HWDATA01(28) => VCC_net_1, 
        F_WDATA_HWDATA01(27) => VCC_net_1, F_WDATA_HWDATA01(26)
         => VCC_net_1, F_WDATA_HWDATA01(25) => VCC_net_1, 
        F_WDATA_HWDATA01(24) => VCC_net_1, F_WDATA_HWDATA01(23)
         => VCC_net_1, F_WDATA_HWDATA01(22) => VCC_net_1, 
        F_WDATA_HWDATA01(21) => VCC_net_1, F_WDATA_HWDATA01(20)
         => VCC_net_1, F_WDATA_HWDATA01(19) => VCC_net_1, 
        F_WDATA_HWDATA01(18) => VCC_net_1, F_WDATA_HWDATA01(17)
         => VCC_net_1, F_WDATA_HWDATA01(16) => VCC_net_1, 
        F_WDATA_HWDATA01(15) => VCC_net_1, F_WDATA_HWDATA01(14)
         => VCC_net_1, F_WDATA_HWDATA01(13) => VCC_net_1, 
        F_WDATA_HWDATA01(12) => VCC_net_1, F_WDATA_HWDATA01(11)
         => VCC_net_1, F_WDATA_HWDATA01(10) => VCC_net_1, 
        F_WDATA_HWDATA01(9) => VCC_net_1, F_WDATA_HWDATA01(8) => 
        VCC_net_1, F_WDATA_HWDATA01(7) => VCC_net_1, 
        F_WDATA_HWDATA01(6) => VCC_net_1, F_WDATA_HWDATA01(5) => 
        VCC_net_1, F_WDATA_HWDATA01(4) => VCC_net_1, 
        F_WDATA_HWDATA01(3) => VCC_net_1, F_WDATA_HWDATA01(2) => 
        VCC_net_1, F_WDATA_HWDATA01(1) => VCC_net_1, 
        F_WDATA_HWDATA01(0) => VCC_net_1, F_WID_HREADY01(3) => 
        GND_net_1, F_WID_HREADY01(2) => GND_net_1, 
        F_WID_HREADY01(1) => GND_net_1, F_WID_HREADY01(0) => 
        GND_net_1, F_WLAST => GND_net_1, F_WSTRB(7) => GND_net_1, 
        F_WSTRB(6) => GND_net_1, F_WSTRB(5) => GND_net_1, 
        F_WSTRB(4) => GND_net_1, F_WSTRB(3) => GND_net_1, 
        F_WSTRB(2) => GND_net_1, F_WSTRB(1) => GND_net_1, 
        F_WSTRB(0) => GND_net_1, F_WVALID => GND_net_1, 
        FPGA_MDDR_ARESET_N => VCC_net_1, MDDR_FABRIC_PADDR(10)
         => CORECONFIGP_0_MDDR_APBmslave_PADDR(10), 
        MDDR_FABRIC_PADDR(9) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(9), 
        MDDR_FABRIC_PADDR(8) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(8), 
        MDDR_FABRIC_PADDR(7) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(7), 
        MDDR_FABRIC_PADDR(6) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(6), 
        MDDR_FABRIC_PADDR(5) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(5), 
        MDDR_FABRIC_PADDR(4) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(4), 
        MDDR_FABRIC_PADDR(3) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(3), 
        MDDR_FABRIC_PADDR(2) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(2), 
        MDDR_FABRIC_PENABLE => 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE, MDDR_FABRIC_PSEL
         => CORECONFIGP_0_MDDR_APBmslave_PSELx, 
        MDDR_FABRIC_PWDATA(15) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(15), 
        MDDR_FABRIC_PWDATA(14) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(14), 
        MDDR_FABRIC_PWDATA(13) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(13), 
        MDDR_FABRIC_PWDATA(12) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(12), 
        MDDR_FABRIC_PWDATA(11) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(11), 
        MDDR_FABRIC_PWDATA(10) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(10), 
        MDDR_FABRIC_PWDATA(9) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(9), 
        MDDR_FABRIC_PWDATA(8) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(8), 
        MDDR_FABRIC_PWDATA(7) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(7), 
        MDDR_FABRIC_PWDATA(6) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(6), 
        MDDR_FABRIC_PWDATA(5) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(5), 
        MDDR_FABRIC_PWDATA(4) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(4), 
        MDDR_FABRIC_PWDATA(3) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(3), 
        MDDR_FABRIC_PWDATA(2) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(2), 
        MDDR_FABRIC_PWDATA(1) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(1), 
        MDDR_FABRIC_PWDATA(0) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(0), 
        MDDR_FABRIC_PWRITE => CORECONFIGP_0_MDDR_APBmslave_PWRITE, 
        PRESET_N => \CORECONFIGP_0_APB_S_PRESET_N\, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_IN => GPIO_GPIO_3_BI_PAD_Y, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN => GPIO_GPIO_4_BI_PAD_Y, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_IN => GND_net_1, DM_IN(2)
         => GND_net_1, DM_IN(1) => MDDR_DM_RDQS_1_PAD_Y, DM_IN(0)
         => MDDR_DM_RDQS_0_PAD_Y, DRAM_DQ_IN(17) => GND_net_1, 
        DRAM_DQ_IN(16) => GND_net_1, DRAM_DQ_IN(15) => 
        MDDR_DQ_15_PAD_Y, DRAM_DQ_IN(14) => MDDR_DQ_14_PAD_Y, 
        DRAM_DQ_IN(13) => MDDR_DQ_13_PAD_Y, DRAM_DQ_IN(12) => 
        MDDR_DQ_12_PAD_Y, DRAM_DQ_IN(11) => MDDR_DQ_11_PAD_Y, 
        DRAM_DQ_IN(10) => MDDR_DQ_10_PAD_Y, DRAM_DQ_IN(9) => 
        MDDR_DQ_9_PAD_Y, DRAM_DQ_IN(8) => MDDR_DQ_8_PAD_Y, 
        DRAM_DQ_IN(7) => MDDR_DQ_7_PAD_Y, DRAM_DQ_IN(6) => 
        MDDR_DQ_6_PAD_Y, DRAM_DQ_IN(5) => MDDR_DQ_5_PAD_Y, 
        DRAM_DQ_IN(4) => MDDR_DQ_4_PAD_Y, DRAM_DQ_IN(3) => 
        MDDR_DQ_3_PAD_Y, DRAM_DQ_IN(2) => MDDR_DQ_2_PAD_Y, 
        DRAM_DQ_IN(1) => MDDR_DQ_1_PAD_Y, DRAM_DQ_IN(0) => 
        MDDR_DQ_0_PAD_Y, DRAM_DQS_IN(2) => GND_net_1, 
        DRAM_DQS_IN(1) => MDDR_DQS_1_PAD_Y, DRAM_DQS_IN(0) => 
        MDDR_DQS_0_PAD_Y, DRAM_FIFO_WE_IN(1) => GND_net_1, 
        DRAM_FIFO_WE_IN(0) => MDDR_DQS_TMATCH_0_IN_PAD_Y, 
        I2C0_SCL_USBC_DATA1_MGPIO31B_IN => GND_net_1, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_IN => GND_net_1, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_IN => I2C_1_SCL_PAD_Y, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_IN => I2C_1_SDA_PAD_Y, 
        MGPIO0B_IN => GPIO_GPIO_0_BI_PAD_Y, MGPIO10B_IN => 
        GND_net_1, MGPIO1B_IN => GND_net_1, MGPIO25A_IN => 
        GPIO_GPIO_25_BI_PAD_Y, MGPIO26A_IN => 
        GPIO_GPIO_26_BI_PAD_Y, MGPIO27A_IN => GND_net_1, 
        MGPIO28A_IN => GND_net_1, MGPIO29A_IN => GND_net_1, 
        MGPIO2B_IN => GND_net_1, MGPIO30A_IN => GND_net_1, 
        MGPIO31A_IN => GPIO_GPIO_31_BI_PAD_Y, MGPIO3B_IN => 
        GND_net_1, MGPIO4B_IN => GND_net_1, MGPIO5B_IN => 
        GND_net_1, MGPIO6B_IN => GND_net_1, MGPIO7B_IN => 
        GND_net_1, MGPIO8B_IN => GND_net_1, MGPIO9B_IN => 
        GND_net_1, MMUART0_CTS_USBC_DATA7_MGPIO19B_IN => 
        GND_net_1, MMUART0_DCD_MGPIO22B_IN => GND_net_1, 
        MMUART0_DSR_MGPIO20B_IN => GND_net_1, 
        MMUART0_DTR_USBC_DATA6_MGPIO18B_IN => GND_net_1, 
        MMUART0_RI_MGPIO21B_IN => GND_net_1, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_IN => GND_net_1, 
        MMUART0_RXD_USBC_STP_MGPIO28B_IN => GND_net_1, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_IN => GND_net_1, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_IN => GND_net_1, 
        MMUART1_CTS_MGPIO13B_IN => GND_net_1, 
        MMUART1_DCD_MGPIO16B_IN => GPIO_GPIO_16_BI_PAD_Y, 
        MMUART1_DSR_MGPIO14B_IN => GPIO_GPIO_14_BI_PAD_Y, 
        MMUART1_DTR_MGPIO12B_IN => GPIO_GPIO_12_BI_PAD_Y, 
        MMUART1_RI_MGPIO15B_IN => GPIO_GPIO_15_BI_PAD_Y, 
        MMUART1_RTS_MGPIO11B_IN => GND_net_1, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_IN => MMUART_1_RXD_PAD_Y, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_IN => GND_net_1, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_IN => GND_net_1, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN => GND_net_1, 
        RGMII_MDC_RMII_MDC_IN => GND_net_1, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN => GND_net_1, 
        RGMII_RX_CLK_IN => GND_net_1, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN => GND_net_1, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN => GND_net_1, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN => GND_net_1, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN => GND_net_1, 
        RGMII_RXD3_USBB_DATA4_IN => GND_net_1, RGMII_TX_CLK_IN
         => GND_net_1, RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN => 
        GND_net_1, RGMII_TXD0_RMII_TXD0_USBB_DIR_IN => GND_net_1, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_IN => GND_net_1, 
        RGMII_TXD2_USBB_DATA5_IN => GND_net_1, 
        RGMII_TXD3_USBB_DATA6_IN => GND_net_1, 
        SPI0_SCK_USBA_XCLK_IN => SPI_0_CLK_PAD_Y, 
        SPI0_SDI_USBA_DIR_MGPIO5A_IN => SPI_0_DI_PAD_Y, 
        SPI0_SDO_USBA_STP_MGPIO6A_IN => GND_net_1, 
        SPI0_SS0_USBA_NXT_MGPIO7A_IN => SPI_0_SS0_PAD_Y, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_IN => GND_net_1, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_IN => GND_net_1, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_IN => GND_net_1, 
        SPI0_SS4_MGPIO19A_IN => GND_net_1, SPI0_SS5_MGPIO20A_IN
         => GND_net_1, SPI0_SS6_MGPIO21A_IN => GND_net_1, 
        SPI0_SS7_MGPIO22A_IN => GND_net_1, SPI1_SCK_IN => 
        GND_net_1, SPI1_SDI_MGPIO11A_IN => GND_net_1, 
        SPI1_SDO_MGPIO12A_IN => GND_net_1, SPI1_SS0_MGPIO13A_IN
         => GND_net_1, SPI1_SS1_MGPIO14A_IN => GND_net_1, 
        SPI1_SS2_MGPIO15A_IN => GND_net_1, SPI1_SS3_MGPIO16A_IN
         => GND_net_1, SPI1_SS4_MGPIO17A_IN => 
        GPIO_GPIO_17_BI_PAD_Y, SPI1_SS5_MGPIO18A_IN => 
        GPIO_GPIO_18_BI_PAD_Y, SPI1_SS6_MGPIO23A_IN => GND_net_1, 
        SPI1_SS7_MGPIO24A_IN => GND_net_1, USBC_XCLK_IN => 
        GND_net_1, USBD_DATA0_IN => GND_net_1, USBD_DATA1_IN => 
        GND_net_1, USBD_DATA2_IN => GND_net_1, USBD_DATA3_IN => 
        GND_net_1, USBD_DATA4_IN => GND_net_1, USBD_DATA5_IN => 
        GND_net_1, USBD_DATA6_IN => GND_net_1, 
        USBD_DATA7_MGPIO23B_IN => GND_net_1, USBD_DIR_IN => 
        GND_net_1, USBD_NXT_IN => GND_net_1, USBD_STP_IN => 
        GND_net_1, USBD_XCLK_IN => GND_net_1, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT => 
        MSS_ADLIB_INST_CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT => 
        MSS_ADLIB_INST_CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT => OPEN, DRAM_ADDR(15)
         => \DRAM_ADDR_net_0[15]\, DRAM_ADDR(14) => 
        \DRAM_ADDR_net_0[14]\, DRAM_ADDR(13) => 
        \DRAM_ADDR_net_0[13]\, DRAM_ADDR(12) => 
        \DRAM_ADDR_net_0[12]\, DRAM_ADDR(11) => 
        \DRAM_ADDR_net_0[11]\, DRAM_ADDR(10) => 
        \DRAM_ADDR_net_0[10]\, DRAM_ADDR(9) => 
        \DRAM_ADDR_net_0[9]\, DRAM_ADDR(8) => 
        \DRAM_ADDR_net_0[8]\, DRAM_ADDR(7) => 
        \DRAM_ADDR_net_0[7]\, DRAM_ADDR(6) => 
        \DRAM_ADDR_net_0[6]\, DRAM_ADDR(5) => 
        \DRAM_ADDR_net_0[5]\, DRAM_ADDR(4) => 
        \DRAM_ADDR_net_0[4]\, DRAM_ADDR(3) => 
        \DRAM_ADDR_net_0[3]\, DRAM_ADDR(2) => 
        \DRAM_ADDR_net_0[2]\, DRAM_ADDR(1) => 
        \DRAM_ADDR_net_0[1]\, DRAM_ADDR(0) => 
        \DRAM_ADDR_net_0[0]\, DRAM_BA(2) => \DRAM_BA_net_0[2]\, 
        DRAM_BA(1) => \DRAM_BA_net_0[1]\, DRAM_BA(0) => 
        \DRAM_BA_net_0[0]\, DRAM_CASN => MSS_ADLIB_INST_DRAM_CASN, 
        DRAM_CKE => MSS_ADLIB_INST_DRAM_CKE, DRAM_CLK => 
        MSS_ADLIB_INST_DRAM_CLK, DRAM_CSN => 
        MSS_ADLIB_INST_DRAM_CSN, DRAM_DM_RDQS_OUT(2) => nc22, 
        DRAM_DM_RDQS_OUT(1) => \DRAM_DM_RDQS_OUT_net_0[1]\, 
        DRAM_DM_RDQS_OUT(0) => \DRAM_DM_RDQS_OUT_net_0[0]\, 
        DRAM_DQ_OUT(17) => nc210, DRAM_DQ_OUT(16) => nc185, 
        DRAM_DQ_OUT(15) => \DRAM_DQ_OUT_net_0[15]\, 
        DRAM_DQ_OUT(14) => \DRAM_DQ_OUT_net_0[14]\, 
        DRAM_DQ_OUT(13) => \DRAM_DQ_OUT_net_0[13]\, 
        DRAM_DQ_OUT(12) => \DRAM_DQ_OUT_net_0[12]\, 
        DRAM_DQ_OUT(11) => \DRAM_DQ_OUT_net_0[11]\, 
        DRAM_DQ_OUT(10) => \DRAM_DQ_OUT_net_0[10]\, 
        DRAM_DQ_OUT(9) => \DRAM_DQ_OUT_net_0[9]\, DRAM_DQ_OUT(8)
         => \DRAM_DQ_OUT_net_0[8]\, DRAM_DQ_OUT(7) => 
        \DRAM_DQ_OUT_net_0[7]\, DRAM_DQ_OUT(6) => 
        \DRAM_DQ_OUT_net_0[6]\, DRAM_DQ_OUT(5) => 
        \DRAM_DQ_OUT_net_0[5]\, DRAM_DQ_OUT(4) => 
        \DRAM_DQ_OUT_net_0[4]\, DRAM_DQ_OUT(3) => 
        \DRAM_DQ_OUT_net_0[3]\, DRAM_DQ_OUT(2) => 
        \DRAM_DQ_OUT_net_0[2]\, DRAM_DQ_OUT(1) => 
        \DRAM_DQ_OUT_net_0[1]\, DRAM_DQ_OUT(0) => 
        \DRAM_DQ_OUT_net_0[0]\, DRAM_DQS_OUT(2) => nc143, 
        DRAM_DQS_OUT(1) => \DRAM_DQS_OUT_net_0[1]\, 
        DRAM_DQS_OUT(0) => \DRAM_DQS_OUT_net_0[0]\, 
        DRAM_FIFO_WE_OUT(1) => nc77, DRAM_FIFO_WE_OUT(0) => 
        \DRAM_FIFO_WE_OUT_net_0[0]\, DRAM_ODT => 
        MSS_ADLIB_INST_DRAM_ODT, DRAM_RASN => 
        MSS_ADLIB_INST_DRAM_RASN, DRAM_RSTN => 
        MSS_ADLIB_INST_DRAM_RSTN, DRAM_WEN => 
        MSS_ADLIB_INST_DRAM_WEN, I2C0_SCL_USBC_DATA1_MGPIO31B_OUT
         => OPEN, I2C0_SDA_USBC_DATA0_MGPIO30B_OUT => OPEN, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_OUT => 
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OUT, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_OUT => 
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OUT, 
        MGPIO0B_OUT => MSS_ADLIB_INST_MGPIO0B_OUT, MGPIO10B_OUT
         => OPEN, MGPIO1B_OUT => OPEN, MGPIO25A_OUT => 
        MSS_ADLIB_INST_MGPIO25A_OUT, MGPIO26A_OUT => 
        MSS_ADLIB_INST_MGPIO26A_OUT, MGPIO27A_OUT => OPEN, 
        MGPIO28A_OUT => OPEN, MGPIO29A_OUT => OPEN, MGPIO2B_OUT
         => OPEN, MGPIO30A_OUT => OPEN, MGPIO31A_OUT => 
        MSS_ADLIB_INST_MGPIO31A_OUT, MGPIO3B_OUT => OPEN, 
        MGPIO4B_OUT => OPEN, MGPIO5B_OUT => OPEN, MGPIO6B_OUT => 
        OPEN, MGPIO7B_OUT => OPEN, MGPIO8B_OUT => OPEN, 
        MGPIO9B_OUT => OPEN, MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT
         => OPEN, MMUART0_DCD_MGPIO22B_OUT => OPEN, 
        MMUART0_DSR_MGPIO20B_OUT => OPEN, 
        MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT => OPEN, 
        MMUART0_RI_MGPIO21B_OUT => OPEN, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT => OPEN, 
        MMUART0_RXD_USBC_STP_MGPIO28B_OUT => OPEN, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OUT => OPEN, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_OUT => OPEN, 
        MMUART1_CTS_MGPIO13B_OUT => OPEN, 
        MMUART1_DCD_MGPIO16B_OUT => 
        MSS_ADLIB_INST_MMUART1_DCD_MGPIO16B_OUT, 
        MMUART1_DSR_MGPIO14B_OUT => 
        MSS_ADLIB_INST_MMUART1_DSR_MGPIO14B_OUT, 
        MMUART1_DTR_MGPIO12B_OUT => 
        MSS_ADLIB_INST_MMUART1_DTR_MGPIO12B_OUT, 
        MMUART1_RI_MGPIO15B_OUT => 
        MSS_ADLIB_INST_MMUART1_RI_MGPIO15B_OUT, 
        MMUART1_RTS_MGPIO11B_OUT => OPEN, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT => OPEN, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT => OPEN, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT => 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT => OPEN, 
        RGMII_MDC_RMII_MDC_OUT => OPEN, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT => OPEN, 
        RGMII_RX_CLK_OUT => OPEN, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT => OPEN, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT => OPEN, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT => OPEN, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT => OPEN, 
        RGMII_RXD3_USBB_DATA4_OUT => OPEN, RGMII_TX_CLK_OUT => 
        OPEN, RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT => OPEN, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT => OPEN, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_OUT => OPEN, 
        RGMII_TXD2_USBB_DATA5_OUT => OPEN, 
        RGMII_TXD3_USBB_DATA6_OUT => OPEN, SPI0_SCK_USBA_XCLK_OUT
         => MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT, 
        SPI0_SDI_USBA_DIR_MGPIO5A_OUT => OPEN, 
        SPI0_SDO_USBA_STP_MGPIO6A_OUT => 
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT, 
        SPI0_SS0_USBA_NXT_MGPIO7A_OUT => 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OUT => 
        MSS_ADLIB_INST_SPI0_SS1_USBA_DATA5_MGPIO8A_OUT, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OUT => OPEN, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OUT => OPEN, 
        SPI0_SS4_MGPIO19A_OUT => OPEN, SPI0_SS5_MGPIO20A_OUT => 
        MSS_ADLIB_INST_SPI0_SS5_MGPIO20A_OUT, 
        SPI0_SS6_MGPIO21A_OUT => OPEN, SPI0_SS7_MGPIO22A_OUT => 
        OPEN, SPI1_SCK_OUT => OPEN, SPI1_SDI_MGPIO11A_OUT => OPEN, 
        SPI1_SDO_MGPIO12A_OUT => OPEN, SPI1_SS0_MGPIO13A_OUT => 
        OPEN, SPI1_SS1_MGPIO14A_OUT => OPEN, 
        SPI1_SS2_MGPIO15A_OUT => OPEN, SPI1_SS3_MGPIO16A_OUT => 
        OPEN, SPI1_SS4_MGPIO17A_OUT => 
        MSS_ADLIB_INST_SPI1_SS4_MGPIO17A_OUT, 
        SPI1_SS5_MGPIO18A_OUT => 
        MSS_ADLIB_INST_SPI1_SS5_MGPIO18A_OUT, 
        SPI1_SS6_MGPIO23A_OUT => OPEN, SPI1_SS7_MGPIO24A_OUT => 
        OPEN, USBC_XCLK_OUT => OPEN, USBD_DATA0_OUT => OPEN, 
        USBD_DATA1_OUT => OPEN, USBD_DATA2_OUT => OPEN, 
        USBD_DATA3_OUT => OPEN, USBD_DATA4_OUT => OPEN, 
        USBD_DATA5_OUT => OPEN, USBD_DATA6_OUT => OPEN, 
        USBD_DATA7_MGPIO23B_OUT => OPEN, USBD_DIR_OUT => OPEN, 
        USBD_NXT_OUT => OPEN, USBD_STP_OUT => OPEN, USBD_XCLK_OUT
         => OPEN, CAN_RXBUS_USBA_DATA1_MGPIO3A_OE => 
        MSS_ADLIB_INST_CAN_RXBUS_USBA_DATA1_MGPIO3A_OE, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE => 
        MSS_ADLIB_INST_CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OE => OPEN, DM_OE(2) => nc6, 
        DM_OE(1) => \DM_OE_net_0[1]\, DM_OE(0) => 
        \DM_OE_net_0[0]\, DRAM_DQ_OE(17) => nc109, DRAM_DQ_OE(16)
         => nc87, DRAM_DQ_OE(15) => \DRAM_DQ_OE_net_0[15]\, 
        DRAM_DQ_OE(14) => \DRAM_DQ_OE_net_0[14]\, DRAM_DQ_OE(13)
         => \DRAM_DQ_OE_net_0[13]\, DRAM_DQ_OE(12) => 
        \DRAM_DQ_OE_net_0[12]\, DRAM_DQ_OE(11) => 
        \DRAM_DQ_OE_net_0[11]\, DRAM_DQ_OE(10) => 
        \DRAM_DQ_OE_net_0[10]\, DRAM_DQ_OE(9) => 
        \DRAM_DQ_OE_net_0[9]\, DRAM_DQ_OE(8) => 
        \DRAM_DQ_OE_net_0[8]\, DRAM_DQ_OE(7) => 
        \DRAM_DQ_OE_net_0[7]\, DRAM_DQ_OE(6) => 
        \DRAM_DQ_OE_net_0[6]\, DRAM_DQ_OE(5) => 
        \DRAM_DQ_OE_net_0[5]\, DRAM_DQ_OE(4) => 
        \DRAM_DQ_OE_net_0[4]\, DRAM_DQ_OE(3) => 
        \DRAM_DQ_OE_net_0[3]\, DRAM_DQ_OE(2) => 
        \DRAM_DQ_OE_net_0[2]\, DRAM_DQ_OE(1) => 
        \DRAM_DQ_OE_net_0[1]\, DRAM_DQ_OE(0) => 
        \DRAM_DQ_OE_net_0[0]\, DRAM_DQS_OE(2) => nc123, 
        DRAM_DQS_OE(1) => \DRAM_DQS_OE_net_0[1]\, DRAM_DQS_OE(0)
         => \DRAM_DQS_OE_net_0[0]\, 
        I2C0_SCL_USBC_DATA1_MGPIO31B_OE => OPEN, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_OE => OPEN, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_OE => 
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OE, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_OE => 
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OE, MGPIO0B_OE
         => MSS_ADLIB_INST_MGPIO0B_OE, MGPIO10B_OE => OPEN, 
        MGPIO1B_OE => OPEN, MGPIO25A_OE => 
        MSS_ADLIB_INST_MGPIO25A_OE, MGPIO26A_OE => 
        MSS_ADLIB_INST_MGPIO26A_OE, MGPIO27A_OE => OPEN, 
        MGPIO28A_OE => OPEN, MGPIO29A_OE => OPEN, MGPIO2B_OE => 
        OPEN, MGPIO30A_OE => OPEN, MGPIO31A_OE => 
        MSS_ADLIB_INST_MGPIO31A_OE, MGPIO3B_OE => OPEN, 
        MGPIO4B_OE => OPEN, MGPIO5B_OE => OPEN, MGPIO6B_OE => 
        OPEN, MGPIO7B_OE => OPEN, MGPIO8B_OE => OPEN, MGPIO9B_OE
         => OPEN, MMUART0_CTS_USBC_DATA7_MGPIO19B_OE => OPEN, 
        MMUART0_DCD_MGPIO22B_OE => OPEN, MMUART0_DSR_MGPIO20B_OE
         => OPEN, MMUART0_DTR_USBC_DATA6_MGPIO18B_OE => OPEN, 
        MMUART0_RI_MGPIO21B_OE => OPEN, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OE => OPEN, 
        MMUART0_RXD_USBC_STP_MGPIO28B_OE => OPEN, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OE => OPEN, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_OE => OPEN, 
        MMUART1_CTS_MGPIO13B_OE => OPEN, MMUART1_DCD_MGPIO16B_OE
         => MSS_ADLIB_INST_MMUART1_DCD_MGPIO16B_OE, 
        MMUART1_DSR_MGPIO14B_OE => 
        MSS_ADLIB_INST_MMUART1_DSR_MGPIO14B_OE, 
        MMUART1_DTR_MGPIO12B_OE => 
        MSS_ADLIB_INST_MMUART1_DTR_MGPIO12B_OE, 
        MMUART1_RI_MGPIO15B_OE => 
        MSS_ADLIB_INST_MMUART1_RI_MGPIO15B_OE, 
        MMUART1_RTS_MGPIO11B_OE => OPEN, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OE => OPEN, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OE => OPEN, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_OE => 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE => OPEN, 
        RGMII_MDC_RMII_MDC_OE => OPEN, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE => OPEN, 
        RGMII_RX_CLK_OE => OPEN, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE => OPEN, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE => OPEN, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE => OPEN, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE => OPEN, 
        RGMII_RXD3_USBB_DATA4_OE => OPEN, RGMII_TX_CLK_OE => OPEN, 
        RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE => OPEN, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OE => OPEN, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_OE => OPEN, 
        RGMII_TXD2_USBB_DATA5_OE => OPEN, 
        RGMII_TXD3_USBB_DATA6_OE => OPEN, SPI0_SCK_USBA_XCLK_OE
         => MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE, 
        SPI0_SDI_USBA_DIR_MGPIO5A_OE => OPEN, 
        SPI0_SDO_USBA_STP_MGPIO6A_OE => 
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE, 
        SPI0_SS0_USBA_NXT_MGPIO7A_OE => 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OE => 
        MSS_ADLIB_INST_SPI0_SS1_USBA_DATA5_MGPIO8A_OE, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OE => OPEN, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OE => OPEN, 
        SPI0_SS4_MGPIO19A_OE => OPEN, SPI0_SS5_MGPIO20A_OE => 
        OPEN, SPI0_SS6_MGPIO21A_OE => OPEN, SPI0_SS7_MGPIO22A_OE
         => OPEN, SPI1_SCK_OE => OPEN, SPI1_SDI_MGPIO11A_OE => 
        OPEN, SPI1_SDO_MGPIO12A_OE => OPEN, SPI1_SS0_MGPIO13A_OE
         => OPEN, SPI1_SS1_MGPIO14A_OE => OPEN, 
        SPI1_SS2_MGPIO15A_OE => OPEN, SPI1_SS3_MGPIO16A_OE => 
        OPEN, SPI1_SS4_MGPIO17A_OE => 
        MSS_ADLIB_INST_SPI1_SS4_MGPIO17A_OE, SPI1_SS5_MGPIO18A_OE
         => MSS_ADLIB_INST_SPI1_SS5_MGPIO18A_OE, 
        SPI1_SS6_MGPIO23A_OE => OPEN, SPI1_SS7_MGPIO24A_OE => 
        OPEN, USBC_XCLK_OE => OPEN, USBD_DATA0_OE => OPEN, 
        USBD_DATA1_OE => OPEN, USBD_DATA2_OE => OPEN, 
        USBD_DATA3_OE => OPEN, USBD_DATA4_OE => OPEN, 
        USBD_DATA5_OE => OPEN, USBD_DATA6_OE => OPEN, 
        USBD_DATA7_MGPIO23B_OE => OPEN, USBD_DIR_OE => OPEN, 
        USBD_NXT_OE => OPEN, USBD_STP_OE => OPEN, USBD_XCLK_OE
         => OPEN);
    
    MDDR_RAS_N_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => MSS_ADLIB_INST_DRAM_RASN, PAD => MDDR_RAS_N);
    
    SPI_0_CLK_PAD : BIBUF
      port map(PAD => SPI_0_CLK, D => 
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT, E => 
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE, Y => 
        SPI_0_CLK_PAD_Y);
    
    MDDR_DQ_4_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(4), D => \DRAM_DQ_OUT_net_0[4]\, E
         => \DRAM_DQ_OE_net_0[4]\, Y => MDDR_DQ_4_PAD_Y);
    
    GPIO_GPIO_18_BI_PAD : BIBUF
      port map(PAD => GPIO_18_BI, D => 
        MSS_ADLIB_INST_SPI1_SS5_MGPIO18A_OUT, E => 
        MSS_ADLIB_INST_SPI1_SS5_MGPIO18A_OE, Y => 
        GPIO_GPIO_18_BI_PAD_Y);
    
    GPIO_GPIO_16_BI_PAD : BIBUF
      port map(PAD => GPIO_16_BI, D => 
        MSS_ADLIB_INST_MMUART1_DCD_MGPIO16B_OUT, E => 
        MSS_ADLIB_INST_MMUART1_DCD_MGPIO16B_OE, Y => 
        GPIO_GPIO_16_BI_PAD_Y);
    
    MDDR_ADDR_10_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[10]\, PAD => MDDR_ADDR(10));
    
    MDDR_DQS_TMATCH_0_IN_PAD : INBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQS_TMATCH_0_IN, Y => 
        MDDR_DQS_TMATCH_0_IN_PAD_Y);
    
    MDDR_CS_N_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => MSS_ADLIB_INST_DRAM_CSN, PAD => MDDR_CS_N);
    
    MDDR_ADDR_4_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[4]\, PAD => MDDR_ADDR(4));
    
    SPI_0_SS0_PAD : BIBUF
      port map(PAD => SPI_0_SS0, D => 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT, E => 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE, Y => 
        SPI_0_SS0_PAD_Y);
    
    MDDR_DQ_7_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(7), D => \DRAM_DQ_OUT_net_0[7]\, E
         => \DRAM_DQ_OE_net_0[7]\, Y => MDDR_DQ_7_PAD_Y);
    
    MDDR_WE_N_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => MSS_ADLIB_INST_DRAM_WEN, PAD => MDDR_WE_N);
    
    MDDR_ADDR_8_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[8]\, PAD => MDDR_ADDR(8));
    
    GPIO_GPIO_3_BI_PAD : BIBUF
      port map(PAD => GPIO_3_BI, D => 
        MSS_ADLIB_INST_CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT, E => 
        MSS_ADLIB_INST_CAN_RXBUS_USBA_DATA1_MGPIO3A_OE, Y => 
        GPIO_GPIO_3_BI_PAD_Y);
    
    MDDR_ADDR_15_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[15]\, PAD => MDDR_ADDR(15));
    
    MDDR_ADDR_0_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[0]\, PAD => MDDR_ADDR(0));
    
    MDDR_ADDR_1_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[1]\, PAD => MDDR_ADDR(1));
    
    GPIO_GPIO_20_OUT_PAD : OUTBUF
      port map(D => MSS_ADLIB_INST_SPI0_SS5_MGPIO20A_OUT, PAD => 
        GPIO_20_OUT);
    
    SPI_0_SS1_PAD : TRIBUFF
      port map(D => 
        MSS_ADLIB_INST_SPI0_SS1_USBA_DATA5_MGPIO8A_OUT, E => 
        MSS_ADLIB_INST_SPI0_SS1_USBA_DATA5_MGPIO8A_OE, PAD => 
        SPI_0_SS1);
    
    FIC_2_APB_M_PCLK_inferred_clock_RNIPG5 : CLKINT
      port map(A => FIC_2_APB_M_PCLK, Y => 
        \CORECONFIGP_0_APB_S_PCLK\);
    
    MDDR_DQ_13_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(13), D => \DRAM_DQ_OUT_net_0[13]\, 
        E => \DRAM_DQ_OE_net_0[13]\, Y => MDDR_DQ_13_PAD_Y);
    
    MDDR_ADDR_3_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[3]\, PAD => MDDR_ADDR(3));
    
    MMUART_1_RXD_PAD : INBUF
      port map(PAD => MMUART_1_RXD, Y => MMUART_1_RXD_PAD_Y);
    
    MDDR_BA_0_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_BA_net_0[0]\, PAD => MDDR_BA(0));
    
    GPIO_GPIO_26_BI_PAD : BIBUF
      port map(PAD => GPIO_26_BI, D => 
        MSS_ADLIB_INST_MGPIO26A_OUT, E => 
        MSS_ADLIB_INST_MGPIO26A_OE, Y => GPIO_GPIO_26_BI_PAD_Y);
    
    MDDR_DQ_6_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(6), D => \DRAM_DQ_OUT_net_0[6]\, E
         => \DRAM_DQ_OE_net_0[6]\, Y => MDDR_DQ_6_PAD_Y);
    
    MDDR_CLK_PAD : OUTBUF_DIFF
      generic map(IOSTD => "LPDDRI")

      port map(D => MSS_ADLIB_INST_DRAM_CLK, PADP => MDDR_CLK, 
        PADN => MDDR_CLK_N);
    
    MDDR_DQ_14_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(14), D => \DRAM_DQ_OUT_net_0[14]\, 
        E => \DRAM_DQ_OE_net_0[14]\, Y => MDDR_DQ_14_PAD_Y);
    
    GPIO_GPIO_15_BI_PAD : BIBUF
      port map(PAD => GPIO_15_BI, D => 
        MSS_ADLIB_INST_MMUART1_RI_MGPIO15B_OUT, E => 
        MSS_ADLIB_INST_MMUART1_RI_MGPIO15B_OE, Y => 
        GPIO_GPIO_15_BI_PAD_Y);
    
    MDDR_DQS_TMATCH_0_OUT_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_FIFO_WE_OUT_net_0[0]\, PAD => 
        MDDR_DQS_TMATCH_0_OUT);
    
    MDDR_BA_1_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_BA_net_0[1]\, PAD => MDDR_BA(1));
    
    MDDR_DQ_5_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(5), D => \DRAM_DQ_OUT_net_0[5]\, E
         => \DRAM_DQ_OE_net_0[5]\, Y => MDDR_DQ_5_PAD_Y);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreResetP is

    port( CORECONFIGP_0_CONFIG2_DONE              : in    std_logic;
          CORECONFIGP_0_CONFIG1_DONE              : in    std_logic;
          CORECONFIGP_0_APB_S_PRESET_N            : in    std_logic;
          m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F : in    std_logic;
          m2s010_som_sb_0_POWER_ON_RESET_N        : in    std_logic;
          INIT_DONE                               : out   std_logic;
          FABOSC_0_RCOSC_25_50MHZ_O2F             : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz               : in    std_logic
        );

end CoreResetP;

architecture DEF_ARCH of CoreResetP is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \sm0_areset_n_rcosc\, sm0_areset_n_rcosc_0, 
        \sm0_areset_n_clk_base\, sm0_areset_n_clk_base_0, 
        \count_ddr[0]_net_1\, \count_ddr_s[0]\, \mss_ready_state\, 
        VCC_net_1, \POWER_ON_RESET_N_clk_base\, 
        \RESET_N_M2F_clk_base\, GND_net_1, \ddr_settled\, 
        \un14_count_ddr\, \count_ddr_enable\, 
        next_count_ddr_enable_0_sqmuxa, 
        \un1_next_ddr_ready_0_sqmuxa\, \mss_ready_select\, 
        \un6_fic_2_apb_m_preset_n_clk_base\, \sm0_state[0]_net_1\, 
        \sm0_state[6]_net_1\, \sm0_state[5]_net_1\, 
        \sm0_state[4]_net_1\, \sm0_state_ns[2]_net_1\, 
        \sm0_state[3]_net_1\, \sm0_state_ns[3]_net_1\, 
        \sm0_state[2]_net_1\, \sm0_state_ns[4]_net_1\, 
        \sm0_state[1]_net_1\, \sm0_state_ns[5]_net_1\, 
        \sm0_state_ns_a3[6]_net_1\, \MSS_HPMS_READY_int\, 
        \MSS_HPMS_READY_int_3\, sm0_areset_n_rcosc_q1, 
        sm0_areset_n_i_i, \release_sdif0_core_q1\, 
        \release_sdif0_core\, \POWER_ON_RESET_N_q1\, 
        \RESET_N_M2F_q1\, \FIC_2_APB_M_PRESET_N_q1\, 
        \sdif3_spll_lock_q1\, \count_ddr_enable_rcosc\, 
        \count_ddr_enable_q1\, \ddr_settled_clk_base\, 
        \ddr_settled_q1\, \release_sdif0_core_clk_base\, 
        \FIC_2_APB_M_PRESET_N_clk_base\, \sm0_areset_n_q1\, 
        \CONFIG1_DONE_clk_base\, \CONFIG1_DONE_q1\, 
        \CONFIG2_DONE_clk_base\, \CONFIG2_DONE_q1\, 
        \sdif3_spll_lock_q2\, \count_ddr[1]_net_1\, 
        \count_ddr_s[1]\, \count_ddr[2]_net_1\, \count_ddr_s[2]\, 
        \count_ddr[3]_net_1\, \count_ddr_s[3]\, 
        \count_ddr[4]_net_1\, \count_ddr_s[4]\, 
        \count_ddr[5]_net_1\, \count_ddr_s[5]\, 
        \count_ddr[6]_net_1\, \count_ddr_s[6]\, 
        \count_ddr[7]_net_1\, \count_ddr_s[7]\, 
        \count_ddr[8]_net_1\, \count_ddr_s[8]\, 
        \count_ddr[9]_net_1\, \count_ddr_s[9]\, 
        \count_ddr[10]_net_1\, \count_ddr_s[10]\, 
        \count_ddr[11]_net_1\, \count_ddr_s[11]\, 
        \count_ddr[12]_net_1\, \count_ddr_s[12]\, 
        \count_ddr[13]_net_1\, \count_ddr_s[13]_net_1\, 
        count_ddr_s_373_FCO, \count_ddr_cry[1]_net_1\, 
        \count_ddr_cry[2]_net_1\, \count_ddr_cry[3]_net_1\, 
        \count_ddr_cry[4]_net_1\, \count_ddr_cry[5]_net_1\, 
        \count_ddr_cry[6]_net_1\, \count_ddr_cry[7]_net_1\, 
        \count_ddr_cry[8]_net_1\, \count_ddr_cry[9]_net_1\, 
        \count_ddr_cry[10]_net_1\, \count_ddr_cry[11]_net_1\, 
        \count_ddr_cry[12]_net_1\, \un14_count_ddr_6\, 
        \un8_ddr_settled_clk_base\, \un14_count_ddr_9\, 
        \un14_count_ddr_8\, \un14_count_ddr_7\ : std_logic;

begin 


    un14_count_ddr : CFG4
      generic map(INIT => x"8000")

      port map(A => \un14_count_ddr_7\, B => \un14_count_ddr_6\, 
        C => \un14_count_ddr_8\, D => \un14_count_ddr_9\, Y => 
        \un14_count_ddr\);
    
    \sm0_state_ns[4]\ : CFG4
      generic map(INIT => x"FF70")

      port map(A => \release_sdif0_core_clk_base\, B => 
        \ddr_settled_clk_base\, C => \sm0_state[2]_net_1\, D => 
        next_count_ddr_enable_0_sqmuxa, Y => 
        \sm0_state_ns[4]_net_1\);
    
    sm0_areset_n_rcosc : SLE
      port map(D => sm0_areset_n_rcosc_q1, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => VCC_net_1, ALn => 
        sm0_areset_n_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        sm0_areset_n_rcosc_0);
    
    \count_ddr[3]\ : SLE
      port map(D => \count_ddr_s[3]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[3]_net_1\);
    
    sm0_areset_n_q1 : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => sm0_areset_n_i_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sm0_areset_n_q1\);
    
    MSS_HPMS_READY_int_RNINOKG : CFG2
      generic map(INIT => x"8")

      port map(A => \MSS_HPMS_READY_int\, B => 
        m2s010_som_sb_0_POWER_ON_RESET_N, Y => sm0_areset_n_i_i);
    
    count_ddr_s_373 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => count_ddr_s_373_FCO);
    
    count_ddr_enable_q1 : SLE
      port map(D => \count_ddr_enable\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => VCC_net_1, ALn => 
        \sm0_areset_n_rcosc\, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \count_ddr_enable_q1\);
    
    \sm0_state[6]\ : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => \sm0_areset_n_clk_base\, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sm0_state[6]_net_1\);
    
    \sm0_state[2]\ : SLE
      port map(D => \sm0_state_ns[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sm0_state[2]_net_1\);
    
    FIC_2_APB_M_PRESET_N_clk_base : SLE
      port map(D => \FIC_2_APB_M_PRESET_N_q1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \FIC_2_APB_M_PRESET_N_clk_base\);
    
    \count_ddr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[3]_net_1\, S => \count_ddr_s[4]\, Y => 
        OPEN, FCO => \count_ddr_cry[4]_net_1\);
    
    un8_ddr_settled_clk_base : CFG2
      generic map(INIT => x"8")

      port map(A => \ddr_settled_clk_base\, B => 
        \release_sdif0_core_clk_base\, Y => 
        \un8_ddr_settled_clk_base\);
    
    INIT_DONE_int : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \sm0_state[0]_net_1\, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        INIT_DONE);
    
    \count_ddr[9]\ : SLE
      port map(D => \count_ddr_s[9]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[9]_net_1\);
    
    MSS_HPMS_READY_int : SLE
      port map(D => \MSS_HPMS_READY_int_3\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \POWER_ON_RESET_N_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \MSS_HPMS_READY_int\);
    
    count_ddr_enable_rcosc : SLE
      port map(D => \count_ddr_enable_q1\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => VCC_net_1, ALn => 
        \sm0_areset_n_rcosc\, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \count_ddr_enable_rcosc\);
    
    sm0_areset_n_clk_base_RNIEFM9 : CLKINT
      port map(A => sm0_areset_n_clk_base_0, Y => 
        \sm0_areset_n_clk_base\);
    
    \count_ddr[7]\ : SLE
      port map(D => \count_ddr_s[7]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[7]_net_1\);
    
    \sm0_state_ns_a3[6]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \CONFIG2_DONE_clk_base\, B => 
        \sm0_state[1]_net_1\, Y => \sm0_state_ns_a3[6]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sm0_state[4]\ : SLE
      port map(D => \sm0_state_ns[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sm0_state[4]_net_1\);
    
    MSS_HPMS_READY_int_3 : CFG3
      generic map(INIT => x"E0")

      port map(A => \RESET_N_M2F_clk_base\, B => 
        \mss_ready_select\, C => \FIC_2_APB_M_PRESET_N_clk_base\, 
        Y => \MSS_HPMS_READY_int_3\);
    
    count_ddr_enable : SLE
      port map(D => next_count_ddr_enable_0_sqmuxa, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        \un1_next_ddr_ready_0_sqmuxa\, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \count_ddr_enable\);
    
    \count_ddr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[9]_net_1\, S => \count_ddr_s[10]\, Y => 
        OPEN, FCO => \count_ddr_cry[10]_net_1\);
    
    \sm0_state[5]\ : SLE
      port map(D => \sm0_state[6]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sm0_state[5]_net_1\);
    
    \count_ddr_cry[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[10]_net_1\, S => \count_ddr_s[11]\, Y => 
        OPEN, FCO => \count_ddr_cry[11]_net_1\);
    
    \count_ddr[8]\ : SLE
      port map(D => \count_ddr_s[8]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[8]_net_1\);
    
    \sm0_state_ns[2]\ : CFG3
      generic map(INIT => x"AE")

      port map(A => \sm0_state[5]_net_1\, B => 
        \sm0_state[4]_net_1\, C => \CONFIG1_DONE_clk_base\, Y => 
        \sm0_state_ns[2]_net_1\);
    
    sm0_areset_n_clk_base : SLE
      port map(D => \sm0_areset_n_q1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        sm0_areset_n_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        sm0_areset_n_clk_base_0);
    
    \count_ddr_cry[12]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[12]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[11]_net_1\, S => \count_ddr_s[12]\, Y => 
        OPEN, FCO => \count_ddr_cry[12]_net_1\);
    
    mss_ready_state : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \RESET_N_M2F_clk_base\, ALn => 
        \POWER_ON_RESET_N_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mss_ready_state\);
    
    \sm0_state[1]\ : SLE
      port map(D => \sm0_state_ns[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sm0_state[1]_net_1\);
    
    next_count_ddr_enable_0_sqmuxa_0_a3 : CFG2
      generic map(INIT => x"8")

      port map(A => \sdif3_spll_lock_q2\, B => 
        \sm0_state[3]_net_1\, Y => next_count_ddr_enable_0_sqmuxa);
    
    ddr_settled_clk_base : SLE
      port map(D => \ddr_settled_q1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ddr_settled_clk_base\);
    
    FIC_2_APB_M_PRESET_N_q1 : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \FIC_2_APB_M_PRESET_N_q1\);
    
    un14_count_ddr_7 : CFG4
      generic map(INIT => x"8000")

      port map(A => \count_ddr[10]_net_1\, B => 
        \count_ddr[9]_net_1\, C => \count_ddr[8]_net_1\, D => 
        \count_ddr[4]_net_1\, Y => \un14_count_ddr_7\);
    
    \count_ddr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[7]_net_1\, S => \count_ddr_s[8]\, Y => 
        OPEN, FCO => \count_ddr_cry[8]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \count_ddr_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \count_ddr[0]_net_1\, Y => \count_ddr_s[0]\);
    
    POWER_ON_RESET_N_clk_base : SLE
      port map(D => \POWER_ON_RESET_N_q1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        m2s010_som_sb_0_POWER_ON_RESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \POWER_ON_RESET_N_clk_base\);
    
    \count_ddr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => count_ddr_s_373_FCO, S
         => \count_ddr_s[1]\, Y => OPEN, FCO => 
        \count_ddr_cry[1]_net_1\);
    
    RESET_N_M2F_q1 : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => 
        m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \RESET_N_M2F_q1\);
    
    release_sdif0_core_q1 : SLE
      port map(D => \release_sdif0_core\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \release_sdif0_core_q1\);
    
    \count_ddr[10]\ : SLE
      port map(D => \count_ddr_s[10]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[10]_net_1\);
    
    \count_ddr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[5]_net_1\, S => \count_ddr_s[6]\, Y => 
        OPEN, FCO => \count_ddr_cry[6]_net_1\);
    
    \count_ddr_s[13]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[13]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[12]_net_1\, S => \count_ddr_s[13]_net_1\, 
        Y => OPEN, FCO => OPEN);
    
    \count_ddr[5]\ : SLE
      port map(D => \count_ddr_s[5]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[5]_net_1\);
    
    \count_ddr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[2]_net_1\, S => \count_ddr_s[3]\, Y => 
        OPEN, FCO => \count_ddr_cry[3]_net_1\);
    
    \count_ddr[2]\ : SLE
      port map(D => \count_ddr_s[2]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[2]_net_1\);
    
    sdif0_areset_n_rcosc_q1 : SLE
      port map(D => VCC_net_1, CLK => FABOSC_0_RCOSC_25_50MHZ_O2F, 
        EN => VCC_net_1, ALn => sm0_areset_n_i_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => sm0_areset_n_rcosc_q1);
    
    \count_ddr[1]\ : SLE
      port map(D => \count_ddr_s[1]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[1]_net_1\);
    
    \sm0_state[0]\ : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \sm0_state_ns_a3[6]_net_1\, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sm0_state[0]_net_1\);
    
    un14_count_ddr_8 : CFG4
      generic map(INIT => x"0001")

      port map(A => \count_ddr[7]_net_1\, B => 
        \count_ddr[6]_net_1\, C => \count_ddr[5]_net_1\, D => 
        \count_ddr[3]_net_1\, Y => \un14_count_ddr_8\);
    
    \count_ddr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[1]_net_1\, S => \count_ddr_s[2]\, Y => 
        OPEN, FCO => \count_ddr_cry[2]_net_1\);
    
    \count_ddr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[4]_net_1\, S => \count_ddr_s[5]\, Y => 
        OPEN, FCO => \count_ddr_cry[5]_net_1\);
    
    ddr_settled_q1 : SLE
      port map(D => \ddr_settled\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ddr_settled_q1\);
    
    \count_ddr[11]\ : SLE
      port map(D => \count_ddr_s[11]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[11]_net_1\);
    
    un14_count_ddr_9 : CFG4
      generic map(INIT => x"0001")

      port map(A => \count_ddr[12]_net_1\, B => 
        \count_ddr[11]_net_1\, C => \count_ddr[2]_net_1\, D => 
        \count_ddr[1]_net_1\, Y => \un14_count_ddr_9\);
    
    \sm0_state[3]\ : SLE
      port map(D => \sm0_state_ns[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sm0_state[3]_net_1\);
    
    \sm0_state_ns[3]\ : CFG4
      generic map(INIT => x"F222")

      port map(A => \sm0_state[3]_net_1\, B => 
        \sdif3_spll_lock_q2\, C => \sm0_state[4]_net_1\, D => 
        \CONFIG1_DONE_clk_base\, Y => \sm0_state_ns[3]_net_1\);
    
    \count_ddr[0]\ : SLE
      port map(D => \count_ddr_s[0]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[0]_net_1\);
    
    CONFIG2_DONE_q1 : SLE
      port map(D => CORECONFIGP_0_CONFIG2_DONE, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \CONFIG2_DONE_q1\);
    
    CONFIG2_DONE_clk_base : SLE
      port map(D => \CONFIG2_DONE_q1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \CONFIG2_DONE_clk_base\);
    
    CONFIG1_DONE_clk_base : SLE
      port map(D => \CONFIG1_DONE_q1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \CONFIG1_DONE_clk_base\);
    
    sm0_areset_n_rcosc_RNIKFSA : CLKINT
      port map(A => sm0_areset_n_rcosc_0, Y => 
        \sm0_areset_n_rcosc\);
    
    mss_ready_select : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \un6_fic_2_apb_m_preset_n_clk_base\, ALn => 
        \POWER_ON_RESET_N_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mss_ready_select\);
    
    un6_fic_2_apb_m_preset_n_clk_base : CFG2
      generic map(INIT => x"8")

      port map(A => \FIC_2_APB_M_PRESET_N_clk_base\, B => 
        \mss_ready_state\, Y => 
        \un6_fic_2_apb_m_preset_n_clk_base\);
    
    \count_ddr[4]\ : SLE
      port map(D => \count_ddr_s[4]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[4]_net_1\);
    
    \count_ddr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[6]_net_1\, S => \count_ddr_s[7]\, Y => 
        OPEN, FCO => \count_ddr_cry[7]_net_1\);
    
    release_sdif0_core : SLE
      port map(D => VCC_net_1, CLK => FABOSC_0_RCOSC_25_50MHZ_O2F, 
        EN => VCC_net_1, ALn => \sm0_areset_n_rcosc\, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \release_sdif0_core\);
    
    POWER_ON_RESET_N_q1 : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => m2s010_som_sb_0_POWER_ON_RESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \POWER_ON_RESET_N_q1\);
    
    \count_ddr[12]\ : SLE
      port map(D => \count_ddr_s[12]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[12]_net_1\);
    
    ddr_settled : SLE
      port map(D => VCC_net_1, CLK => FABOSC_0_RCOSC_25_50MHZ_O2F, 
        EN => \un14_count_ddr\, ALn => \sm0_areset_n_rcosc\, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \ddr_settled\);
    
    \count_ddr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[8]_net_1\, S => \count_ddr_s[9]\, Y => 
        OPEN, FCO => \count_ddr_cry[9]_net_1\);
    
    \count_ddr[6]\ : SLE
      port map(D => \count_ddr_s[6]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[6]_net_1\);
    
    CONFIG1_DONE_q1 : SLE
      port map(D => CORECONFIGP_0_CONFIG1_DONE, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \CONFIG1_DONE_q1\);
    
    un14_count_ddr_6 : CFG2
      generic map(INIT => x"4")

      port map(A => \count_ddr[0]_net_1\, B => 
        \count_ddr[13]_net_1\, Y => \un14_count_ddr_6\);
    
    sdif3_spll_lock_q1 : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => \sm0_areset_n_clk_base\, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sdif3_spll_lock_q1\);
    
    release_sdif0_core_clk_base : SLE
      port map(D => \release_sdif0_core_q1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \release_sdif0_core_clk_base\);
    
    sdif3_spll_lock_q2 : SLE
      port map(D => \sdif3_spll_lock_q1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sdif3_spll_lock_q2\);
    
    RESET_N_M2F_clk_base : SLE
      port map(D => \RESET_N_M2F_q1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \RESET_N_M2F_clk_base\);
    
    un1_next_ddr_ready_0_sqmuxa : CFG4
      generic map(INIT => x"F888")

      port map(A => \sdif3_spll_lock_q2\, B => 
        \sm0_state[3]_net_1\, C => \ddr_settled_clk_base\, D => 
        \sm0_state[2]_net_1\, Y => \un1_next_ddr_ready_0_sqmuxa\);
    
    \count_ddr[13]\ : SLE
      port map(D => \count_ddr_s[13]_net_1\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[13]_net_1\);
    
    \sm0_state_ns[5]\ : CFG4
      generic map(INIT => x"F444")

      port map(A => \CONFIG2_DONE_clk_base\, B => 
        \sm0_state[1]_net_1\, C => \un8_ddr_settled_clk_base\, D
         => \sm0_state[2]_net_1\, Y => \sm0_state_ns[5]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb_GPIO_6_IO is

    port( GPIO_6_PAD_0                      : inout std_logic := 'Z';
          GPIO_6_Y_0                        : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_6_M2F_OE : in    std_logic;
          m2s010_som_sb_MSS_0_GPIO_6_M2F    : in    std_logic
        );

end m2s010_som_sb_GPIO_6_IO;

architecture DEF_ARCH of m2s010_som_sb_GPIO_6_IO is 

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    U0_0 : BIBUF
      generic map(IOSTD => "LVCMOS33")

      port map(PAD => GPIO_6_PAD_0, D => 
        m2s010_som_sb_MSS_0_GPIO_6_M2F, E => 
        m2s010_som_sb_MSS_0_GPIO_6_M2F_OE, Y => GPIO_6_Y_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreConfigP is

    port( CORECONFIGP_0_MDDR_APBmslave_PRDATA              : in    std_logic_vector(15 downto 1);
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA  : out   std_logic_vector(17 downto 0);
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR   : in    std_logic_vector(15 downto 2);
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA  : in    std_logic_vector(16 downto 0);
          CORECONFIGP_0_MDDR_APBmslave_PADDR               : out   std_logic_vector(10 downto 2);
          CORECONFIGP_0_MDDR_APBmslave_PWDATA              : out   std_logic_vector(15 downto 0);
          CORECONFIGP_0_MDDR_APBmslave_PRDATA_reto_0       : in    std_logic;
          state_0                                          : out   std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PSLVERR             : in    std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx   : in    std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE : in    std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PREADY              : in    std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PSELx               : out   std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PENABLE             : out   std_logic;
          INIT_DONE                                        : in    std_logic;
          CORECONFIGP_0_APB_S_PCLK_i                       : in    std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE  : in    std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PWRITE              : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY  : out   std_logic;
          CORECONFIGP_0_CONFIG2_DONE                       : out   std_logic;
          CORECONFIGP_0_CONFIG1_DONE                       : out   std_logic;
          CORECONFIGP_0_APB_S_PCLK                         : in    std_logic;
          CORECONFIGP_0_APB_S_PRESET_N                     : in    std_logic
        );

end CoreConfigP;

architecture DEF_ARCH of CoreConfigP is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \state_d[2]\, GND_net_1, \paddr[12]_net_1\, 
        \paddr_60\, \paddr[13]_net_1\, \paddr_61\, 
        \paddr[15]_net_1\, \paddr_63\, 
        \CORECONFIGP_0_CONFIG1_DONE\, \un8_int_psel\, 
        \CORECONFIGP_0_CONFIG2_DONE\, \prdata[13]\, \state_0\, 
        \prdata[14]\, \prdata[15]\, \prdata[16]\, 
        \prdata_0_iv_1[16]\, \soft_reset_reg[15]_net_1\, 
        \un17_int_psel\, \soft_reset_reg[16]_net_1\, \prdata[1]\, 
        \prdata[2]\, \prdata[3]\, \prdata[4]\, \prdata[5]\, 
        \prdata[6]\, \prdata[7]\, \prdata[8]\, \prdata[9]\, 
        \prdata[10]\, \prdata[11]\, \prdata[12]\, 
        \soft_reset_reg[0]_net_1\, \soft_reset_reg[1]_net_1\, 
        \soft_reset_reg[2]_net_1\, \soft_reset_reg[3]_net_1\, 
        \soft_reset_reg[4]_net_1\, \soft_reset_reg[5]_net_1\, 
        \soft_reset_reg[6]_net_1\, \soft_reset_reg[7]_net_1\, 
        \soft_reset_reg[8]_net_1\, \soft_reset_reg[9]_net_1\, 
        \soft_reset_reg[10]_net_1\, \soft_reset_reg[11]_net_1\, 
        \soft_reset_reg[12]_net_1\, \soft_reset_reg[13]_net_1\, 
        \soft_reset_reg[14]_net_1\, 
        un1_next_FIC_2_APB_M_PREADY_0_sqmuxa, pslverr, 
        \state[0]_net_1\, \state_ns[0]\, \state_ns[1]\, \psel\, 
        \state_d_i[2]\, \INIT_DONE_q2\, \INIT_DONE_q1\, 
        \MDDR_PENABLE_0_1\, \prdata_0_iv_1_reto[0]\, 
        \prdata_0_iv_1[0]_net_1\, \soft_reset_reg_m_reto[0]\, 
        \soft_reset_reg_m[0]\, 
        CORECONFIGP_0_MDDR_APBmslave_PSELx_reto, 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, 
        \un1_fic_2_apb_m_psel\, pready, \prdata_0_iv_1_N_3L3\, 
        \prdata_0_iv_1_1[0]\, \prdata_0_iv_1_N_4L6\, N_486, 
        \control_reg_1_m_1[0]\, \paddr_RNI09N31[12]_net_1\, 
        \int_prdata_3_sqmuxa_0\, \un6_int_psel_1\, N_471, N_468, 
        soft_N_6_0, \FIC_2_APB_M_PRDATA_0_ret_1_RNO_0\, 
        int_prdata_4_sqmuxa_out_0, \soft_reset_reg_m_0[10]\, 
        \soft_reset_reg_m_0[4]\, \soft_reset_reg_m_0[6]\, 
        \soft_reset_reg_m_0[11]\, \int_prdata_3_sqmuxa\, 
        \soft_reset_reg_m[1]\, \soft_reset_reg_m[9]\, 
        \soft_reset_reg_m[7]\, \soft_reset_reg_m[5]\, 
        \soft_reset_reg_m[3]\, \soft_reset_reg_m[13]\, 
        \soft_reset_reg_m[2]\, \soft_reset_reg_m[12]\, 
        \soft_reset_reg_m[14]\, \soft_reset_reg_m[15]\, 
        \soft_reset_reg_m[8]\, \control_reg_1_m[1]\ : std_logic;

begin 

    state_0 <= \state_0\;
    CORECONFIGP_0_MDDR_APBmslave_PSELx <= 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\;
    CORECONFIGP_0_CONFIG2_DONE <= \CORECONFIGP_0_CONFIG2_DONE\;
    CORECONFIGP_0_CONFIG1_DONE <= \CORECONFIGP_0_CONFIG1_DONE\;

    \state[0]\ : SLE
      port map(D => \state_ns[0]\, CLK => 
        CORECONFIGP_0_APB_S_PCLK, EN => VCC_net_1, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \state[0]_net_1\);
    
    psel_RNI30HQ1 : CFG3
      generic map(INIT => x"DF")

      port map(A => \paddr_RNI09N31[12]_net_1\, B => 
        CORECONFIGP_0_MDDR_APBmslave_PREADY, C => \psel\, Y => 
        pready);
    
    \FIC_2_APB_M_PRDATA_0[9]\ : SLE
      port map(D => \prdata[9]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state_0\, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(9));
    
    FIC_2_APB_M_PSLVERR_0_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => CORECONFIGP_0_MDDR_APBmslave_PSLVERR, B => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, Y => pslverr);
    
    \FIC_2_APB_M_PRDATA_0[5]\ : SLE
      port map(D => \prdata[5]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state_0\, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(5));
    
    \paddr[5]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(5), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(5));
    
    \FIC_2_APB_M_PRDATA_0[4]\ : SLE
      port map(D => \prdata[4]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state_0\, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(4));
    
    \paddr[2]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(2));
    
    \FIC_2_APB_M_PRDATA_0[13]\ : SLE
      port map(D => \prdata[13]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state_0\, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(13));
    
    FIC_2_APB_M_PRDATA_0_ret_1_RNO_0 : CFG2
      generic map(INIT => x"4")

      port map(A => \paddr[15]_net_1\, B => \paddr[13]_net_1\, Y
         => \FIC_2_APB_M_PRDATA_0_ret_1_RNO_0\);
    
    \prdata_0_iv_RNO[15]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \control_reg_1_m_1[0]\, B => N_486, C => 
        N_471, D => \soft_reset_reg[15]_net_1\, Y => 
        \soft_reset_reg_m[15]\);
    
    FIC_2_APB_M_PREADY_0 : SLE
      port map(D => \state_0\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => un1_next_FIC_2_APB_M_PREADY_0_sqmuxa, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY);
    
    \control_reg_1[1]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(1), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un8_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \CORECONFIGP_0_CONFIG2_DONE\);
    
    \pwdata[8]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(8), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(8));
    
    \prdata_0_iv[11]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \soft_reset_reg_m_0[11]\, B => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(11), C => 
        int_prdata_4_sqmuxa_out_0, D => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, Y => \prdata[11]\);
    
    int_prdata_4_sqmuxa_s_0 : CFG4
      generic map(INIT => x"A8AA")

      port map(A => N_471, B => \paddr[13]_net_1\, C => 
        \paddr[15]_net_1\, D => \psel\, Y => 
        int_prdata_4_sqmuxa_out_0);
    
    FIC_2_APB_M_PRDATA_0_ret_2 : SLE
      port map(D => \CORECONFIGP_0_MDDR_APBmslave_PSELx\, CLK => 
        CORECONFIGP_0_APB_S_PCLK, EN => \state_0\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PSELx_reto);
    
    paddr_63 : CFG3
      generic map(INIT => x"D8")

      port map(A => \state_d[2]\, B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(15), C => 
        \paddr[15]_net_1\, Y => \paddr_63\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \FIC_2_APB_M_PRDATA_0[8]\ : SLE
      port map(D => \prdata[8]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state_0\, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(8));
    
    \prdata_0_iv_RNO[3]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \control_reg_1_m_1[0]\, B => N_486, C => 
        N_471, D => \soft_reset_reg[3]_net_1\, Y => 
        \soft_reset_reg_m[3]\);
    
    \pwdata[10]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(10), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(10));
    
    \pwdata[4]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(4), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(4));
    
    \soft_reset_reg[6]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(6), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[6]_net_1\);
    
    \FIC_2_APB_M_PRDATA_0[6]\ : SLE
      port map(D => \prdata[6]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state_0\, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(6));
    
    \pwdata[7]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(7), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(7));
    
    \paddr[7]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(7), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(7));
    
    \pwdata[0]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(0), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(0));
    
    \FIC_2_APB_M_PRDATA_0[16]\ : SLE
      port map(D => \prdata[16]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state_0\, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(16));
    
    \pwdata[13]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(13), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(13));
    
    \soft_reset_reg[3]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(3), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[3]_net_1\);
    
    FIC_2_APB_M_PRDATA_0_ret_1 : SLE
      port map(D => \soft_reset_reg_m[0]\, CLK => 
        CORECONFIGP_0_APB_S_PCLK, EN => \state_0\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg_m_reto[0]\);
    
    \soft_reset_reg[15]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(15), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[15]_net_1\);
    
    \prdata_0_iv_RNO[11]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \control_reg_1_m_1[0]\, B => 
        \soft_reset_reg[11]_net_1\, Y => \soft_reset_reg_m_0[11]\);
    
    \paddr[12]\ : SLE
      port map(D => \paddr_60\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => VCC_net_1, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \paddr[12]_net_1\);
    
    \FIC_2_APB_M_PRDATA_0[10]\ : SLE
      port map(D => \prdata[10]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state_0\, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(10));
    
    psel : SLE
      port map(D => \state_d_i[2]\, CLK => 
        CORECONFIGP_0_APB_S_PCLK_i, EN => VCC_net_1, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => \psel\);
    
    \soft_reset_reg[2]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(2), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[2]_net_1\);
    
    \paddr[13]\ : SLE
      port map(D => \paddr_61\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => VCC_net_1, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \paddr[13]_net_1\);
    
    \FIC_2_APB_M_PRDATA_0[7]\ : SLE
      port map(D => \prdata[7]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state_0\, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(7));
    
    un11_int_psel : CFG3
      generic map(INIT => x"01")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), C => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), Y => 
        N_468);
    
    \soft_reset_reg[14]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(14), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[14]_net_1\);
    
    prdata_0_iv_1_N_3L3 : CFG4
      generic map(INIT => x"FEFF")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), C => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), D => 
        \CORECONFIGP_0_CONFIG1_DONE\, Y => \prdata_0_iv_1_N_3L3\);
    
    \prdata_0_iv[1]\ : CFG4
      generic map(INIT => x"FFEA")

      port map(A => \soft_reset_reg_m[1]\, B => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, C => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(1), D => 
        \control_reg_1_m[1]\, Y => \prdata[1]\);
    
    \prdata_0_iv[3]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => CORECONFIGP_0_MDDR_APBmslave_PRDATA(3), B => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, C => 
        \soft_reset_reg_m[3]\, Y => \prdata[3]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    un6_int_psel_1 : CFG3
      generic map(INIT => x"80")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE, B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE, C => 
        \paddr[13]_net_1\, Y => \un6_int_psel_1\);
    
    \FIC_2_APB_M_PRDATA_0[15]\ : SLE
      port map(D => \prdata[15]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state_0\, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(15));
    
    \prdata_0_iv_RNO[14]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \control_reg_1_m_1[0]\, B => N_486, C => 
        N_471, D => \soft_reset_reg[14]_net_1\, Y => 
        \soft_reset_reg_m[14]\);
    
    un8_int_psel : CFG4
      generic map(INIT => x"4000")

      port map(A => \paddr[15]_net_1\, B => N_468, C => \psel\, D
         => \un6_int_psel_1\, Y => \un8_int_psel\);
    
    \soft_reset_reg[8]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(8), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[8]_net_1\);
    
    \prdata_0_iv_RNO[10]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \control_reg_1_m_1[0]\, B => 
        \soft_reset_reg[10]_net_1\, Y => \soft_reset_reg_m_0[10]\);
    
    \prdata_0_iv[10]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \soft_reset_reg_m_0[10]\, B => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(10), C => 
        int_prdata_4_sqmuxa_out_0, D => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, Y => \prdata[10]\);
    
    un20_int_psel : CFG3
      generic map(INIT => x"02")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), C => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), Y => 
        N_471);
    
    un1_next_FIC_2_APB_M_PREADY_0_sqmuxa_0 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \un1_fic_2_apb_m_psel\, B => \state_0\, C => 
        \state_d[2]\, D => pready, Y => 
        un1_next_FIC_2_APB_M_PREADY_0_sqmuxa);
    
    \prdata_0_iv_RNO[6]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \control_reg_1_m_1[0]\, B => 
        \soft_reset_reg[6]_net_1\, Y => \soft_reset_reg_m_0[6]\);
    
    \prdata_0_iv_RNO[7]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \control_reg_1_m_1[0]\, B => N_486, C => 
        N_471, D => \soft_reset_reg[7]_net_1\, Y => 
        \soft_reset_reg_m[7]\);
    
    MDDR_PENABLE_0_1 : CFG4
      generic map(INIT => x"0100")

      port map(A => \paddr[12]_net_1\, B => \paddr[13]_net_1\, C
         => \paddr[15]_net_1\, D => \state_0\, Y => 
        \MDDR_PENABLE_0_1\);
    
    \FIC_2_APB_M_PRDATA_0[11]\ : SLE
      port map(D => \prdata[11]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state_0\, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(11));
    
    \soft_reset_reg[0]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(0), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[0]_net_1\);
    
    \pwdata[1]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(1), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(1));
    
    \prdata_0_iv_RNO[4]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \control_reg_1_m_1[0]\, B => 
        \soft_reset_reg[4]_net_1\, Y => \soft_reset_reg_m_0[4]\);
    
    un1_fic_2_apb_m_psel : CFG2
      generic map(INIT => x"4")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE, B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx, Y => 
        \un1_fic_2_apb_m_psel\);
    
    \soft_reset_reg[1]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(1), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[1]_net_1\);
    
    \paddr[9]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(9), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(9));
    
    un1_next_FIC_2_APB_M_PREADY_0_sqmuxa_0_a3 : CFG2
      generic map(INIT => x"8")

      port map(A => \state_d[2]\, B => \un1_fic_2_apb_m_psel\, Y
         => \state_ns[0]\);
    
    \prdata_0_iv[9]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => CORECONFIGP_0_MDDR_APBmslave_PRDATA(9), B => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, C => 
        \soft_reset_reg_m[9]\, Y => \prdata[9]\);
    
    \paddr[15]\ : SLE
      port map(D => \paddr_63\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => VCC_net_1, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \paddr[15]_net_1\);
    
    \prdata_0_iv[12]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => CORECONFIGP_0_MDDR_APBmslave_PRDATA(12), B
         => \CORECONFIGP_0_MDDR_APBmslave_PSELx\, C => 
        \soft_reset_reg_m[12]\, Y => \prdata[12]\);
    
    int_prdata_3_sqmuxa_0 : CFG2
      generic map(INIT => x"8")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), Y => 
        \int_prdata_3_sqmuxa_0\);
    
    \FIC_2_APB_M_PRDATA_0[12]\ : SLE
      port map(D => \prdata[12]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state_0\, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(12));
    
    \control_reg_1[0]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(0), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un8_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \CORECONFIGP_0_CONFIG1_DONE\);
    
    \soft_reset_reg[5]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(5), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[5]_net_1\);
    
    \prdata_0_iv[14]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => CORECONFIGP_0_MDDR_APBmslave_PRDATA(14), B
         => \CORECONFIGP_0_MDDR_APBmslave_PSELx\, C => 
        \soft_reset_reg_m[14]\, Y => \prdata[14]\);
    
    \FIC_2_APB_M_PRDATA_0[14]\ : SLE
      port map(D => \prdata[14]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state_0\, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(14));
    
    psel_RNIPF3R : CFG2
      generic map(INIT => x"7")

      port map(A => \psel\, B => \paddr[15]_net_1\, Y => 
        \control_reg_1_m_1[0]\);
    
    \paddr[3]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(3));
    
    INIT_DONE_q2 : SLE
      port map(D => \INIT_DONE_q1\, CLK => 
        CORECONFIGP_0_APB_S_PCLK, EN => VCC_net_1, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INIT_DONE_q2\);
    
    \prdata_0_iv[5]\ : CFG4
      generic map(INIT => x"FFEA")

      port map(A => \soft_reset_reg_m[5]\, B => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, C => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(5), D => 
        \int_prdata_3_sqmuxa\, Y => \prdata[5]\);
    
    \paddr_RNI09N31[12]\ : CFG3
      generic map(INIT => x"01")

      port map(A => \paddr[12]_net_1\, B => \paddr[13]_net_1\, C
         => \paddr[15]_net_1\, Y => \paddr_RNI09N31[12]_net_1\);
    
    state_s0_0_a2_i : CFG2
      generic map(INIT => x"E")

      port map(A => \state_0\, B => \state[0]_net_1\, Y => 
        \state_d_i[2]\);
    
    pwrite : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE, CLK => 
        CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWRITE);
    
    MDDR_PENABLE_0 : SLE
      port map(D => \MDDR_PENABLE_0_1\, CLK => 
        CORECONFIGP_0_APB_S_PCLK_i, EN => VCC_net_1, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE);
    
    \soft_reset_reg[10]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(10), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[10]_net_1\);
    
    \soft_reset_reg[4]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(4), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[4]_net_1\);
    
    \prdata_0_iv[13]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => CORECONFIGP_0_MDDR_APBmslave_PRDATA(13), B
         => \CORECONFIGP_0_MDDR_APBmslave_PSELx\, C => 
        \soft_reset_reg_m[13]\, Y => \prdata[13]\);
    
    \pwdata[6]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(6), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(6));
    
    \prdata_0_iv_RNO[8]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \control_reg_1_m_1[0]\, B => N_486, C => 
        N_471, D => \soft_reset_reg[8]_net_1\, Y => 
        \soft_reset_reg_m[8]\);
    
    \prdata_0_iv[16]\ : CFG4
      generic map(INIT => x"ECCC")

      port map(A => int_prdata_4_sqmuxa_out_0, B => 
        \prdata_0_iv_1[16]\, C => \soft_reset_reg[16]_net_1\, D
         => \control_reg_1_m_1[0]\, Y => \prdata[16]\);
    
    \prdata_0_iv_RNO[12]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \control_reg_1_m_1[0]\, B => N_486, C => 
        N_471, D => \soft_reset_reg[12]_net_1\, Y => 
        \soft_reset_reg_m[12]\);
    
    int_prdata_5_sqmuxa : CFG4
      generic map(INIT => x"0080")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), C => 
        \prdata_0_iv_1_1[0]\, D => N_486, Y => 
        \prdata_0_iv_1[16]\);
    
    \state_ns_0[1]\ : CFG3
      generic map(INIT => x"F2")

      port map(A => \state_0\, B => pready, C => \state[0]_net_1\, 
        Y => \state_ns[1]\);
    
    \pwdata[11]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(11), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(11));
    
    \paddr[6]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(6), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(6));
    
    FIC_2_APB_M_PSLVERR_0 : SLE
      port map(D => pslverr, CLK => CORECONFIGP_0_APB_S_PCLK, EN
         => \state_0\, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR);
    
    \pwdata[12]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(12), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(12));
    
    \prdata_0_iv[0]\ : CFG4
      generic map(INIT => x"FFF8")

      port map(A => CORECONFIGP_0_MDDR_APBmslave_PSELx_reto, B
         => CORECONFIGP_0_MDDR_APBmslave_PRDATA_reto_0, C => 
        \soft_reset_reg_m_reto[0]\, D => \prdata_0_iv_1_reto[0]\, 
        Y => m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(0));
    
    \paddr_RNIEI071[13]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \paddr[13]_net_1\, B => \paddr[15]_net_1\, C
         => \psel\, Y => N_486);
    
    \prdata_0_iv_RNO[5]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \control_reg_1_m_1[0]\, B => N_486, C => 
        N_471, D => \soft_reset_reg[5]_net_1\, Y => 
        \soft_reset_reg_m[5]\);
    
    \paddr[4]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(4));
    
    \pwdata[9]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(9), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(9));
    
    \prdata_0_iv[15]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => CORECONFIGP_0_MDDR_APBmslave_PRDATA(15), B
         => \CORECONFIGP_0_MDDR_APBmslave_PSELx\, C => 
        \soft_reset_reg_m[15]\, Y => \prdata[15]\);
    
    \prdata_0_iv[7]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => CORECONFIGP_0_MDDR_APBmslave_PRDATA(7), B => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, C => 
        \soft_reset_reg_m[7]\, Y => \prdata[7]\);
    
    \state[1]\ : SLE
      port map(D => \state_ns[1]\, CLK => 
        CORECONFIGP_0_APB_S_PCLK, EN => VCC_net_1, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \state_0\);
    
    \soft_reset_reg[13]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(13), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[13]_net_1\);
    
    \FIC_2_APB_M_PRDATA_0[17]\ : SLE
      port map(D => \prdata_0_iv_1[16]\, CLK => 
        CORECONFIGP_0_APB_S_PCLK, EN => \state_0\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(17));
    
    psel_RNIQRM21 : CFG3
      generic map(INIT => x"15")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), B => 
        \paddr[15]_net_1\, C => \psel\, Y => \prdata_0_iv_1_1[0]\);
    
    \prdata_0_iv_RNO[2]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \control_reg_1_m_1[0]\, B => N_486, C => 
        N_471, D => \soft_reset_reg[2]_net_1\, Y => 
        \soft_reset_reg_m[2]\);
    
    \pwdata[15]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(15), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(15));
    
    \pwdata[5]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(5), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(5));
    
    INIT_DONE_q1 : SLE
      port map(D => INIT_DONE, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => VCC_net_1, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \INIT_DONE_q1\);
    
    FIC_2_APB_M_PRDATA_0_ret : SLE
      port map(D => \prdata_0_iv_1[0]_net_1\, CLK => 
        CORECONFIGP_0_APB_S_PCLK, EN => \state_0\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \prdata_0_iv_1_reto[0]\);
    
    \prdata_0_iv_RNO_1[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \psel\, B => \paddr[15]_net_1\, Y => 
        soft_N_6_0);
    
    state_s0_0_a2 : CFG2
      generic map(INIT => x"1")

      port map(A => \state_0\, B => \state[0]_net_1\, Y => 
        \state_d[2]\);
    
    \prdata_0_iv[6]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \soft_reset_reg_m_0[6]\, B => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(6), C => 
        int_prdata_4_sqmuxa_out_0, D => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, Y => \prdata[6]\);
    
    \prdata_0_iv[2]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => CORECONFIGP_0_MDDR_APBmslave_PRDATA(2), B => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, C => 
        \soft_reset_reg_m[2]\, Y => \prdata[2]\);
    
    un17_int_psel : CFG4
      generic map(INIT => x"4000")

      port map(A => \paddr[15]_net_1\, B => N_471, C => \psel\, D
         => \un6_int_psel_1\, Y => \un17_int_psel\);
    
    \prdata_0_iv[8]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => CORECONFIGP_0_MDDR_APBmslave_PRDATA(8), B => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, C => 
        \soft_reset_reg_m[8]\, Y => \prdata[8]\);
    
    \prdata_0_iv[4]\ : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \soft_reset_reg_m_0[4]\, B => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(4), C => 
        int_prdata_4_sqmuxa_out_0, D => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, Y => \prdata[4]\);
    
    \paddr[10]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(10), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(10));
    
    paddr_61 : CFG3
      generic map(INIT => x"D8")

      port map(A => \state_d[2]\, B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(13), C => 
        \paddr[13]_net_1\, Y => \paddr_61\);
    
    \soft_reset_reg[9]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(9), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[9]_net_1\);
    
    \soft_reset_reg[11]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(11), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[11]_net_1\);
    
    \pwdata[2]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(2), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(2));
    
    prdata_0_iv_1_N_4L6 : CFG4
      generic map(INIT => x"DFFF")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), C => 
        \prdata_0_iv_1_1[0]\, D => \INIT_DONE_q2\, Y => 
        \prdata_0_iv_1_N_4L6\);
    
    \soft_reset_reg[16]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(16), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[16]_net_1\);
    
    int_prdata_3_sqmuxa : CFG4
      generic map(INIT => x"0020")

      port map(A => \control_reg_1_m_1[0]\, B => N_486, C => 
        \int_prdata_3_sqmuxa_0\, D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), Y => 
        \int_prdata_3_sqmuxa\);
    
    \FIC_2_APB_M_PRDATA_0[2]\ : SLE
      port map(D => \prdata[2]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state_0\, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(2));
    
    \pwdata[14]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(14), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(14));
    
    \prdata_0_iv_RNO_0[1]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \control_reg_1_m_1[0]\, B => N_486, C => 
        N_468, D => \CORECONFIGP_0_CONFIG2_DONE\, Y => 
        \control_reg_1_m[1]\);
    
    \pwdata[3]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(3), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(3));
    
    \prdata_0_iv_1[0]\ : CFG4
      generic map(INIT => x"1511")

      port map(A => N_486, B => \prdata_0_iv_1_N_4L6\, C => 
        \prdata_0_iv_1_N_3L3\, D => \control_reg_1_m_1[0]\, Y => 
        \prdata_0_iv_1[0]_net_1\);
    
    FIC_2_APB_M_PRDATA_0_ret_1_RNO : CFG4
      generic map(INIT => x"B000")

      port map(A => \FIC_2_APB_M_PRDATA_0_ret_1_RNO_0\, B => 
        \psel\, C => N_471, D => \soft_reset_reg[0]_net_1\, Y => 
        \soft_reset_reg_m[0]\);
    
    \prdata_0_iv_RNO[9]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \control_reg_1_m_1[0]\, B => N_486, C => 
        N_471, D => \soft_reset_reg[9]_net_1\, Y => 
        \soft_reset_reg_m[9]\);
    
    \FIC_2_APB_M_PRDATA_0[3]\ : SLE
      port map(D => \prdata[3]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state_0\, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(3));
    
    \paddr[8]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(8), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(8));
    
    \prdata_0_iv_RNO[1]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => soft_N_6_0, B => N_486, C => N_471, D => 
        \soft_reset_reg[1]_net_1\, Y => \soft_reset_reg_m[1]\);
    
    \FIC_2_APB_M_PRDATA_0[1]\ : SLE
      port map(D => \prdata[1]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state_0\, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(1));
    
    \prdata_0_iv_RNO[13]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => \control_reg_1_m_1[0]\, B => N_486, C => 
        N_471, D => \soft_reset_reg[13]_net_1\, Y => 
        \soft_reset_reg_m[13]\);
    
    \soft_reset_reg[7]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(7), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[7]_net_1\);
    
    \soft_reset_reg[12]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(12), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[12]_net_1\);
    
    \paddr_RNI2KTI1[12]\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \paddr[12]_net_1\, B => \paddr[13]_net_1\, C
         => \paddr[15]_net_1\, D => \psel\, Y => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\);
    
    paddr_60 : CFG3
      generic map(INIT => x"D8")

      port map(A => \state_d[2]\, B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(12), C => 
        \paddr[12]_net_1\, Y => \paddr_60\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb_CCC_0_FCCC is

    port( m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC : in    std_logic;
          FAB_CCC_LOCK                              : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz                 : out   std_logic
        );

end m2s010_som_sb_CCC_0_FCCC;

architecture DEF_ARCH of m2s010_som_sb_CCC_0_FCCC is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CCC

            generic (INIT:std_logic_vector(209 downto 0) := "00" & x"0000000000000000000000000000000000000000000000000000"; 
        VCOFREQUENCY:real := 0.0);

    port( Y0              : out   std_logic;
          Y1              : out   std_logic;
          Y2              : out   std_logic;
          Y3              : out   std_logic;
          PRDATA          : out   std_logic_vector(7 downto 0);
          LOCK            : out   std_logic;
          BUSY            : out   std_logic;
          CLK0            : in    std_logic := 'U';
          CLK1            : in    std_logic := 'U';
          CLK2            : in    std_logic := 'U';
          CLK3            : in    std_logic := 'U';
          NGMUX0_SEL      : in    std_logic := 'U';
          NGMUX1_SEL      : in    std_logic := 'U';
          NGMUX2_SEL      : in    std_logic := 'U';
          NGMUX3_SEL      : in    std_logic := 'U';
          NGMUX0_HOLD_N   : in    std_logic := 'U';
          NGMUX1_HOLD_N   : in    std_logic := 'U';
          NGMUX2_HOLD_N   : in    std_logic := 'U';
          NGMUX3_HOLD_N   : in    std_logic := 'U';
          NGMUX0_ARST_N   : in    std_logic := 'U';
          NGMUX1_ARST_N   : in    std_logic := 'U';
          NGMUX2_ARST_N   : in    std_logic := 'U';
          NGMUX3_ARST_N   : in    std_logic := 'U';
          PLL_BYPASS_N    : in    std_logic := 'U';
          PLL_ARST_N      : in    std_logic := 'U';
          PLL_POWERDOWN_N : in    std_logic := 'U';
          GPD0_ARST_N     : in    std_logic := 'U';
          GPD1_ARST_N     : in    std_logic := 'U';
          GPD2_ARST_N     : in    std_logic := 'U';
          GPD3_ARST_N     : in    std_logic := 'U';
          PRESET_N        : in    std_logic := 'U';
          PCLK            : in    std_logic := 'U';
          PSEL            : in    std_logic := 'U';
          PENABLE         : in    std_logic := 'U';
          PWRITE          : in    std_logic := 'U';
          PADDR           : in    std_logic_vector(7 downto 2) := (others => 'U');
          PWDATA          : in    std_logic_vector(7 downto 0) := (others => 'U');
          CLK0_PAD        : in    std_logic := 'U';
          CLK1_PAD        : in    std_logic := 'U';
          CLK2_PAD        : in    std_logic := 'U';
          CLK3_PAD        : in    std_logic := 'U';
          GL0             : out   std_logic;
          GL1             : out   std_logic;
          GL2             : out   std_logic;
          GL3             : out   std_logic;
          RCOSC_25_50MHZ  : in    std_logic := 'U';
          RCOSC_1MHZ      : in    std_logic := 'U';
          XTLOSC          : in    std_logic := 'U'
        );
  end component;

    signal GL0_net, VCC_net_1, GND_net_1 : std_logic;
    signal nc8, nc7, nc6, nc2, nc5, nc4, nc3, nc1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    GL0_INST : CLKINT
      port map(A => GL0_net, Y => m2s010_som_sb_0_CCC_71MHz);
    
    CCC_INST : CCC

              generic map(INIT => "00" & x"000007F88000044D64000318C6318C1F18C61E40404040404613",
         VCOFREQUENCY => 568.0)

      port map(Y0 => OPEN, Y1 => OPEN, Y2 => OPEN, Y3 => OPEN, 
        PRDATA(7) => nc8, PRDATA(6) => nc7, PRDATA(5) => nc6, 
        PRDATA(4) => nc2, PRDATA(3) => nc5, PRDATA(2) => nc4, 
        PRDATA(1) => nc3, PRDATA(0) => nc1, LOCK => FAB_CCC_LOCK, 
        BUSY => OPEN, CLK0 => VCC_net_1, CLK1 => VCC_net_1, CLK2
         => VCC_net_1, CLK3 => VCC_net_1, NGMUX0_SEL => GND_net_1, 
        NGMUX1_SEL => GND_net_1, NGMUX2_SEL => GND_net_1, 
        NGMUX3_SEL => GND_net_1, NGMUX0_HOLD_N => VCC_net_1, 
        NGMUX1_HOLD_N => VCC_net_1, NGMUX2_HOLD_N => VCC_net_1, 
        NGMUX3_HOLD_N => VCC_net_1, NGMUX0_ARST_N => VCC_net_1, 
        NGMUX1_ARST_N => VCC_net_1, NGMUX2_ARST_N => VCC_net_1, 
        NGMUX3_ARST_N => VCC_net_1, PLL_BYPASS_N => VCC_net_1, 
        PLL_ARST_N => VCC_net_1, PLL_POWERDOWN_N => VCC_net_1, 
        GPD0_ARST_N => VCC_net_1, GPD1_ARST_N => VCC_net_1, 
        GPD2_ARST_N => VCC_net_1, GPD3_ARST_N => VCC_net_1, 
        PRESET_N => GND_net_1, PCLK => VCC_net_1, PSEL => 
        VCC_net_1, PENABLE => VCC_net_1, PWRITE => VCC_net_1, 
        PADDR(7) => VCC_net_1, PADDR(6) => VCC_net_1, PADDR(5)
         => VCC_net_1, PADDR(4) => VCC_net_1, PADDR(3) => 
        VCC_net_1, PADDR(2) => VCC_net_1, PWDATA(7) => VCC_net_1, 
        PWDATA(6) => VCC_net_1, PWDATA(5) => VCC_net_1, PWDATA(4)
         => VCC_net_1, PWDATA(3) => VCC_net_1, PWDATA(2) => 
        VCC_net_1, PWDATA(1) => VCC_net_1, PWDATA(0) => VCC_net_1, 
        CLK0_PAD => GND_net_1, CLK1_PAD => GND_net_1, CLK2_PAD
         => GND_net_1, CLK3_PAD => GND_net_1, GL0 => GL0_net, GL1
         => OPEN, GL2 => OPEN, GL3 => OPEN, RCOSC_25_50MHZ => 
        GND_net_1, RCOSC_1MHZ => GND_net_1, XTLOSC => 
        m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb_OTH_SPI_1_SS0_IO is

    port( SPI_1_SS0_OTH_0                      : inout std_logic := 'Z';
          OTH_SPI_1_SS0_Y_0                    : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE : in    std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F    : in    std_logic
        );

end m2s010_som_sb_OTH_SPI_1_SS0_IO;

architecture DEF_ARCH of m2s010_som_sb_OTH_SPI_1_SS0_IO is 

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    U0_0 : BIBUF
      port map(PAD => SPI_1_SS0_OTH_0, D => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F, E => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE, Y => 
        OTH_SPI_1_SS0_Y_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb_FABOSC_0_OSC is

    port( XTL                                       : in    std_logic;
          m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC : out   std_logic;
          FABOSC_0_RCOSC_25_50MHZ_O2F               : out   std_logic
        );

end m2s010_som_sb_FABOSC_0_OSC;

architecture DEF_ARCH of m2s010_som_sb_FABOSC_0_OSC is 

  component RCOSC_25_50MHZ_FAB
    port( A      : in    std_logic := 'U';
          CLKOUT : out   std_logic
        );
  end component;

  component RCOSC_25_50MHZ
    generic (FREQUENCY:real := 50.0);

    port( CLKOUT : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component XTLOSC
    generic (MODE:std_logic_vector(1 downto 0) := "11"; 
        FREQUENCY:real := 20.0);

    port( XTL    : in    std_logic := 'U';
          CLKOUT : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal N_RCOSC_25_50MHZ_CLKINT, N_RCOSC_25_50MHZ_CLKOUT, 
        GND_net_1, VCC_net_1 : std_logic;

begin 


    I_RCOSC_25_50MHZ_FAB : RCOSC_25_50MHZ_FAB
      port map(A => N_RCOSC_25_50MHZ_CLKOUT, CLKOUT => 
        N_RCOSC_25_50MHZ_CLKINT);
    
    I_RCOSC_25_50MHZ : RCOSC_25_50MHZ
      generic map(FREQUENCY => 50.0)

      port map(CLKOUT => N_RCOSC_25_50MHZ_CLKOUT);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    I_XTLOSC : XTLOSC
      generic map(MODE => "11", FREQUENCY => 20.0)

      port map(XTL => XTL, CLKOUT => 
        m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC);
    
    I_RCOSC_25_50MHZ_FAB_CLKINT : CLKINT
      port map(A => N_RCOSC_25_50MHZ_CLKINT, Y => 
        FABOSC_0_RCOSC_25_50MHZ_O2F);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb is

    port( MDDR_DQS                                  : inout std_logic_vector(1 downto 0) := (others => 'Z');
          MDDR_DQ                                   : inout std_logic_vector(15 downto 0) := (others => 'Z');
          MDDR_DM_RDQS                              : inout std_logic_vector(1 downto 0) := (others => 'Z');
          MDDR_BA                                   : out   std_logic_vector(2 downto 0);
          MDDR_ADDR                                 : out   std_logic_vector(15 downto 0);
          CoreAPB3_0_APBmslave0_PADDR               : out   std_logic_vector(7 downto 0);
          m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR    : out   std_logic_vector(15 downto 12);
          CoreAPB3_0_APBmslave0_PWDATA              : out   std_logic_vector(7 downto 0);
          MAC_MII_TXD_c                             : out   std_logic_vector(3 downto 0);
          CoreAPB3_0_APBmslave0_PRDATA_m            : in    std_logic_vector(7 downto 0);
          Y_net_0                                   : in    std_logic_vector(3 downto 0);
          MAC_MII_RXD_c                             : in    std_logic_vector(3 downto 0);
          SPI_1_SS0_OTH_0                           : inout std_logic := 'Z';
          DEBOUNCE_OUT_net_0_0                      : in    std_logic;
          GPIO_7_PADI_0                             : inout std_logic := 'Z';
          GPIO_6_PAD_0                              : inout std_logic := 'Z';
          GPIO_1_BI_0                               : inout std_logic := 'Z';
          SPI_1_SS0_CAM_0                           : inout std_logic := 'Z';
          SPI_1_CLK_0                               : inout std_logic := 'Z';
          SPI_0_SS1                                 : out   std_logic;
          SPI_0_SS0                                 : inout std_logic := 'Z';
          SPI_0_DO                                  : out   std_logic;
          SPI_0_DI                                  : in    std_logic;
          SPI_0_CLK                                 : inout std_logic := 'Z';
          MMUART_1_TXD                              : out   std_logic;
          MMUART_1_RXD                              : in    std_logic;
          MDDR_WE_N                                 : out   std_logic;
          MDDR_RESET_N                              : out   std_logic;
          MDDR_RAS_N                                : out   std_logic;
          MDDR_ODT                                  : out   std_logic;
          MDDR_DQS_TMATCH_0_OUT                     : out   std_logic;
          MDDR_DQS_TMATCH_0_IN                      : in    std_logic;
          MDDR_CS_N                                 : out   std_logic;
          MDDR_CKE                                  : out   std_logic;
          MDDR_CAS_N                                : out   std_logic;
          I2C_1_SDA                                 : inout std_logic := 'Z';
          I2C_1_SCL                                 : inout std_logic := 'Z';
          GPIO_31_BI                                : inout std_logic := 'Z';
          GPIO_26_BI                                : inout std_logic := 'Z';
          GPIO_25_BI                                : inout std_logic := 'Z';
          GPIO_20_OUT                               : out   std_logic;
          GPIO_18_BI                                : inout std_logic := 'Z';
          GPIO_17_BI                                : inout std_logic := 'Z';
          GPIO_16_BI                                : inout std_logic := 'Z';
          GPIO_15_BI                                : inout std_logic := 'Z';
          GPIO_14_BI                                : inout std_logic := 'Z';
          GPIO_12_BI                                : inout std_logic := 'Z';
          GPIO_4_BI                                 : inout std_logic := 'Z';
          GPIO_3_BI                                 : inout std_logic := 'Z';
          GPIO_0_BI                                 : inout std_logic := 'Z';
          CoreAPB3_0_APBmslave0_PENABLE             : out   std_logic;
          m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx    : out   std_logic;
          CoreAPB3_0_APBmslave0_PWRITE              : out   std_logic;
          MAC_MII_MDC_c                             : out   std_logic;
          GPIO_22_M2F_c                             : out   std_logic;
          GPIO_21_M2F_c                             : out   std_logic;
          m2s010_som_sb_0_GPIO_28_SW_RESET          : out   std_logic;
          MMUART_0_TXD_M2F_c                        : out   std_logic;
          GPIO_24_M2F_c                             : out   std_logic;
          GPIO_5_M2F_c                              : out   std_logic;
          GPIO_8_M2F_c                              : out   std_logic;
          GPIO_11_M2F_c                             : out   std_logic;
          MAC_MII_TX_EN_c                           : out   std_logic;
          MAC_MII_COL_c                             : in    std_logic;
          MAC_MII_CRS_c                             : in    std_logic;
          CommsFPGA_top_0_INT                       : in    std_logic;
          CoreAPB3_0_APBmslave0_PREADY_i_m_i        : in    std_logic;
          DEBOUNCE_OUT_1_c                          : in    std_logic;
          DEBOUNCE_OUT_2_c                          : in    std_logic;
          MMUART_0_RXD_F2M_c                        : in    std_logic;
          MAC_MII_RX_CLK_c                          : in    std_logic;
          MAC_MII_RX_DV_c                           : in    std_logic;
          MAC_MII_RX_ER_c                           : in    std_logic;
          MAC_MII_TX_CLK_c                          : in    std_logic;
          MDDR_CLK_N                                : out   std_logic;
          MDDR_CLK                                  : out   std_logic;
          XTL                                       : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz                 : out   std_logic;
          m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC : inout std_logic := 'Z';
          SPI_1_DI_CAM_c                            : in    std_logic;
          SPI_1_DI_OTH_c                            : in    std_logic;
          CommsFPGA_top_0_CAMERA_NODE               : in    std_logic;
          DEVRST_N                                  : in    std_logic;
          m2s010_som_sb_0_POWER_ON_RESET_N          : out   std_logic;
          MAC_MII_MDIO                              : inout std_logic := 'Z';
          SPI_1_DO_CAM_c                            : inout std_logic := 'Z';
          SPI_1_DO_OTH                              : out   std_logic
        );

end m2s010_som_sb;

architecture DEF_ARCH of m2s010_som_sb is 

  component m2s010_som_sb_GPIO_1_IO
    port( GPIO_1_BI_0                       : inout   std_logic;
          GPIO_1_in_0                       : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_1_M2F_OE : in    std_logic := 'U';
          GPIO_1_M2F                        : in    std_logic := 'U'
        );
  end component;

  component m2s010_som_sb_CAM_SPI_1_CLK_IO
    port( CAM_SPI_1_CLK_Y_0                    : out   std_logic;
          SPI_1_CLK_0                          : inout   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE : in    std_logic := 'U';
          m2s010_som_sb_MSS_0_SPI_1_CLK_M2F    : in    std_logic := 'U'
        );
  end component;

  component m2s010_som_sb_GPIO_7_IO
    port( GPIO_7_PADI_0                     : inout   std_logic;
          GPIO_7_Y_0                        : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_7_M2F_OE : in    std_logic := 'U';
          m2s010_som_sb_MSS_0_GPIO_7_M2F    : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component m2s010_som_sb_CAM_SPI_1_SS0_IO
    port( SPI_1_SS0_CAM_0                      : inout   std_logic;
          CAM_SPI_1_SS0_Y_0                    : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE : in    std_logic := 'U';
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F    : in    std_logic := 'U'
        );
  end component;

  component m2s010_som_sb_MSS
    port( CORECONFIGP_0_MDDR_APBmslave_PWDATA              : in    std_logic_vector(15 downto 0) := (others => 'U');
          CORECONFIGP_0_MDDR_APBmslave_PADDR               : in    std_logic_vector(10 downto 2) := (others => 'U');
          MAC_MII_RXD_c                                    : in    std_logic_vector(3 downto 0) := (others => 'U');
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA  : in    std_logic_vector(17 downto 0) := (others => 'U');
          Y_net_0                                          : in    std_logic_vector(3 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PRDATA_m                   : in    std_logic_vector(7 downto 0) := (others => 'U');
          CORECONFIGP_0_MDDR_APBmslave_PRDATA              : out   std_logic_vector(15 downto 1);
          MAC_MII_TXD_c                                    : out   std_logic_vector(3 downto 0);
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA  : out   std_logic_vector(16 downto 0);
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR   : out   std_logic_vector(15 downto 2);
          CoreAPB3_0_APBmslave0_PWDATA                     : out   std_logic_vector(7 downto 0);
          m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR           : out   std_logic_vector(15 downto 12);
          CoreAPB3_0_APBmslave0_PADDR                      : out   std_logic_vector(7 downto 0);
          MDDR_ADDR                                        : out   std_logic_vector(15 downto 0);
          MDDR_BA                                          : out   std_logic_vector(2 downto 0);
          MDDR_DM_RDQS                                     : inout   std_logic_vector(1 downto 0);
          MDDR_DQ                                          : inout   std_logic_vector(15 downto 0);
          MDDR_DQS                                         : inout   std_logic_vector(1 downto 0);
          CAM_SPI_1_CLK_Y_0                                : in    std_logic := 'U';
          GPIO_7_Y_0                                       : in    std_logic := 'U';
          GPIO_6_Y_0                                       : in    std_logic := 'U';
          DEBOUNCE_OUT_net_0_0                             : in    std_logic := 'U';
          GPIO_1_in_0                                      : in    std_logic := 'U';
          state_0                                          : in    std_logic := 'U';
          CORECONFIGP_0_MDDR_APBmslave_PRDATA_reto_0       : out   std_logic;
          MDDR_CLK                                         : out   std_logic;
          MDDR_CLK_N                                       : out   std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PWRITE              : in    std_logic := 'U';
          CORECONFIGP_0_MDDR_APBmslave_PSELx               : in    std_logic := 'U';
          CORECONFIGP_0_MDDR_APBmslave_PENABLE             : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz                        : in    std_logic := 'U';
          MAC_MII_TX_CLK_c                                 : in    std_logic := 'U';
          SPI_1_SS0_MX_Y                                   : in    std_logic := 'U';
          SPI_1_DI                                         : in    std_logic := 'U';
          MAC_MII_RX_ER_c                                  : in    std_logic := 'U';
          MAC_MII_RX_DV_c                                  : in    std_logic := 'U';
          MAC_MII_RX_CLK_c                                 : in    std_logic := 'U';
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR : in    std_logic := 'U';
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY  : in    std_logic := 'U';
          MMUART_0_RXD_F2M_c                               : in    std_logic := 'U';
          DEBOUNCE_OUT_2_c                                 : in    std_logic := 'U';
          DEBOUNCE_OUT_1_c                                 : in    std_logic := 'U';
          BIBUF_0_Y                                        : in    std_logic := 'U';
          FAB_CCC_LOCK                                     : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PREADY_i_m_i               : in    std_logic := 'U';
          CommsFPGA_top_0_INT                              : in    std_logic := 'U';
          MAC_MII_CRS_c                                    : in    std_logic := 'U';
          MAC_MII_COL_c                                    : in    std_logic := 'U';
          CORECONFIGP_0_MDDR_APBmslave_PSLVERR             : out   std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PREADY              : out   std_logic;
          MAC_MII_TX_EN_c                                  : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE             : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F                : out   std_logic;
          SPI_1_DO_CAM_c                                   : out   std_logic;
          GPIO_11_M2F_c                                    : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_CLK_M2F                : out   std_logic;
          GPIO_8_M2F_c                                     : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_7_M2F                   : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_7_M2F_OE                : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_6_M2F                   : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_6_M2F_OE                : out   std_logic;
          GPIO_5_M2F_c                                     : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE  : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx   : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE : out   std_logic;
          GPIO_24_M2F_c                                    : out   std_logic;
          MMUART_0_TXD_M2F_c                               : out   std_logic;
          m2s010_som_sb_0_GPIO_28_SW_RESET                 : out   std_logic;
          GPIO_21_M2F_c                                    : out   std_logic;
          GPIO_22_M2F_c                                    : out   std_logic;
          m2s010_som_sb_MSS_0_MAC_MII_MDO                  : out   std_logic;
          m2s010_som_sb_MSS_0_MAC_MII_MDO_EN               : out   std_logic;
          MAC_MII_MDC_c                                    : out   std_logic;
          GPIO_1_M2F                                       : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_1_M2F_OE                : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F          : out   std_logic;
          CoreAPB3_0_APBmslave0_PWRITE                     : out   std_logic;
          m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx           : out   std_logic;
          CoreAPB3_0_APBmslave0_PENABLE                    : out   std_logic;
          GPIO_0_BI                                        : inout   std_logic;
          GPIO_3_BI                                        : inout   std_logic;
          GPIO_4_BI                                        : inout   std_logic;
          GPIO_12_BI                                       : inout   std_logic;
          GPIO_14_BI                                       : inout   std_logic;
          GPIO_15_BI                                       : inout   std_logic;
          GPIO_16_BI                                       : inout   std_logic;
          GPIO_17_BI                                       : inout   std_logic;
          GPIO_18_BI                                       : inout   std_logic;
          GPIO_20_OUT                                      : out   std_logic;
          GPIO_25_BI                                       : inout   std_logic;
          GPIO_26_BI                                       : inout   std_logic;
          GPIO_31_BI                                       : inout   std_logic;
          I2C_1_SCL                                        : inout   std_logic;
          I2C_1_SDA                                        : inout   std_logic;
          MDDR_CAS_N                                       : out   std_logic;
          MDDR_CKE                                         : out   std_logic;
          MDDR_CS_N                                        : out   std_logic;
          MDDR_DQS_TMATCH_0_IN                             : in    std_logic := 'U';
          MDDR_DQS_TMATCH_0_OUT                            : out   std_logic;
          MDDR_ODT                                         : out   std_logic;
          MDDR_RAS_N                                       : out   std_logic;
          MDDR_RESET_N                                     : out   std_logic;
          MDDR_WE_N                                        : out   std_logic;
          MMUART_1_RXD                                     : in    std_logic := 'U';
          MMUART_1_TXD                                     : out   std_logic;
          SPI_0_CLK                                        : inout   std_logic;
          SPI_0_DI                                         : in    std_logic := 'U';
          SPI_0_DO                                         : out   std_logic;
          SPI_0_SS0                                        : inout   std_logic;
          SPI_0_SS1                                        : out   std_logic;
          CORECONFIGP_0_APB_S_PCLK_i                       : out   std_logic;
          CORECONFIGP_0_APB_S_PRESET_N                     : out   std_logic;
          CORECONFIGP_0_APB_S_PCLK                         : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CoreResetP
    port( CORECONFIGP_0_CONFIG2_DONE              : in    std_logic := 'U';
          CORECONFIGP_0_CONFIG1_DONE              : in    std_logic := 'U';
          CORECONFIGP_0_APB_S_PRESET_N            : in    std_logic := 'U';
          m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F : in    std_logic := 'U';
          m2s010_som_sb_0_POWER_ON_RESET_N        : in    std_logic := 'U';
          INIT_DONE                               : out   std_logic;
          FABOSC_0_RCOSC_25_50MHZ_O2F             : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz               : in    std_logic := 'U'
        );
  end component;

  component SYSRESET
    port( POWER_ON_RESET_N : out   std_logic;
          DEVRST_N         : in    std_logic := 'U'
        );
  end component;

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component OUTBUF
    generic (IOSTD:string := "");

    port( D   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component m2s010_som_sb_GPIO_6_IO
    port( GPIO_6_PAD_0                      : inout   std_logic;
          GPIO_6_Y_0                        : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_6_M2F_OE : in    std_logic := 'U';
          m2s010_som_sb_MSS_0_GPIO_6_M2F    : in    std_logic := 'U'
        );
  end component;

  component CoreConfigP
    port( CORECONFIGP_0_MDDR_APBmslave_PRDATA              : in    std_logic_vector(15 downto 1) := (others => 'U');
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA  : out   std_logic_vector(17 downto 0);
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR   : in    std_logic_vector(15 downto 2) := (others => 'U');
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA  : in    std_logic_vector(16 downto 0) := (others => 'U');
          CORECONFIGP_0_MDDR_APBmslave_PADDR               : out   std_logic_vector(10 downto 2);
          CORECONFIGP_0_MDDR_APBmslave_PWDATA              : out   std_logic_vector(15 downto 0);
          CORECONFIGP_0_MDDR_APBmslave_PRDATA_reto_0       : in    std_logic := 'U';
          state_0                                          : out   std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PSLVERR             : in    std_logic := 'U';
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx   : in    std_logic := 'U';
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE : in    std_logic := 'U';
          CORECONFIGP_0_MDDR_APBmslave_PREADY              : in    std_logic := 'U';
          CORECONFIGP_0_MDDR_APBmslave_PSELx               : out   std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PENABLE             : out   std_logic;
          INIT_DONE                                        : in    std_logic := 'U';
          CORECONFIGP_0_APB_S_PCLK_i                       : in    std_logic := 'U';
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE  : in    std_logic := 'U';
          CORECONFIGP_0_MDDR_APBmslave_PWRITE              : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY  : out   std_logic;
          CORECONFIGP_0_CONFIG2_DONE                       : out   std_logic;
          CORECONFIGP_0_CONFIG1_DONE                       : out   std_logic;
          CORECONFIGP_0_APB_S_PCLK                         : in    std_logic := 'U';
          CORECONFIGP_0_APB_S_PRESET_N                     : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component m2s010_som_sb_CCC_0_FCCC
    port( m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC : in    std_logic := 'U';
          FAB_CCC_LOCK                              : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz                 : out   std_logic
        );
  end component;

  component m2s010_som_sb_OTH_SPI_1_SS0_IO
    port( SPI_1_SS0_OTH_0                      : inout   std_logic;
          OTH_SPI_1_SS0_Y_0                    : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE : in    std_logic := 'U';
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F    : in    std_logic := 'U'
        );
  end component;

  component m2s010_som_sb_FABOSC_0_OSC
    port( XTL                                       : in    std_logic := 'U';
          m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC : out   std_logic;
          FABOSC_0_RCOSC_25_50MHZ_O2F               : out   std_logic
        );
  end component;

    signal BIBUF_0_Y, m2s010_som_sb_MSS_0_MAC_MII_MDO, 
        m2s010_som_sb_MSS_0_MAC_MII_MDO_EN, 
        \m2s010_som_sb_0_POWER_ON_RESET_N\, SPI_1_SS0_MX_Y, 
        \OTH_SPI_1_SS0_Y[0]\, \CAM_SPI_1_SS0_Y[0]\, SPI_1_DI, 
        \CAM_SPI_1_CLK_Y[0]\, 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE, 
        m2s010_som_sb_MSS_0_SPI_1_CLK_M2F, 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F, FAB_CCC_LOCK, 
        \m2s010_som_sb_0_CCC_71MHz\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[1]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[2]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[3]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[4]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[5]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[6]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[7]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[8]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[9]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[10]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[11]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[12]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[13]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[14]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[15]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[0]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[1]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[2]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[3]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[4]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[5]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[6]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[7]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[8]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[9]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[10]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[11]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[12]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[13]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[14]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[15]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[16]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[17]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA_reto[0]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[2]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[3]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[4]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[5]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[6]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[7]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[8]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[9]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[10]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[12]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[13]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[15]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[0]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[1]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[2]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[3]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[4]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[5]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[6]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[7]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[8]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[9]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[10]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[11]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[12]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[13]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[14]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[15]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[16]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[2]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[3]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[4]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[5]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[6]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[7]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[8]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[9]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[10]\, \state[1]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[0]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[1]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[2]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[3]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[4]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[5]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[6]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[7]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[8]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[9]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[10]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[11]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[12]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[13]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[14]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[15]\, 
        CORECONFIGP_0_MDDR_APBmslave_PSLVERR, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE, 
        CORECONFIGP_0_MDDR_APBmslave_PREADY, 
        CORECONFIGP_0_MDDR_APBmslave_PSELx, 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE, INIT_DONE, 
        CORECONFIGP_0_APB_S_PCLK_i, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE, 
        CORECONFIGP_0_MDDR_APBmslave_PWRITE, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY, 
        CORECONFIGP_0_CONFIG2_DONE, CORECONFIGP_0_CONFIG1_DONE, 
        CORECONFIGP_0_APB_S_PCLK, CORECONFIGP_0_APB_S_PRESET_N, 
        m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        FABOSC_0_RCOSC_25_50MHZ_O2F, \GPIO_1_in[0]\, 
        m2s010_som_sb_MSS_0_GPIO_1_M2F_OE, GPIO_1_M2F, 
        \GPIO_6_Y[0]\, m2s010_som_sb_MSS_0_GPIO_6_M2F_OE, 
        m2s010_som_sb_MSS_0_GPIO_6_M2F, \GPIO_7_Y[0]\, 
        m2s010_som_sb_MSS_0_GPIO_7_M2F_OE, 
        m2s010_som_sb_MSS_0_GPIO_7_M2F, GND_net_1, VCC_net_1
         : std_logic;
    signal nc2, nc4, nc3, nc1 : std_logic;

    for all : m2s010_som_sb_GPIO_1_IO
	Use entity work.m2s010_som_sb_GPIO_1_IO(DEF_ARCH);
    for all : m2s010_som_sb_CAM_SPI_1_CLK_IO
	Use entity work.m2s010_som_sb_CAM_SPI_1_CLK_IO(DEF_ARCH);
    for all : m2s010_som_sb_GPIO_7_IO
	Use entity work.m2s010_som_sb_GPIO_7_IO(DEF_ARCH);
    for all : m2s010_som_sb_CAM_SPI_1_SS0_IO
	Use entity work.m2s010_som_sb_CAM_SPI_1_SS0_IO(DEF_ARCH);
    for all : m2s010_som_sb_MSS
	Use entity work.m2s010_som_sb_MSS(DEF_ARCH);
    for all : CoreResetP
	Use entity work.CoreResetP(DEF_ARCH);
    for all : m2s010_som_sb_GPIO_6_IO
	Use entity work.m2s010_som_sb_GPIO_6_IO(DEF_ARCH);
    for all : CoreConfigP
	Use entity work.CoreConfigP(DEF_ARCH);
    for all : m2s010_som_sb_CCC_0_FCCC
	Use entity work.m2s010_som_sb_CCC_0_FCCC(DEF_ARCH);
    for all : m2s010_som_sb_OTH_SPI_1_SS0_IO
	Use entity work.m2s010_som_sb_OTH_SPI_1_SS0_IO(DEF_ARCH);
    for all : m2s010_som_sb_FABOSC_0_OSC
	Use entity work.m2s010_som_sb_FABOSC_0_OSC(DEF_ARCH);
begin 

    m2s010_som_sb_0_CCC_71MHz <= \m2s010_som_sb_0_CCC_71MHz\;
    m2s010_som_sb_0_POWER_ON_RESET_N <= 
        \m2s010_som_sb_0_POWER_ON_RESET_N\;

    GPIO_1 : m2s010_som_sb_GPIO_1_IO
      port map(GPIO_1_BI_0 => GPIO_1_BI_0, GPIO_1_in_0 => 
        \GPIO_1_in[0]\, m2s010_som_sb_MSS_0_GPIO_1_M2F_OE => 
        m2s010_som_sb_MSS_0_GPIO_1_M2F_OE, GPIO_1_M2F => 
        GPIO_1_M2F);
    
    CAM_SPI_1_CLK : m2s010_som_sb_CAM_SPI_1_CLK_IO
      port map(CAM_SPI_1_CLK_Y_0 => \CAM_SPI_1_CLK_Y[0]\, 
        SPI_1_CLK_0 => SPI_1_CLK_0, 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE, 
        m2s010_som_sb_MSS_0_SPI_1_CLK_M2F => 
        m2s010_som_sb_MSS_0_SPI_1_CLK_M2F);
    
    GPIO_7 : m2s010_som_sb_GPIO_7_IO
      port map(GPIO_7_PADI_0 => GPIO_7_PADI_0, GPIO_7_Y_0 => 
        \GPIO_7_Y[0]\, m2s010_som_sb_MSS_0_GPIO_7_M2F_OE => 
        m2s010_som_sb_MSS_0_GPIO_7_M2F_OE, 
        m2s010_som_sb_MSS_0_GPIO_7_M2F => 
        m2s010_som_sb_MSS_0_GPIO_7_M2F);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    CAM_SPI_1_SS0 : m2s010_som_sb_CAM_SPI_1_SS0_IO
      port map(SPI_1_SS0_CAM_0 => SPI_1_SS0_CAM_0, 
        CAM_SPI_1_SS0_Y_0 => \CAM_SPI_1_SS0_Y[0]\, 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE, 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F);
    
    m2s010_som_sb_MSS_0 : m2s010_som_sb_MSS
      port map(CORECONFIGP_0_MDDR_APBmslave_PWDATA(15) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[15]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(14) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[14]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(13) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[13]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(12) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[12]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(11) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[11]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(10) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[10]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(9) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[9]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(8) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[8]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(7) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[7]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(6) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[6]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(5) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[5]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(4) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[4]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(3) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[3]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(2) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[2]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(1) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[1]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(0) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[0]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(10) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[10]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(9) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[9]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(8) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[8]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(7) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[7]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(6) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[6]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(5) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[5]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(4) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[4]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(3) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[3]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(2) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[2]\, MAC_MII_RXD_c(3)
         => MAC_MII_RXD_c(3), MAC_MII_RXD_c(2) => 
        MAC_MII_RXD_c(2), MAC_MII_RXD_c(1) => MAC_MII_RXD_c(1), 
        MAC_MII_RXD_c(0) => MAC_MII_RXD_c(0), 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(17) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[17]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(16) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[16]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(15) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[15]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(14) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[14]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(13) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[13]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(12) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[12]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(11) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[11]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(10) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[10]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(9) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[9]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(8) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[8]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(7) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[7]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(6) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[6]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(5) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[5]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(4) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[4]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(3) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[3]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(2) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[2]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(1) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[1]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(0) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[0]\, 
        Y_net_0(3) => Y_net_0(3), Y_net_0(2) => Y_net_0(2), 
        Y_net_0(1) => Y_net_0(1), Y_net_0(0) => Y_net_0(0), 
        CoreAPB3_0_APBmslave0_PRDATA_m(7) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(7), 
        CoreAPB3_0_APBmslave0_PRDATA_m(6) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(6), 
        CoreAPB3_0_APBmslave0_PRDATA_m(5) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(5), 
        CoreAPB3_0_APBmslave0_PRDATA_m(4) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(4), 
        CoreAPB3_0_APBmslave0_PRDATA_m(3) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(3), 
        CoreAPB3_0_APBmslave0_PRDATA_m(2) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(2), 
        CoreAPB3_0_APBmslave0_PRDATA_m(1) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(1), 
        CoreAPB3_0_APBmslave0_PRDATA_m(0) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(0), 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(15) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[15]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(14) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[14]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(13) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[13]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(12) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[12]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(11) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[11]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(10) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[10]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(9) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[9]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(8) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[8]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(7) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[7]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(6) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[6]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(5) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[5]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(4) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[4]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(3) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[3]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(2) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[2]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(1) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[1]\, 
        MAC_MII_TXD_c(3) => MAC_MII_TXD_c(3), MAC_MII_TXD_c(2)
         => MAC_MII_TXD_c(2), MAC_MII_TXD_c(1) => 
        MAC_MII_TXD_c(1), MAC_MII_TXD_c(0) => MAC_MII_TXD_c(0), 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(16) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[16]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(15) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[15]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(14) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[14]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(13) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[13]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(12) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[12]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(11) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[11]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(10) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[10]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(9) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[9]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(8) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[8]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(7) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[7]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(6) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[6]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(5) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[5]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(4) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[4]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(3) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[3]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(2) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[2]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(1) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[1]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(0) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[0]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(15) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[15]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(14) => nc2, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(13) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[13]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(12) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[12]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(11) => nc4, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(10) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[10]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(9) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[9]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(8) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[8]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(7) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[7]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(6) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[6]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(5) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[5]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[4]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[3]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[2]\, 
        CoreAPB3_0_APBmslave0_PWDATA(7) => 
        CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(15) => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(15), 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(14) => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(14), 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(13) => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(13), 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(12) => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(12), 
        CoreAPB3_0_APBmslave0_PADDR(7) => 
        CoreAPB3_0_APBmslave0_PADDR(7), 
        CoreAPB3_0_APBmslave0_PADDR(6) => 
        CoreAPB3_0_APBmslave0_PADDR(6), 
        CoreAPB3_0_APBmslave0_PADDR(5) => 
        CoreAPB3_0_APBmslave0_PADDR(5), 
        CoreAPB3_0_APBmslave0_PADDR(4) => 
        CoreAPB3_0_APBmslave0_PADDR(4), 
        CoreAPB3_0_APBmslave0_PADDR(3) => 
        CoreAPB3_0_APBmslave0_PADDR(3), 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        CoreAPB3_0_APBmslave0_PADDR(2), 
        CoreAPB3_0_APBmslave0_PADDR(1) => 
        CoreAPB3_0_APBmslave0_PADDR(1), 
        CoreAPB3_0_APBmslave0_PADDR(0) => 
        CoreAPB3_0_APBmslave0_PADDR(0), MDDR_ADDR(15) => 
        MDDR_ADDR(15), MDDR_ADDR(14) => MDDR_ADDR(14), 
        MDDR_ADDR(13) => MDDR_ADDR(13), MDDR_ADDR(12) => 
        MDDR_ADDR(12), MDDR_ADDR(11) => MDDR_ADDR(11), 
        MDDR_ADDR(10) => MDDR_ADDR(10), MDDR_ADDR(9) => 
        MDDR_ADDR(9), MDDR_ADDR(8) => MDDR_ADDR(8), MDDR_ADDR(7)
         => MDDR_ADDR(7), MDDR_ADDR(6) => MDDR_ADDR(6), 
        MDDR_ADDR(5) => MDDR_ADDR(5), MDDR_ADDR(4) => 
        MDDR_ADDR(4), MDDR_ADDR(3) => MDDR_ADDR(3), MDDR_ADDR(2)
         => MDDR_ADDR(2), MDDR_ADDR(1) => MDDR_ADDR(1), 
        MDDR_ADDR(0) => MDDR_ADDR(0), MDDR_BA(2) => MDDR_BA(2), 
        MDDR_BA(1) => MDDR_BA(1), MDDR_BA(0) => MDDR_BA(0), 
        MDDR_DM_RDQS(1) => MDDR_DM_RDQS(1), MDDR_DM_RDQS(0) => 
        MDDR_DM_RDQS(0), MDDR_DQ(15) => MDDR_DQ(15), MDDR_DQ(14)
         => MDDR_DQ(14), MDDR_DQ(13) => MDDR_DQ(13), MDDR_DQ(12)
         => MDDR_DQ(12), MDDR_DQ(11) => MDDR_DQ(11), MDDR_DQ(10)
         => MDDR_DQ(10), MDDR_DQ(9) => MDDR_DQ(9), MDDR_DQ(8) => 
        MDDR_DQ(8), MDDR_DQ(7) => MDDR_DQ(7), MDDR_DQ(6) => 
        MDDR_DQ(6), MDDR_DQ(5) => MDDR_DQ(5), MDDR_DQ(4) => 
        MDDR_DQ(4), MDDR_DQ(3) => MDDR_DQ(3), MDDR_DQ(2) => 
        MDDR_DQ(2), MDDR_DQ(1) => MDDR_DQ(1), MDDR_DQ(0) => 
        MDDR_DQ(0), MDDR_DQS(1) => MDDR_DQS(1), MDDR_DQS(0) => 
        MDDR_DQS(0), CAM_SPI_1_CLK_Y_0 => \CAM_SPI_1_CLK_Y[0]\, 
        GPIO_7_Y_0 => \GPIO_7_Y[0]\, GPIO_6_Y_0 => \GPIO_6_Y[0]\, 
        DEBOUNCE_OUT_net_0_0 => DEBOUNCE_OUT_net_0_0, GPIO_1_in_0
         => \GPIO_1_in[0]\, state_0 => \state[1]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA_reto_0 => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA_reto[0]\, MDDR_CLK
         => MDDR_CLK, MDDR_CLK_N => MDDR_CLK_N, 
        CORECONFIGP_0_MDDR_APBmslave_PWRITE => 
        CORECONFIGP_0_MDDR_APBmslave_PWRITE, 
        CORECONFIGP_0_MDDR_APBmslave_PSELx => 
        CORECONFIGP_0_MDDR_APBmslave_PSELx, 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE => 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE, 
        m2s010_som_sb_0_CCC_71MHz => \m2s010_som_sb_0_CCC_71MHz\, 
        MAC_MII_TX_CLK_c => MAC_MII_TX_CLK_c, SPI_1_SS0_MX_Y => 
        SPI_1_SS0_MX_Y, SPI_1_DI => SPI_1_DI, MAC_MII_RX_ER_c => 
        MAC_MII_RX_ER_c, MAC_MII_RX_DV_c => MAC_MII_RX_DV_c, 
        MAC_MII_RX_CLK_c => MAC_MII_RX_CLK_c, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY, 
        MMUART_0_RXD_F2M_c => MMUART_0_RXD_F2M_c, 
        DEBOUNCE_OUT_2_c => DEBOUNCE_OUT_2_c, DEBOUNCE_OUT_1_c
         => DEBOUNCE_OUT_1_c, BIBUF_0_Y => BIBUF_0_Y, 
        FAB_CCC_LOCK => FAB_CCC_LOCK, 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i => 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i, CommsFPGA_top_0_INT
         => CommsFPGA_top_0_INT, MAC_MII_CRS_c => MAC_MII_CRS_c, 
        MAC_MII_COL_c => MAC_MII_COL_c, 
        CORECONFIGP_0_MDDR_APBmslave_PSLVERR => 
        CORECONFIGP_0_MDDR_APBmslave_PSLVERR, 
        CORECONFIGP_0_MDDR_APBmslave_PREADY => 
        CORECONFIGP_0_MDDR_APBmslave_PREADY, MAC_MII_TX_EN_c => 
        MAC_MII_TX_EN_c, m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE, 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F, SPI_1_DO_CAM_c => 
        SPI_1_DO_CAM_c, GPIO_11_M2F_c => GPIO_11_M2F_c, 
        m2s010_som_sb_MSS_0_SPI_1_CLK_M2F => 
        m2s010_som_sb_MSS_0_SPI_1_CLK_M2F, GPIO_8_M2F_c => 
        GPIO_8_M2F_c, m2s010_som_sb_MSS_0_GPIO_7_M2F => 
        m2s010_som_sb_MSS_0_GPIO_7_M2F, 
        m2s010_som_sb_MSS_0_GPIO_7_M2F_OE => 
        m2s010_som_sb_MSS_0_GPIO_7_M2F_OE, 
        m2s010_som_sb_MSS_0_GPIO_6_M2F => 
        m2s010_som_sb_MSS_0_GPIO_6_M2F, 
        m2s010_som_sb_MSS_0_GPIO_6_M2F_OE => 
        m2s010_som_sb_MSS_0_GPIO_6_M2F_OE, GPIO_5_M2F_c => 
        GPIO_5_M2F_c, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE, 
        GPIO_24_M2F_c => GPIO_24_M2F_c, MMUART_0_TXD_M2F_c => 
        MMUART_0_TXD_M2F_c, m2s010_som_sb_0_GPIO_28_SW_RESET => 
        m2s010_som_sb_0_GPIO_28_SW_RESET, GPIO_21_M2F_c => 
        GPIO_21_M2F_c, GPIO_22_M2F_c => GPIO_22_M2F_c, 
        m2s010_som_sb_MSS_0_MAC_MII_MDO => 
        m2s010_som_sb_MSS_0_MAC_MII_MDO, 
        m2s010_som_sb_MSS_0_MAC_MII_MDO_EN => 
        m2s010_som_sb_MSS_0_MAC_MII_MDO_EN, MAC_MII_MDC_c => 
        MAC_MII_MDC_c, GPIO_1_M2F => GPIO_1_M2F, 
        m2s010_som_sb_MSS_0_GPIO_1_M2F_OE => 
        m2s010_som_sb_MSS_0_GPIO_1_M2F_OE, 
        m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F => 
        m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        CoreAPB3_0_APBmslave0_PWRITE => 
        CoreAPB3_0_APBmslave0_PWRITE, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx, 
        CoreAPB3_0_APBmslave0_PENABLE => 
        CoreAPB3_0_APBmslave0_PENABLE, GPIO_0_BI => GPIO_0_BI, 
        GPIO_3_BI => GPIO_3_BI, GPIO_4_BI => GPIO_4_BI, 
        GPIO_12_BI => GPIO_12_BI, GPIO_14_BI => GPIO_14_BI, 
        GPIO_15_BI => GPIO_15_BI, GPIO_16_BI => GPIO_16_BI, 
        GPIO_17_BI => GPIO_17_BI, GPIO_18_BI => GPIO_18_BI, 
        GPIO_20_OUT => GPIO_20_OUT, GPIO_25_BI => GPIO_25_BI, 
        GPIO_26_BI => GPIO_26_BI, GPIO_31_BI => GPIO_31_BI, 
        I2C_1_SCL => I2C_1_SCL, I2C_1_SDA => I2C_1_SDA, 
        MDDR_CAS_N => MDDR_CAS_N, MDDR_CKE => MDDR_CKE, MDDR_CS_N
         => MDDR_CS_N, MDDR_DQS_TMATCH_0_IN => 
        MDDR_DQS_TMATCH_0_IN, MDDR_DQS_TMATCH_0_OUT => 
        MDDR_DQS_TMATCH_0_OUT, MDDR_ODT => MDDR_ODT, MDDR_RAS_N
         => MDDR_RAS_N, MDDR_RESET_N => MDDR_RESET_N, MDDR_WE_N
         => MDDR_WE_N, MMUART_1_RXD => MMUART_1_RXD, MMUART_1_TXD
         => MMUART_1_TXD, SPI_0_CLK => SPI_0_CLK, SPI_0_DI => 
        SPI_0_DI, SPI_0_DO => SPI_0_DO, SPI_0_SS0 => SPI_0_SS0, 
        SPI_0_SS1 => SPI_0_SS1, CORECONFIGP_0_APB_S_PCLK_i => 
        CORECONFIGP_0_APB_S_PCLK_i, CORECONFIGP_0_APB_S_PRESET_N
         => CORECONFIGP_0_APB_S_PRESET_N, 
        CORECONFIGP_0_APB_S_PCLK => CORECONFIGP_0_APB_S_PCLK);
    
    SPI_1_SS0_MX : MX2
      port map(A => \OTH_SPI_1_SS0_Y[0]\, B => 
        \CAM_SPI_1_SS0_Y[0]\, S => CommsFPGA_top_0_CAMERA_NODE, Y
         => SPI_1_SS0_MX_Y);
    
    CORERESETP_0 : CoreResetP
      port map(CORECONFIGP_0_CONFIG2_DONE => 
        CORECONFIGP_0_CONFIG2_DONE, CORECONFIGP_0_CONFIG1_DONE
         => CORECONFIGP_0_CONFIG1_DONE, 
        CORECONFIGP_0_APB_S_PRESET_N => 
        CORECONFIGP_0_APB_S_PRESET_N, 
        m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F => 
        m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        m2s010_som_sb_0_POWER_ON_RESET_N => 
        \m2s010_som_sb_0_POWER_ON_RESET_N\, INIT_DONE => 
        INIT_DONE, FABOSC_0_RCOSC_25_50MHZ_O2F => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, m2s010_som_sb_0_CCC_71MHz
         => \m2s010_som_sb_0_CCC_71MHz\);
    
    SYSRESET_POR : SYSRESET
      port map(POWER_ON_RESET_N => 
        \m2s010_som_sb_0_POWER_ON_RESET_N\, DEVRST_N => DEVRST_N);
    
    BIBUF_0 : BIBUF
      port map(PAD => MAC_MII_MDIO, D => 
        m2s010_som_sb_MSS_0_MAC_MII_MDO, E => 
        m2s010_som_sb_MSS_0_MAC_MII_MDO_EN, Y => BIBUF_0_Y);
    
    SPI_1_D0_OUT : OUTBUF
      port map(D => SPI_1_DO_CAM_c, PAD => SPI_1_DO_OTH);
    
    GPIO_6 : m2s010_som_sb_GPIO_6_IO
      port map(GPIO_6_PAD_0 => GPIO_6_PAD_0, GPIO_6_Y_0 => 
        \GPIO_6_Y[0]\, m2s010_som_sb_MSS_0_GPIO_6_M2F_OE => 
        m2s010_som_sb_MSS_0_GPIO_6_M2F_OE, 
        m2s010_som_sb_MSS_0_GPIO_6_M2F => 
        m2s010_som_sb_MSS_0_GPIO_6_M2F);
    
    CORECONFIGP_0 : CoreConfigP
      port map(CORECONFIGP_0_MDDR_APBmslave_PRDATA(15) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[15]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(14) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[14]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(13) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[13]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(12) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[12]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(11) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[11]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(10) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[10]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(9) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[9]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(8) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[8]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(7) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[7]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(6) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[6]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(5) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[5]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(4) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[4]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(3) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[3]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(2) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[2]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(1) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[1]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(17) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[17]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(16) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[16]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(15) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[15]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(14) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[14]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(13) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[13]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(12) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[12]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(11) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[11]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(10) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[10]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(9) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[9]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(8) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[8]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(7) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[7]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(6) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[6]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(5) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[5]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(4) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[4]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(3) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[3]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(2) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[2]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(1) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[1]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(0) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[0]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(15) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[15]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(14) => nc3, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(13) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[13]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(12) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[12]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(11) => nc1, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(10) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[10]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(9) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[9]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(8) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[8]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(7) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[7]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(6) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[6]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(5) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[5]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[4]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[3]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[2]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(16) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[16]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(15) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[15]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(14) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[14]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(13) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[13]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(12) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[12]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(11) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[11]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(10) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[10]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(9) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[9]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(8) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[8]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(7) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[7]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(6) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[6]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(5) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[5]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(4) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[4]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(3) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[3]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(2) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[2]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(1) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[1]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(0) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[0]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(10) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[10]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(9) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[9]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(8) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[8]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(7) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[7]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(6) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[6]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(5) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[5]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(4) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[4]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(3) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[3]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(2) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[2]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(15) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[15]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(14) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[14]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(13) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[13]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(12) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[12]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(11) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[11]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(10) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[10]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(9) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[9]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(8) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[8]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(7) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[7]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(6) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[6]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(5) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[5]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(4) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[4]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(3) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[3]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(2) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[2]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(1) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[1]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(0) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[0]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA_reto_0 => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA_reto[0]\, state_0
         => \state[1]\, CORECONFIGP_0_MDDR_APBmslave_PSLVERR => 
        CORECONFIGP_0_MDDR_APBmslave_PSLVERR, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE, 
        CORECONFIGP_0_MDDR_APBmslave_PREADY => 
        CORECONFIGP_0_MDDR_APBmslave_PREADY, 
        CORECONFIGP_0_MDDR_APBmslave_PSELx => 
        CORECONFIGP_0_MDDR_APBmslave_PSELx, 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE => 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE, INIT_DONE => 
        INIT_DONE, CORECONFIGP_0_APB_S_PCLK_i => 
        CORECONFIGP_0_APB_S_PCLK_i, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE, 
        CORECONFIGP_0_MDDR_APBmslave_PWRITE => 
        CORECONFIGP_0_MDDR_APBmslave_PWRITE, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY, 
        CORECONFIGP_0_CONFIG2_DONE => CORECONFIGP_0_CONFIG2_DONE, 
        CORECONFIGP_0_CONFIG1_DONE => CORECONFIGP_0_CONFIG1_DONE, 
        CORECONFIGP_0_APB_S_PCLK => CORECONFIGP_0_APB_S_PCLK, 
        CORECONFIGP_0_APB_S_PRESET_N => 
        CORECONFIGP_0_APB_S_PRESET_N);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    CCC_0 : m2s010_som_sb_CCC_0_FCCC
      port map(m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC => 
        m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC, FAB_CCC_LOCK
         => FAB_CCC_LOCK, m2s010_som_sb_0_CCC_71MHz => 
        \m2s010_som_sb_0_CCC_71MHz\);
    
    SPI_1_DI_MX : MX2
      port map(A => SPI_1_DI_OTH_c, B => SPI_1_DI_CAM_c, S => 
        CommsFPGA_top_0_CAMERA_NODE, Y => SPI_1_DI);
    
    OTH_SPI_1_SS0 : m2s010_som_sb_OTH_SPI_1_SS0_IO
      port map(SPI_1_SS0_OTH_0 => SPI_1_SS0_OTH_0, 
        OTH_SPI_1_SS0_Y_0 => \OTH_SPI_1_SS0_Y[0]\, 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE, 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F);
    
    FABOSC_0 : m2s010_som_sb_FABOSC_0_OSC
      port map(XTL => XTL, 
        m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC => 
        m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC, 
        FABOSC_0_RCOSC_25_50MHZ_O2F => 
        FABOSC_0_RCOSC_25_50MHZ_O2F);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity Debounce_1 is

    port( DEBOUNCE_IN_c_0    : in    std_logic;
          un2_apb3_reset     : in    std_logic;
          DEBOUNCE_OUT_2_c   : out   std_logic;
          un2_apb3_reset_set : in    std_logic;
          BIT_CLK            : in    std_logic
        );

end Debounce_1;

architecture DEF_ARCH of Debounce_1 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \debounce_cntr[1]_net_1\, VCC_net_1, N_1068_i_i, 
        un3_debounce_cntr_1_cry_1_S_1, GND_net_1, 
        \debounce_cntr[2]_net_1\, un3_debounce_cntr_1_cry_2_S_1, 
        \debounce_cntr[3]_net_1\, un3_debounce_cntr_1_cry_3_S_1, 
        \debounce_cntrrs[4]\, un3_debounce_in_rs_1, 
        \debounce_cntr[4]\, un3_debounce_in_i, 
        un3_debounce_cntr_1_cry_4_S_1, \debounce_cntrrs[6]\, 
        \debounce_cntr[6]\, un3_debounce_cntr_1_cry_6_S_1, 
        \debounce_cntr[5]\, un3_debounce_cntr_1_cry_5_S_1, 
        \debounce_cntr[7]\, un3_debounce_cntr_1_cry_7_S_1, 
        \debounce_cntrrs[8]\, \debounce_cntr[8]_net_1\, 
        un3_debounce_cntr_1_cry_8_S_1, \debounce_cntrrs[9]\, 
        \debounce_cntr[9]_net_1\, un3_debounce_cntr_1_cry_9_S_1, 
        \debounce_cntr[10]_net_1\, un3_debounce_cntr_1_cry_10_S_1, 
        \debounce_cntr[11]_net_1\, un3_debounce_cntr_1_cry_11_S_1, 
        \debounce_cntr[12]_net_1\, un3_debounce_cntr_1_cry_12_S_1, 
        \debounce_cntr[13]_net_1\, un3_debounce_cntr_1_cry_13_S_1, 
        \debounce_cntrrs[14]\, \debounce_cntr[14]_net_1\, 
        un3_debounce_cntr_1_cry_14_S_1, \debounce_cntrrs[15]\, 
        \debounce_cntr[15]_net_1\, un3_debounce_cntr_1_s_15_S_1, 
        \debounce_cntr[0]_net_1\, \debounce_cntr_4[0]_net_1\, 
        DEBOUNCE_OUT_2_crs, un1_debounce_cntr, 
        un3_debounce_cntr_1_s_1_394_FCO, 
        \un3_debounce_cntr_1_cry_1\, \un3_debounce_cntr_1_cry_2\, 
        \un3_debounce_cntr_1_cry_3\, \un3_debounce_cntr_1_cry_4\, 
        \un3_debounce_cntr_1_cry_5\, \un3_debounce_cntr_1_cry_6\, 
        \un3_debounce_cntr_1_cry_7\, \un3_debounce_cntr_1_cry_8\, 
        \un3_debounce_cntr_1_cry_9\, \un3_debounce_cntr_1_cry_10\, 
        \un3_debounce_cntr_1_cry_11\, 
        \un3_debounce_cntr_1_cry_12\, 
        \un3_debounce_cntr_1_cry_13\, 
        \un3_debounce_cntr_1_cry_14\, un1_debounce_cntr_11, 
        un1_debounce_cntr_10, un1_debounce_cntr_9, 
        un1_debounce_cntr_8 : std_logic;

begin 


    \debounce_cntr_0_0[0]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_5_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => N_1068_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \debounce_cntr[5]\);
    
    un3_debounce_cntr_1_cry_9 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[9]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_8\, S => 
        un3_debounce_cntr_1_cry_9_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_9\);
    
    \debounce_cntr[12]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_12_S_1, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => N_1068_i_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[12]_net_1\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_8\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \debounce_cntr[2]_net_1\, B => 
        \debounce_cntr[1]_net_1\, C => \debounce_cntr[15]_net_1\, 
        D => \debounce_cntr[14]_net_1\, Y => un1_debounce_cntr_8);
    
    \DEBOUNCE_PROC.un3_debounce_in_rs\ : SLE
      port map(D => VCC_net_1, CLK => un2_apb3_reset, EN => 
        VCC_net_1, ALn => un3_debounce_in_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q
         => un3_debounce_in_rs_1);
    
    \debounce_cntr[15]\ : SLE
      port map(D => un3_debounce_cntr_1_s_15_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[15]\);
    
    un3_debounce_cntr_1_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_4\, S => 
        un3_debounce_cntr_1_cry_5_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_5\);
    
    un3_debounce_cntr_1_cry_2 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[2]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_1\, S => 
        un3_debounce_cntr_1_cry_2_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_2\);
    
    \debounce_cntr[3]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_3_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => N_1068_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \debounce_cntr[3]_net_1\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_9\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \debounce_cntr[9]_net_1\, B => 
        \debounce_cntr[8]_net_1\, C => \debounce_cntr[6]\, D => 
        \debounce_cntr[4]\, Y => un1_debounce_cntr_9);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_10\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \debounce_cntr[13]_net_1\, B => 
        \debounce_cntr[12]_net_1\, C => \debounce_cntr[11]_net_1\, 
        D => \debounce_cntr[10]_net_1\, Y => un1_debounce_cntr_10);
    
    debounce_out : SLE
      port map(D => un1_debounce_cntr, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => un3_debounce_in_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => DEBOUNCE_OUT_2_crs);
    
    \debounce_cntr_RNI9QDE[9]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \debounce_cntrrs[9]\, B => 
        un3_debounce_in_rs_1, C => un2_apb3_reset_set, Y => 
        \debounce_cntr[9]_net_1\);
    
    \debounce_cntr[10]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_10_S_1, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => N_1068_i_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[10]_net_1\);
    
    un3_debounce_cntr_1_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_3\, S => 
        un3_debounce_cntr_1_cry_4_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_4\);
    
    \debounce_cntr_RNI8PDE[8]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \debounce_cntrrs[8]\, B => 
        un3_debounce_in_rs_1, C => un2_apb3_reset_set, Y => 
        \debounce_cntr[8]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \debounce_cntr[13]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_13_S_1, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => N_1068_i_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[13]_net_1\);
    
    \debounce_cntr_RNIMRBQ[15]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \debounce_cntrrs[15]\, B => 
        un3_debounce_in_rs_1, C => un2_apb3_reset_set, Y => 
        \debounce_cntr[15]_net_1\);
    
    un3_debounce_cntr_1_cry_14 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[14]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_13\, S => 
        un3_debounce_cntr_1_cry_14_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_14\);
    
    debounce_out_RNIPLAK : CFG3
      generic map(INIT => x"F8")

      port map(A => un3_debounce_in_rs_1, B => un2_apb3_reset_set, 
        C => DEBOUNCE_OUT_2_crs, Y => DEBOUNCE_OUT_2_c);
    
    \debounce_cntr_0_0[1]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_7_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => N_1068_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \debounce_cntr[7]\);
    
    un3_debounce_cntr_1_cry_13 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[13]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_12\, S => 
        un3_debounce_cntr_1_cry_13_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_13\);
    
    \debounce_cntr[9]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_9_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[9]\);
    
    \DEBOUNCE_PROC.un3_debounce_in_0_a3\ : CFG2
      generic map(INIT => x"E")

      port map(A => un2_apb3_reset, B => DEBOUNCE_IN_c_0, Y => 
        un3_debounce_in_i);
    
    un3_debounce_cntr_1_cry_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_6\, S => 
        un3_debounce_cntr_1_cry_7_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_7\);
    
    un3_debounce_cntr_1_s_1_394 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[0]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => 
        OPEN, Y => OPEN, FCO => un3_debounce_cntr_1_s_1_394_FCO);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \debounce_cntr[1]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_1_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => N_1068_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \debounce_cntr[1]_net_1\);
    
    \debounce_cntr_0[0]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_4_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[4]\);
    
    N_1068_i : CFG2
      generic map(INIT => x"4")

      port map(A => un2_apb3_reset, B => DEBOUNCE_IN_c_0, Y => 
        N_1068_i_i);
    
    \debounce_cntr[14]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_14_S_1, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => un3_debounce_in_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[14]\);
    
    un3_debounce_cntr_1_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_5\, S => 
        un3_debounce_cntr_1_cry_6_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_6\);
    
    un3_debounce_cntr_1_cry_11 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[11]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_10\, S => 
        un3_debounce_cntr_1_cry_11_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_11\);
    
    \debounce_cntr_4[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => un1_debounce_cntr, B => 
        \debounce_cntr[0]_net_1\, Y => \debounce_cntr_4[0]_net_1\);
    
    \debounce_cntr_RNILQBQ[14]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \debounce_cntrrs[14]\, B => 
        un3_debounce_in_rs_1, C => un2_apb3_reset_set, Y => 
        \debounce_cntr[14]_net_1\);
    
    \debounce_cntr[8]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_8_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[8]\);
    
    \debounce_cntr[0]\ : SLE
      port map(D => \debounce_cntr_4[0]_net_1\, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => N_1068_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \debounce_cntr[0]_net_1\);
    
    \debounce_cntr_0[1]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_6_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[6]\);
    
    un3_debounce_cntr_1_cry_8 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[8]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_7\, S => 
        un3_debounce_cntr_1_cry_8_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_8\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr\ : CFG4
      generic map(INIT => x"8000")

      port map(A => un1_debounce_cntr_11, B => 
        un1_debounce_cntr_10, C => un1_debounce_cntr_8, D => 
        un1_debounce_cntr_9, Y => un1_debounce_cntr);
    
    un3_debounce_cntr_1_cry_12 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[12]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_11\, S => 
        un3_debounce_cntr_1_cry_12_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_12\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_11\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \debounce_cntr[7]\, B => \debounce_cntr[5]\, 
        C => \debounce_cntr[3]_net_1\, D => 
        \debounce_cntr[0]_net_1\, Y => un1_debounce_cntr_11);
    
    un3_debounce_cntr_1_s_15 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[15]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_14\, S => 
        un3_debounce_cntr_1_s_15_S_1, Y => OPEN, FCO => OPEN);
    
    un3_debounce_cntr_1_cry_10 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[10]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_9\, S => 
        un3_debounce_cntr_1_cry_10_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_10\);
    
    \debounce_cntr_0_RNIGGHL[1]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \debounce_cntrrs[6]\, B => 
        un3_debounce_in_rs_1, C => un2_apb3_reset_set, Y => 
        \debounce_cntr[6]\);
    
    \debounce_cntr[2]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_2_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => N_1068_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \debounce_cntr[2]_net_1\);
    
    \debounce_cntr[11]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_11_S_1, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => N_1068_i_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[11]_net_1\);
    
    \debounce_cntr_0_RNIFFHL[0]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \debounce_cntrrs[4]\, B => 
        un3_debounce_in_rs_1, C => un2_apb3_reset_set, Y => 
        \debounce_cntr[4]\);
    
    un3_debounce_cntr_1_cry_1 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[1]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        un3_debounce_cntr_1_s_1_394_FCO, S => 
        un3_debounce_cntr_1_cry_1_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_1\);
    
    un3_debounce_cntr_1_cry_3 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[3]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_2\, S => 
        un3_debounce_cntr_1_cry_3_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_3\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity Debounce_0 is

    port( DEBOUNCE_IN_c_0    : in    std_logic;
          un2_apb3_reset     : in    std_logic;
          DEBOUNCE_OUT_1_c   : out   std_logic;
          un2_apb3_reset_set : in    std_logic;
          BIT_CLK            : in    std_logic
        );

end Debounce_0;

architecture DEF_ARCH of Debounce_0 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \debounce_cntr[1]_net_1\, VCC_net_1, N_1053_i_i, 
        un3_debounce_cntr_1_cry_1_S_0, GND_net_1, 
        \debounce_cntr[2]_net_1\, un3_debounce_cntr_1_cry_2_S_0, 
        \debounce_cntr[3]_net_1\, un3_debounce_cntr_1_cry_3_S_0, 
        \debounce_cntrrs[4]\, un3_debounce_in_rs_0, 
        \debounce_cntr[4]\, un3_debounce_in_i, 
        un3_debounce_cntr_1_cry_4_S_0, \debounce_cntrrs[6]\, 
        \debounce_cntr[6]\, un3_debounce_cntr_1_cry_6_S_0, 
        \debounce_cntr[5]\, un3_debounce_cntr_1_cry_5_S_0, 
        \debounce_cntr[7]\, un3_debounce_cntr_1_cry_7_S_0, 
        \debounce_cntrrs[8]\, \debounce_cntr[8]_net_1\, 
        un3_debounce_cntr_1_cry_8_S_0, \debounce_cntrrs[9]\, 
        \debounce_cntr[9]_net_1\, un3_debounce_cntr_1_cry_9_S_0, 
        \debounce_cntr[10]_net_1\, un3_debounce_cntr_1_cry_10_S_0, 
        \debounce_cntr[11]_net_1\, un3_debounce_cntr_1_cry_11_S_0, 
        \debounce_cntr[12]_net_1\, un3_debounce_cntr_1_cry_12_S_0, 
        \debounce_cntr[13]_net_1\, un3_debounce_cntr_1_cry_13_S_0, 
        \debounce_cntrrs[14]\, \debounce_cntr[14]_net_1\, 
        un3_debounce_cntr_1_cry_14_S_0, \debounce_cntrrs[15]\, 
        \debounce_cntr[15]_net_1\, un3_debounce_cntr_1_s_15_S_0, 
        \debounce_cntr[0]_net_1\, \debounce_cntr_4[0]_net_1\, 
        DEBOUNCE_OUT_1_crs, un1_debounce_cntr, 
        un3_debounce_cntr_1_s_1_393_FCO, 
        \un3_debounce_cntr_1_cry_1\, \un3_debounce_cntr_1_cry_2\, 
        \un3_debounce_cntr_1_cry_3\, \un3_debounce_cntr_1_cry_4\, 
        \un3_debounce_cntr_1_cry_5\, \un3_debounce_cntr_1_cry_6\, 
        \un3_debounce_cntr_1_cry_7\, \un3_debounce_cntr_1_cry_8\, 
        \un3_debounce_cntr_1_cry_9\, \un3_debounce_cntr_1_cry_10\, 
        \un3_debounce_cntr_1_cry_11\, 
        \un3_debounce_cntr_1_cry_12\, 
        \un3_debounce_cntr_1_cry_13\, 
        \un3_debounce_cntr_1_cry_14\, un1_debounce_cntr_11, 
        un1_debounce_cntr_10, un1_debounce_cntr_9, 
        un1_debounce_cntr_8 : std_logic;

begin 


    \debounce_cntr_0_0[0]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_5_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => N_1053_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \debounce_cntr[5]\);
    
    un3_debounce_cntr_1_cry_9 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[9]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_8\, S => 
        un3_debounce_cntr_1_cry_9_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_9\);
    
    \debounce_cntr[12]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_12_S_0, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => N_1053_i_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[12]_net_1\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_8\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \debounce_cntr[2]_net_1\, B => 
        \debounce_cntr[1]_net_1\, C => \debounce_cntr[15]_net_1\, 
        D => \debounce_cntr[14]_net_1\, Y => un1_debounce_cntr_8);
    
    \DEBOUNCE_PROC.un3_debounce_in_rs\ : SLE
      port map(D => VCC_net_1, CLK => un2_apb3_reset, EN => 
        VCC_net_1, ALn => un3_debounce_in_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q
         => un3_debounce_in_rs_0);
    
    \debounce_cntr[15]\ : SLE
      port map(D => un3_debounce_cntr_1_s_15_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[15]\);
    
    un3_debounce_cntr_1_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_4\, S => 
        un3_debounce_cntr_1_cry_5_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_5\);
    
    un3_debounce_cntr_1_cry_2 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[2]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_1\, S => 
        un3_debounce_cntr_1_cry_2_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_2\);
    
    \debounce_cntr[3]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_3_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => N_1053_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \debounce_cntr[3]_net_1\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_9\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \debounce_cntr[9]_net_1\, B => 
        \debounce_cntr[8]_net_1\, C => \debounce_cntr[6]\, D => 
        \debounce_cntr[4]\, Y => un1_debounce_cntr_9);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_10\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \debounce_cntr[13]_net_1\, B => 
        \debounce_cntr[12]_net_1\, C => \debounce_cntr[11]_net_1\, 
        D => \debounce_cntr[10]_net_1\, Y => un1_debounce_cntr_10);
    
    debounce_out : SLE
      port map(D => un1_debounce_cntr, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => un3_debounce_in_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => DEBOUNCE_OUT_1_crs);
    
    \debounce_cntr[10]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_10_S_0, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => N_1053_i_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[10]_net_1\);
    
    un3_debounce_cntr_1_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_3\, S => 
        un3_debounce_cntr_1_cry_4_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_4\);
    
    debounce_out_RNINTGL : CFG3
      generic map(INIT => x"EA")

      port map(A => DEBOUNCE_OUT_1_crs, B => un3_debounce_in_rs_0, 
        C => un2_apb3_reset_set, Y => DEBOUNCE_OUT_1_c);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \debounce_cntr_RNI7U5P[9]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un2_apb3_reset_set, B => \debounce_cntrrs[9]\, 
        C => un3_debounce_in_rs_0, Y => \debounce_cntr[9]_net_1\);
    
    \debounce_cntr[13]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_13_S_0, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => N_1053_i_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[13]_net_1\);
    
    un3_debounce_cntr_1_cry_14 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[14]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_13\, S => 
        un3_debounce_cntr_1_cry_14_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_14\);
    
    \debounce_cntr_0_0[1]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_7_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => N_1053_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \debounce_cntr[7]\);
    
    un3_debounce_cntr_1_cry_13 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[13]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_12\, S => 
        un3_debounce_cntr_1_cry_13_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_13\);
    
    \debounce_cntr[9]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_9_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[9]\);
    
    \DEBOUNCE_PROC.un3_debounce_in_0_a3\ : CFG2
      generic map(INIT => x"E")

      port map(A => un2_apb3_reset, B => DEBOUNCE_IN_c_0, Y => 
        un3_debounce_in_i);
    
    \debounce_cntr_RNIKUDT[15]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un2_apb3_reset_set, B => 
        \debounce_cntrrs[15]\, C => un3_debounce_in_rs_0, Y => 
        \debounce_cntr[15]_net_1\);
    
    un3_debounce_cntr_1_cry_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_6\, S => 
        un3_debounce_cntr_1_cry_7_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_7\);
    
    \debounce_cntr_0_RNIEISQ[1]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un2_apb3_reset_set, B => \debounce_cntrrs[6]\, 
        C => un3_debounce_in_rs_0, Y => \debounce_cntr[6]\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \debounce_cntr_RNI6T5P[8]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un2_apb3_reset_set, B => \debounce_cntrrs[8]\, 
        C => un3_debounce_in_rs_0, Y => \debounce_cntr[8]_net_1\);
    
    \debounce_cntr[1]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_1_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => N_1053_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \debounce_cntr[1]_net_1\);
    
    \debounce_cntr_0[0]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_4_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[4]\);
    
    \debounce_cntr[14]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_14_S_0, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => un3_debounce_in_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[14]\);
    
    un3_debounce_cntr_1_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_5\, S => 
        un3_debounce_cntr_1_cry_6_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_6\);
    
    N_1053_i : CFG2
      generic map(INIT => x"4")

      port map(A => un2_apb3_reset, B => DEBOUNCE_IN_c_0, Y => 
        N_1053_i_i);
    
    un3_debounce_cntr_1_cry_11 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[11]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_10\, S => 
        un3_debounce_cntr_1_cry_11_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_11\);
    
    \debounce_cntr_4[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => un1_debounce_cntr, B => 
        \debounce_cntr[0]_net_1\, Y => \debounce_cntr_4[0]_net_1\);
    
    \debounce_cntr[8]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_8_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[8]\);
    
    \debounce_cntr[0]\ : SLE
      port map(D => \debounce_cntr_4[0]_net_1\, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => N_1053_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \debounce_cntr[0]_net_1\);
    
    \debounce_cntr_0[1]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_6_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[6]\);
    
    un3_debounce_cntr_1_cry_8 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[8]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_7\, S => 
        un3_debounce_cntr_1_cry_8_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_8\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr\ : CFG4
      generic map(INIT => x"8000")

      port map(A => un1_debounce_cntr_11, B => 
        un1_debounce_cntr_10, C => un1_debounce_cntr_8, D => 
        un1_debounce_cntr_9, Y => un1_debounce_cntr);
    
    un3_debounce_cntr_1_cry_12 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[12]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_11\, S => 
        un3_debounce_cntr_1_cry_12_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_12\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_11\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \debounce_cntr[7]\, B => \debounce_cntr[5]\, 
        C => \debounce_cntr[3]_net_1\, D => 
        \debounce_cntr[0]_net_1\, Y => un1_debounce_cntr_11);
    
    un3_debounce_cntr_1_s_15 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[15]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_14\, S => 
        un3_debounce_cntr_1_s_15_S_0, Y => OPEN, FCO => OPEN);
    
    un3_debounce_cntr_1_cry_10 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[10]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_9\, S => 
        un3_debounce_cntr_1_cry_10_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_10\);
    
    \debounce_cntr_RNIJTDT[14]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un2_apb3_reset_set, B => 
        \debounce_cntrrs[14]\, C => un3_debounce_in_rs_0, Y => 
        \debounce_cntr[14]_net_1\);
    
    \debounce_cntr_0_RNIDHSQ[0]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un2_apb3_reset_set, B => \debounce_cntrrs[4]\, 
        C => un3_debounce_in_rs_0, Y => \debounce_cntr[4]\);
    
    \debounce_cntr[2]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_2_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => N_1053_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \debounce_cntr[2]_net_1\);
    
    \debounce_cntr[11]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_11_S_0, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => N_1053_i_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[11]_net_1\);
    
    un3_debounce_cntr_1_cry_1 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[1]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        un3_debounce_cntr_1_s_1_393_FCO, S => 
        un3_debounce_cntr_1_cry_1_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_1\);
    
    un3_debounce_cntr_1_cry_3 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[3]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_2\, S => 
        un3_debounce_cntr_1_cry_3_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_3\);
    
    un3_debounce_cntr_1_s_1_393 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[0]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => 
        OPEN, Y => OPEN, FCO => un3_debounce_cntr_1_s_1_393_FCO);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity Debounce is

    port( DEBOUNCE_IN_c_0      : in    std_logic;
          DEBOUNCE_OUT_net_0_0 : out   std_logic;
          un2_apb3_reset       : in    std_logic;
          un2_apb3_reset_set   : in    std_logic;
          BIT_CLK              : in    std_logic
        );

end Debounce;

architecture DEF_ARCH of Debounce is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \debounce_cntr[1]_net_1\, VCC_net_1, N_1052_i_i, 
        un3_debounce_cntr_1_cry_1_S, GND_net_1, 
        \debounce_cntr[2]_net_1\, un3_debounce_cntr_1_cry_2_S, 
        \debounce_cntr[3]_net_1\, un3_debounce_cntr_1_cry_3_S, 
        \debounce_cntrrs[4]\, un3_debounce_in_rs, 
        \debounce_cntr[4]\, un3_debounce_in_i, 
        un3_debounce_cntr_1_cry_4_S, \debounce_cntrrs[6]\, 
        \debounce_cntr[6]\, un3_debounce_cntr_1_cry_6_S, 
        \debounce_cntr[5]\, un3_debounce_cntr_1_cry_5_S, 
        \debounce_cntr[7]\, un3_debounce_cntr_1_cry_7_S, 
        \debounce_cntrrs[8]\, \debounce_cntr[8]_net_1\, 
        un3_debounce_cntr_1_cry_8_S, \debounce_cntrrs[9]\, 
        \debounce_cntr[9]_net_1\, un3_debounce_cntr_1_cry_9_S, 
        \debounce_cntr[10]_net_1\, un3_debounce_cntr_1_cry_10_S, 
        \debounce_cntr[11]_net_1\, un3_debounce_cntr_1_cry_11_S, 
        \debounce_cntr[12]_net_1\, un3_debounce_cntr_1_cry_12_S, 
        \debounce_cntr[13]_net_1\, un3_debounce_cntr_1_cry_13_S, 
        \debounce_cntrrs[14]\, \debounce_cntr[14]_net_1\, 
        un3_debounce_cntr_1_cry_14_S, \debounce_cntrrs[15]\, 
        \debounce_cntr[15]_net_1\, un3_debounce_cntr_1_s_15_S, 
        \debounce_cntr[0]_net_1\, \debounce_cntr_4[0]_net_1\, 
        \DEBOUNCE_OUT_net_0rs[0]\, un1_debounce_cntr, 
        un3_debounce_cntr_1_s_1_392_FCO, 
        \un3_debounce_cntr_1_cry_1\, \un3_debounce_cntr_1_cry_2\, 
        \un3_debounce_cntr_1_cry_3\, \un3_debounce_cntr_1_cry_4\, 
        \un3_debounce_cntr_1_cry_5\, \un3_debounce_cntr_1_cry_6\, 
        \un3_debounce_cntr_1_cry_7\, \un3_debounce_cntr_1_cry_8\, 
        \un3_debounce_cntr_1_cry_9\, \un3_debounce_cntr_1_cry_10\, 
        \un3_debounce_cntr_1_cry_11\, 
        \un3_debounce_cntr_1_cry_12\, 
        \un3_debounce_cntr_1_cry_13\, 
        \un3_debounce_cntr_1_cry_14\, un1_debounce_cntr_11, 
        un1_debounce_cntr_10, un1_debounce_cntr_9, 
        un1_debounce_cntr_8 : std_logic;

begin 


    \debounce_cntr_0_0[0]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_5_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => N_1052_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \debounce_cntr[5]\);
    
    un3_debounce_cntr_1_cry_9 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[9]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_8\, S => 
        un3_debounce_cntr_1_cry_9_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_9\);
    
    \debounce_cntr[12]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_12_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => N_1052_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \debounce_cntr[12]_net_1\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_8\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \debounce_cntr[2]_net_1\, B => 
        \debounce_cntr[1]_net_1\, C => \debounce_cntr[15]_net_1\, 
        D => \debounce_cntr[14]_net_1\, Y => un1_debounce_cntr_8);
    
    \DEBOUNCE_PROC.un3_debounce_in_rs\ : SLE
      port map(D => VCC_net_1, CLK => un2_apb3_reset, EN => 
        VCC_net_1, ALn => un3_debounce_in_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q
         => un3_debounce_in_rs);
    
    \debounce_cntr[15]\ : SLE
      port map(D => un3_debounce_cntr_1_s_15_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[15]\);
    
    un3_debounce_cntr_1_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_4\, S => 
        un3_debounce_cntr_1_cry_5_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_5\);
    
    un3_debounce_cntr_1_cry_2 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[2]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_1\, S => 
        un3_debounce_cntr_1_cry_2_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_2\);
    
    \debounce_cntr[3]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_3_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => N_1052_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \debounce_cntr[3]_net_1\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_9\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \debounce_cntr[9]_net_1\, B => 
        \debounce_cntr[8]_net_1\, C => \debounce_cntr[6]\, D => 
        \debounce_cntr[4]\, Y => un1_debounce_cntr_9);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_10\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \debounce_cntr[13]_net_1\, B => 
        \debounce_cntr[12]_net_1\, C => \debounce_cntr[11]_net_1\, 
        D => \debounce_cntr[10]_net_1\, Y => un1_debounce_cntr_10);
    
    \debounce_cntr_0_RNIBJ7G[0]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un2_apb3_reset_set, B => \debounce_cntrrs[4]\, 
        C => un3_debounce_in_rs, Y => \debounce_cntr[4]\);
    
    debounce_out : SLE
      port map(D => un1_debounce_cntr, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => un3_debounce_in_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \DEBOUNCE_OUT_net_0rs[0]\);
    
    \debounce_cntr[10]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_10_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => N_1052_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \debounce_cntr[10]_net_1\);
    
    un3_debounce_cntr_1_s_1_392 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[0]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => 
        OPEN, Y => OPEN, FCO => un3_debounce_cntr_1_s_1_392_FCO);
    
    un3_debounce_cntr_1_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_3\, S => 
        un3_debounce_cntr_1_cry_4_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_4\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \debounce_cntr[13]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_13_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => N_1052_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \debounce_cntr[13]_net_1\);
    
    un3_debounce_cntr_1_cry_14 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[14]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_13\, S => 
        un3_debounce_cntr_1_cry_14_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_14\);
    
    \debounce_cntr_0_0[1]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_7_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => N_1052_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \debounce_cntr[7]\);
    
    un3_debounce_cntr_1_cry_13 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[13]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_12\, S => 
        un3_debounce_cntr_1_cry_13_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_13\);
    
    \debounce_cntr[9]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_9_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[9]\);
    
    \debounce_cntr_RNI41UJ[8]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un2_apb3_reset_set, B => \debounce_cntrrs[8]\, 
        C => un3_debounce_in_rs, Y => \debounce_cntr[8]_net_1\);
    
    \DEBOUNCE_PROC.un3_debounce_in_0_a3\ : CFG2
      generic map(INIT => x"E")

      port map(A => un2_apb3_reset, B => DEBOUNCE_IN_c_0, Y => 
        un3_debounce_in_i);
    
    un3_debounce_cntr_1_cry_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_6\, S => 
        un3_debounce_cntr_1_cry_7_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_7\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \debounce_cntr[1]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_1_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => N_1052_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \debounce_cntr[1]_net_1\);
    
    \debounce_cntr_0[0]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_4_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[4]\);
    
    \debounce_cntr[14]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_14_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[14]\);
    
    un3_debounce_cntr_1_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_5\, S => 
        un3_debounce_cntr_1_cry_6_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_6\);
    
    un3_debounce_cntr_1_cry_11 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[11]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_10\, S => 
        un3_debounce_cntr_1_cry_11_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_11\);
    
    \debounce_cntr_0_RNICK7G[1]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un2_apb3_reset_set, B => \debounce_cntrrs[6]\, 
        C => un3_debounce_in_rs, Y => \debounce_cntr[6]\);
    
    \debounce_cntr_4[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => un1_debounce_cntr, B => 
        \debounce_cntr[0]_net_1\, Y => \debounce_cntr_4[0]_net_1\);
    
    \debounce_cntr[8]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_8_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[8]\);
    
    \debounce_cntr[0]\ : SLE
      port map(D => \debounce_cntr_4[0]_net_1\, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => N_1052_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \debounce_cntr[0]_net_1\);
    
    \debounce_cntr_0[1]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_6_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[6]\);
    
    N_1052_i : CFG2
      generic map(INIT => x"4")

      port map(A => un2_apb3_reset, B => DEBOUNCE_IN_c_0, Y => 
        N_1052_i_i);
    
    un3_debounce_cntr_1_cry_8 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[8]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_7\, S => 
        un3_debounce_cntr_1_cry_8_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_8\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr\ : CFG4
      generic map(INIT => x"8000")

      port map(A => un1_debounce_cntr_11, B => 
        un1_debounce_cntr_10, C => un1_debounce_cntr_8, D => 
        un1_debounce_cntr_9, Y => un1_debounce_cntr);
    
    un3_debounce_cntr_1_cry_12 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[12]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_11\, S => 
        un3_debounce_cntr_1_cry_12_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_12\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_11\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \debounce_cntr[7]\, B => \debounce_cntr[5]\, 
        C => \debounce_cntr[3]_net_1\, D => 
        \debounce_cntr[0]_net_1\, Y => un1_debounce_cntr_11);
    
    un3_debounce_cntr_1_s_15 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[15]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_14\, S => 
        un3_debounce_cntr_1_s_15_S, Y => OPEN, FCO => OPEN);
    
    un3_debounce_cntr_1_cry_10 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[10]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_9\, S => 
        un3_debounce_cntr_1_cry_10_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_10\);
    
    \debounce_cntr_RNI52UJ[9]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un2_apb3_reset_set, B => \debounce_cntrrs[9]\, 
        C => un3_debounce_in_rs, Y => \debounce_cntr[9]_net_1\);
    
    \debounce_cntr_RNIH0GG[14]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un2_apb3_reset_set, B => 
        \debounce_cntrrs[14]\, C => un3_debounce_in_rs, Y => 
        \debounce_cntr[14]_net_1\);
    
    \debounce_cntr[2]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_2_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => N_1052_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \debounce_cntr[2]_net_1\);
    
    \debounce_cntr[11]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_11_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => N_1052_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \debounce_cntr[11]_net_1\);
    
    un3_debounce_cntr_1_cry_1 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[1]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        un3_debounce_cntr_1_s_1_392_FCO, S => 
        un3_debounce_cntr_1_cry_1_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_1\);
    
    \debounce_cntr_RNII1GG[15]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => un2_apb3_reset_set, B => 
        \debounce_cntrrs[15]\, C => un3_debounce_in_rs, Y => 
        \debounce_cntr[15]_net_1\);
    
    debounce_out_RNIL5NM : CFG3
      generic map(INIT => x"EA")

      port map(A => \DEBOUNCE_OUT_net_0rs[0]\, B => 
        un3_debounce_in_rs, C => un2_apb3_reset_set, Y => 
        DEBOUNCE_OUT_net_0_0);
    
    un3_debounce_cntr_1_cry_3 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[3]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_2\, S => 
        un3_debounce_cntr_1_cry_3_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_3\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity TriDebounce is

    port( DEBOUNCE_IN_c        : in    std_logic_vector(2 downto 0);
          DEBOUNCE_OUT_net_0_0 : out   std_logic;
          DEBOUNCE_OUT_2_c     : out   std_logic;
          DEBOUNCE_OUT_1_c     : out   std_logic;
          BIT_CLK              : in    std_logic;
          un2_apb3_reset_set   : in    std_logic;
          un2_apb3_reset       : in    std_logic
        );

end TriDebounce;

architecture DEF_ARCH of TriDebounce is 

  component Debounce_1
    port( DEBOUNCE_IN_c_0    : in    std_logic := 'U';
          un2_apb3_reset     : in    std_logic := 'U';
          DEBOUNCE_OUT_2_c   : out   std_logic;
          un2_apb3_reset_set : in    std_logic := 'U';
          BIT_CLK            : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component Debounce_0
    port( DEBOUNCE_IN_c_0    : in    std_logic := 'U';
          un2_apb3_reset     : in    std_logic := 'U';
          DEBOUNCE_OUT_1_c   : out   std_logic;
          un2_apb3_reset_set : in    std_logic := 'U';
          BIT_CLK            : in    std_logic := 'U'
        );
  end component;

  component Debounce
    port( DEBOUNCE_IN_c_0      : in    std_logic := 'U';
          DEBOUNCE_OUT_net_0_0 : out   std_logic;
          un2_apb3_reset       : in    std_logic := 'U';
          un2_apb3_reset_set   : in    std_logic := 'U';
          BIT_CLK              : in    std_logic := 'U'
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : Debounce_1
	Use entity work.Debounce_1(DEF_ARCH);
    for all : Debounce_0
	Use entity work.Debounce_0(DEF_ARCH);
    for all : Debounce
	Use entity work.Debounce(DEF_ARCH);
begin 


    DEBOUNCE_2_INST : Debounce_1
      port map(DEBOUNCE_IN_c_0 => DEBOUNCE_IN_c(2), 
        un2_apb3_reset => un2_apb3_reset, DEBOUNCE_OUT_2_c => 
        DEBOUNCE_OUT_2_c, un2_apb3_reset_set => 
        un2_apb3_reset_set, BIT_CLK => BIT_CLK);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    DEBOUNCE_1_INST : Debounce_0
      port map(DEBOUNCE_IN_c_0 => DEBOUNCE_IN_c(1), 
        un2_apb3_reset => un2_apb3_reset, DEBOUNCE_OUT_1_c => 
        DEBOUNCE_OUT_1_c, un2_apb3_reset_set => 
        un2_apb3_reset_set, BIT_CLK => BIT_CLK);
    
    DEBOUNCE_0_INST : Debounce
      port map(DEBOUNCE_IN_c_0 => DEBOUNCE_IN_c(0), 
        DEBOUNCE_OUT_net_0_0 => DEBOUNCE_OUT_net_0_0, 
        un2_apb3_reset => un2_apb3_reset, un2_apb3_reset_set => 
        un2_apb3_reset_set, BIT_CLK => BIT_CLK);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CRC16_Generator_0 is

    port( tx_crc_data    : out   std_logic_vector(15 downto 0);
          N_705          : in    std_logic;
          N_709          : in    std_logic;
          N_710          : in    std_logic;
          N_711          : in    std_logic;
          N_704          : in    std_logic;
          N_707          : in    std_logic;
          N_708          : in    std_logic;
          N_706          : in    std_logic;
          tx_crc_gen     : in    std_logic;
          byte_clk_en    : in    std_logic;
          BIT_CLK        : in    std_logic;
          tx_crc_reset_i : in    std_logic
        );

end CRC16_Generator_0;

architecture DEF_ARCH of CRC16_Generator_0 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \tx_crc_data[13]\, GND_net_1, \tx_crc_data[5]\, 
        \lfsr_q_0_sqmuxa\, VCC_net_1, \tx_crc_data[14]\, 
        \tx_crc_data[6]\, \tx_crc_data[15]\, \lfsr_c[15]\, 
        \tx_crc_data[0]\, \lfsr_c[0]\, \tx_crc_data[1]\, 
        \lfsr_c[1]\, \tx_crc_data[2]\, N_617_i, \tx_crc_data[3]\, 
        N_620_i, \tx_crc_data[4]\, N_619_i, N_618_i, N_621_i, 
        \tx_crc_data[7]\, N_622_i, \tx_crc_data[8]\, N_107_i_i, 
        \tx_crc_data[9]\, \lfsr_c[9]\, \tx_crc_data[10]\, 
        \tx_crc_data[11]\, \tx_crc_data[12]\, N_567_i
         : std_logic;

begin 

    tx_crc_data(15) <= \tx_crc_data[15]\;
    tx_crc_data(14) <= \tx_crc_data[14]\;
    tx_crc_data(13) <= \tx_crc_data[13]\;
    tx_crc_data(12) <= \tx_crc_data[12]\;
    tx_crc_data(11) <= \tx_crc_data[11]\;
    tx_crc_data(10) <= \tx_crc_data[10]\;
    tx_crc_data(9) <= \tx_crc_data[9]\;
    tx_crc_data(8) <= \tx_crc_data[8]\;
    tx_crc_data(7) <= \tx_crc_data[7]\;
    tx_crc_data(6) <= \tx_crc_data[6]\;
    tx_crc_data(5) <= \tx_crc_data[5]\;
    tx_crc_data(4) <= \tx_crc_data[4]\;
    tx_crc_data(3) <= \tx_crc_data[3]\;
    tx_crc_data(2) <= \tx_crc_data[2]\;
    tx_crc_data(1) <= \tx_crc_data[1]\;
    tx_crc_data(0) <= \tx_crc_data[0]\;

    \lfsr_q[9]\ : SLE
      port map(D => \lfsr_c[9]\, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[9]\);
    
    \lfsr_q[6]\ : SLE
      port map(D => N_621_i, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[6]\);
    
    \lfsr_q[3]\ : SLE
      port map(D => N_620_i, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[3]\);
    
    \lfsr_c_0_a2_0_x2_0_x2_0_x2[3]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \tx_crc_data[10]\, B => \tx_crc_data[9]\, C
         => N_711, D => N_710, Y => N_620_i);
    
    \lfsr_q[10]\ : SLE
      port map(D => \tx_crc_data[2]\, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[10]\);
    
    \lfsr_c_0_a2_1_0_x2_0_x2_0_x2[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => N_706, B => \tx_crc_data[15]\, Y => N_567_i);
    
    \lfsr_q[2]\ : SLE
      port map(D => N_617_i, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[2]\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \lfsr_q[1]\ : SLE
      port map(D => \lfsr_c[1]\, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[1]\);
    
    \lfsr_q[7]\ : SLE
      port map(D => N_622_i, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[7]\);
    
    \lfsr_c_0_a2_2_x2_1_x2_2_x2[4]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \tx_crc_data[10]\, B => \tx_crc_data[11]\, C
         => N_710, D => N_709, Y => N_619_i);
    
    \lfsr_q[4]\ : SLE
      port map(D => N_619_i, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[4]\);
    
    \lfsr_q[11]\ : SLE
      port map(D => \tx_crc_data[3]\, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[11]\);
    
    \lfsr_c_0_a2_0_x2_1_x2_1_x2[5]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \tx_crc_data[12]\, B => \tx_crc_data[11]\, C
         => N_709, D => N_704, Y => N_618_i);
    
    \lfsr_q[5]\ : SLE
      port map(D => N_618_i, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[5]\);
    
    \lfsr_c_0_a2[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => N_567_i, B => \tx_crc_data[1]\, Y => 
        \lfsr_c[9]\);
    
    \lfsr_c_0_a2[1]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => N_618_i, B => N_620_i, C => N_567_i, D => 
        N_622_i, Y => \lfsr_c[1]\);
    
    \lfsr_q[0]\ : SLE
      port map(D => \lfsr_c[0]\, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[0]\);
    
    \lfsr_c_0_a2[15]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => N_705, B => \lfsr_c[1]\, C => 
        \tx_crc_data[7]\, D => \tx_crc_data[8]\, Y => 
        \lfsr_c[15]\);
    
    \lfsr_q[12]\ : SLE
      port map(D => \tx_crc_data[4]\, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[12]\);
    
    lfsr_q_0_sqmuxa : CFG2
      generic map(INIT => x"8")

      port map(A => byte_clk_en, B => tx_crc_gen, Y => 
        \lfsr_q_0_sqmuxa\);
    
    \lfsr_c_0_a2_2_x2_1_x2_1_x2[2]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \tx_crc_data[9]\, B => \tx_crc_data[8]\, C
         => N_711, D => N_705, Y => N_617_i);
    
    \lfsr_q[14]\ : SLE
      port map(D => \tx_crc_data[6]\, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[14]\);
    
    \lfsr_c_0_a2_i_x2[8]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \tx_crc_data[14]\, B => \tx_crc_data[0]\, C
         => N_567_i, D => N_707, Y => N_107_i_i);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \lfsr_c_0_a2_2_x2_1_x2_1_x2[6]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \tx_crc_data[13]\, B => \tx_crc_data[12]\, C
         => N_708, D => N_704, Y => N_621_i);
    
    \lfsr_q[8]\ : SLE
      port map(D => N_107_i_i, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[8]\);
    
    \lfsr_q[13]\ : SLE
      port map(D => \tx_crc_data[5]\, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[13]\);
    
    \lfsr_c_0_a2[0]\ : CFG3
      generic map(INIT => x"96")

      port map(A => N_705, B => \lfsr_c[1]\, C => 
        \tx_crc_data[8]\, Y => \lfsr_c[0]\);
    
    \lfsr_q[15]\ : SLE
      port map(D => \lfsr_c[15]\, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[15]\);
    
    \lfsr_c_0_a2_0_x2_2_x2_0_x2[7]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \tx_crc_data[14]\, B => \tx_crc_data[13]\, C
         => N_708, D => N_707, Y => N_622_i);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity TX_Collision_Detector is

    port( un2_apb3_reset      : in    std_logic;
          external_loopback   : in    std_logic;
          internal_loopback   : in    std_logic;
          DRVR_EN_c           : in    std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          tx_col_detect_en    : out   std_logic
        );

end TX_Collision_Detector;

architecture DEF_ARCH of TX_Collision_Detector is 

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \tx_col_detect_en_0\, GND_net_1, 
        un10_reset : std_logic;

begin 


    tx_col_detect_en_0 : CFG2
      generic map(INIT => x"4")

      port map(A => un10_reset, B => DRVR_EN_c, Y => 
        \tx_col_detect_en_0\);
    
    \tx_col_detect_en\ : SLE
      port map(D => \tx_col_detect_en_0\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => tx_col_detect_en);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \SYNCH_PROC.un10_reset\ : CFG3
      generic map(INIT => x"FE")

      port map(A => internal_loopback, B => external_loopback, C
         => un2_apb3_reset, Y => un10_reset);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity IdleLineDetector_0 is

    port( manches_in_dly      : in    std_logic_vector(1 downto 0);
          idle_line5          : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          un2_apb3_reset_i    : in    std_logic;
          tx_idle_line        : out   std_logic
        );

end IdleLineDetector_0;

architecture DEF_ARCH of IdleLineDetector_0 is 

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal VCC_net_1, N_1351_i, GND_net_1, 
        \idle_line_cntr[0]_net_1\, \idle_line_cntr_s[0]\, 
        \idle_line_cntr[1]_net_1\, \idle_line_cntr_s[1]\, 
        \idle_line_cntr[2]_net_1\, \idle_line_cntr_s[2]\, 
        \idle_line_cntr[3]_net_1\, \idle_line_cntr_s[3]\, 
        \idle_line_cntr[4]_net_1\, \idle_line_cntr_s[4]\, 
        \idle_line_cntr[5]_net_1\, \idle_line_cntr_s[5]\, 
        \idle_line_cntr[6]_net_1\, \idle_line_cntr_s[6]\, 
        \idle_line_cntr[7]_net_1\, \idle_line_cntr_s[7]\, 
        \idle_line_cntr[8]_net_1\, \idle_line_cntr_s[8]\, 
        \idle_line_cntr[9]_net_1\, \idle_line_cntr_s[9]\, 
        \idle_line_cntr[10]_net_1\, \idle_line_cntr_s[10]\, 
        \idle_line_cntr[11]_net_1\, \idle_line_cntr_s[11]\, 
        \idle_line_cntr[12]_net_1\, \idle_line_cntr_s[12]\, 
        \idle_line_cntr[13]_net_1\, \idle_line_cntr_s[13]\, 
        \idle_line_cntr[14]_net_1\, \idle_line_cntr_s[14]\, 
        \idle_line_cntr[15]_net_1\, \idle_line_cntr_s[15]\, 
        idle_line_cntr_cry_cy, un5_manches_in_dly_9_RNIQSC51_Y, 
        \idle_line5\, un5_manches_in_dly_9, un5_manches_in_dly_10, 
        un5_manches_in_dly_11, \idle_line_cntr_cry[0]\, 
        \idle_line_cntr_cry[1]\, \idle_line_cntr_cry[2]\, 
        \idle_line_cntr_cry[3]\, \idle_line_cntr_cry[4]\, 
        \idle_line_cntr_cry[5]\, \idle_line_cntr_cry[6]\, 
        \idle_line_cntr_cry[7]\, \idle_line_cntr_cry[8]\, 
        \idle_line_cntr_cry[9]\, \idle_line_cntr_cry[10]\, 
        \idle_line_cntr_cry[11]\, \idle_line_cntr_cry[12]\, 
        \idle_line_cntr_cry[13]\, \idle_line_cntr_cry[14]\, 
        un5_manches_in_dly_8 : std_logic;

begin 

    idle_line5 <= \idle_line5\;

    \idle_line_cntr_RNICPKC7[3]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[3]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[2]\, S => \idle_line_cntr_s[3]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[3]\);
    
    idle_line : SLE
      port map(D => N_1351_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        tx_idle_line);
    
    \IDLE_LINE_DETECT_PROC.un5_manches_in_dly_11\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \idle_line_cntr[11]_net_1\, B => 
        \idle_line_cntr[8]_net_1\, C => \idle_line_cntr[7]_net_1\, 
        D => un5_manches_in_dly_8, Y => un5_manches_in_dly_11);
    
    \idle_line_cntr_RNIE6TJD[7]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[7]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[6]\, S => \idle_line_cntr_s[7]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[7]\);
    
    \idle_line_cntr[4]\ : SLE
      port map(D => \idle_line_cntr_s[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[4]_net_1\);
    
    \idle_line_cntr[14]\ : SLE
      port map(D => \idle_line_cntr_s[14]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[14]_net_1\);
    
    \idle_line_cntr_RNIDQ6N2[0]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[0]_net_1\, D => GND_net_1, FCI => 
        idle_line_cntr_cry_cy, S => \idle_line_cntr_s[0]\, Y => 
        OPEN, FCO => \idle_line_cntr_cry[0]\);
    
    \idle_line_cntr_RNI2800M[11]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[11]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[10]\, S => \idle_line_cntr_s[11]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[11]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \IDLE_LINE_DETECT_PROC.un5_manches_in_dly_9\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \idle_line_cntr[10]_net_1\, B => 
        \idle_line_cntr[9]_net_1\, C => \idle_line_cntr[2]_net_1\, 
        D => \idle_line_cntr[1]_net_1\, Y => un5_manches_in_dly_9);
    
    \IDLE_LINE_DETECT_PROC.un5_manches_in_dly_10\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \idle_line_cntr[6]_net_1\, B => 
        \idle_line_cntr[5]_net_1\, C => \idle_line_cntr[4]_net_1\, 
        D => \idle_line_cntr[3]_net_1\, Y => 
        un5_manches_in_dly_10);
    
    \idle_line_cntr_RNINOFCQ[14]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[14]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[13]\, S => \idle_line_cntr_s[14]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[14]\);
    
    \idle_line_cntr[9]\ : SLE
      port map(D => \idle_line_cntr_s[9]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[9]_net_1\);
    
    \idle_line_cntr[8]\ : SLE
      port map(D => \idle_line_cntr_s[8]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[8]_net_1\);
    
    \idle_line_cntr[7]\ : SLE
      port map(D => \idle_line_cntr_s[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[7]_net_1\);
    
    \idle_line_cntr[15]\ : SLE
      port map(D => \idle_line_cntr_s[15]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[15]_net_1\);
    
    \idle_line_cntr[11]\ : SLE
      port map(D => \idle_line_cntr_s[11]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[11]_net_1\);
    
    \idle_line_cntr[10]\ : SLE
      port map(D => \idle_line_cntr_s[10]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[10]_net_1\);
    
    \idle_line_cntr[1]\ : SLE
      port map(D => \idle_line_cntr_s[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[1]_net_1\);
    
    \idle_line_cntr_RNIK132C[6]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[6]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[5]\, S => \idle_line_cntr_s[6]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[6]\);
    
    \IDLE_LINE_DETECT_PROC.un5_manches_in_dly_8\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \idle_line_cntr[15]_net_1\, B => 
        \idle_line_cntr[14]_net_1\, C => 
        \idle_line_cntr[13]_net_1\, D => 
        \idle_line_cntr[12]_net_1\, Y => un5_manches_in_dly_8);
    
    \idle_line_cntr_RNIF7LTO[13]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[13]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[12]\, S => \idle_line_cntr_s[13]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[13]\);
    
    \idle_line_cntr_RNI9CN5F[8]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[8]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[7]\, S => \idle_line_cntr_s[8]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[8]\);
    
    \idle_line_cntr_RNO[15]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[15]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[14]\, S => \idle_line_cntr_s[15]\, Y
         => OPEN, FCO => OPEN);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \idle_line_cntr_RNITP5HK[10]\ : ARI1
      generic map(INIT => x"4D800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[10]_net_1\, D => N_1351_i, FCI => 
        \idle_line_cntr_cry[9]\, S => \idle_line_cntr_s[10]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[10]\);
    
    \idle_line_cntr_RNIVFUSH[9]\ : ARI1
      generic map(INIT => x"4D800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[9]_net_1\, D => N_1351_i, FCI => 
        \idle_line_cntr_cry[8]\, S => \idle_line_cntr_s[9]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[9]\);
    
    \idle_line_cntr_RNI1P094[1]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[1]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[0]\, S => \idle_line_cntr_s[1]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[1]\);
    
    \idle_line_cntr[6]\ : SLE
      port map(D => \idle_line_cntr_s[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[6]_net_1\);
    
    \idle_line_cntr_RNIMOQQ5[2]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[2]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[1]\, S => \idle_line_cntr_s[2]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[2]\);
    
    \idle_line_cntr_RNI3REU8[4]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[4]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[3]\, S => \idle_line_cntr_s[4]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[4]\);
    
    \idle_line_cntr_RNIRT8GA[5]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[5]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[4]\, S => \idle_line_cntr_s[5]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[5]\);
    
    \idle_line_cntr[13]\ : SLE
      port map(D => \idle_line_cntr_s[13]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[13]_net_1\);
    
    \idle_line_cntr[0]\ : SLE
      port map(D => \idle_line_cntr_s[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[0]_net_1\);
    
    \IDLE_LINE_DETECT_PROC.un5_manches_in_dly_9_RNIQSC51\ : ARI1
      generic map(INIT => x"41555")

      port map(A => un5_manches_in_dly_11, B => \idle_line5\, C
         => un5_manches_in_dly_9, D => un5_manches_in_dly_10, FCI
         => VCC_net_1, S => OPEN, Y => 
        un5_manches_in_dly_9_RNIQSC51_Y, FCO => 
        idle_line_cntr_cry_cy);
    
    \idle_line_cntr_RNI8NQEN[12]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[12]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[11]\, S => \idle_line_cntr_s[12]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[12]\);
    
    \idle_line_cntr[12]\ : SLE
      port map(D => \idle_line_cntr_s[12]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[12]_net_1\);
    
    \idle_line_cntr[3]\ : SLE
      port map(D => \idle_line_cntr_s[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[3]_net_1\);
    
    un4_manches_in_dly : CFG2
      generic map(INIT => x"6")

      port map(A => manches_in_dly(1), B => manches_in_dly(0), Y
         => \idle_line5\);
    
    \IDLE_LINE_DETECT_PROC.un5_manches_in_dly_9_RNIQSC51_0\ : 
        CFG4
      generic map(INIT => x"4000")

      port map(A => \idle_line5\, B => un5_manches_in_dly_11, C
         => un5_manches_in_dly_10, D => un5_manches_in_dly_9, Y
         => N_1351_i);
    
    \idle_line_cntr[5]\ : SLE
      port map(D => \idle_line_cntr_s[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[5]_net_1\);
    
    \idle_line_cntr[2]\ : SLE
      port map(D => \idle_line_cntr_s[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[2]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity TX_SM is

    port( manches_in_dly                  : in    std_logic_vector(1 downto 0);
          CommsFPGA_CCC_0_GL0             : in    std_logic;
          idle_line5                      : out   std_logic;
          TX_FIFO_Empty                   : in    std_logic;
          N_705                           : in    std_logic;
          N_706                           : in    std_logic;
          N_707                           : in    std_logic;
          N_708                           : in    std_logic;
          N_704                           : in    std_logic;
          N_709                           : in    std_logic;
          N_710                           : in    std_logic;
          N_711                           : in    std_logic;
          TX_DataEn                       : out   std_logic;
          TX_PreAmble                     : out   std_logic;
          tx_crc_byte1_en                 : out   std_logic;
          tx_crc_byte2_en                 : out   std_logic;
          tx_packet_complt                : out   std_logic;
          tx_crc_gen                      : out   std_logic;
          TX_DataEn_1_o                   : out   std_logic;
          un1_tx_packet_length_0_sqmuxa_o : out   std_logic;
          start_tx_FIFO                   : in    std_logic;
          DRVR_EN_c                       : out   std_logic;
          byte_clk_en                     : in    std_logic;
          tx_preamble_pat_en              : out   std_logic;
          BIT_CLK                         : in    std_logic;
          un2_apb3_reset_i                : in    std_logic
        );

end TX_SM;

architecture DEF_ARCH of TX_SM is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component IdleLineDetector_0
    port( manches_in_dly      : in    std_logic_vector(1 downto 0) := (others => 'U');
          idle_line5          : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          un2_apb3_reset_i    : in    std_logic := 'U';
          tx_idle_line        : out   std_logic
        );
  end component;

    signal un25_tx_byte_cntr_a_4_cry_9, 
        \un25_tx_byte_cntr_a_4_i[11]\, \TX_STATE[8]_net_1\, 
        \TX_STATE_i_0[8]\, \un25_tx_byte_cntr_a_4[6]\, GND_net_1, 
        \un25_tx_byte_cntr_a_4_i[6]\, un1_byte_clk_en_inv_2_i, 
        VCC_net_1, \un25_tx_byte_cntr_a_4[7]\, 
        \un25_tx_byte_cntr_a_4_i[7]\, \un25_tx_byte_cntr_a_4[8]\, 
        \un25_tx_byte_cntr_a_4_i[8]\, \un25_tx_byte_cntr_a_4[9]\, 
        \un25_tx_byte_cntr_a_4_i[9]\, \un25_tx_byte_cntr_a_4[10]\, 
        \un25_tx_byte_cntr_a_4_i[10]\, 
        \un25_tx_byte_cntr_a_4[11]\, \tx_packet_length[1]_net_1\, 
        \un25_tx_byte_cntr_a_4_i_i[1]\, 
        \tx_packet_length[2]_net_1\, 
        un25_tx_byte_cntr_a_4_axb_1_i, 
        \tx_packet_length[3]_net_1\, 
        un25_tx_byte_cntr_a_4_axb_2_i, 
        \tx_packet_length[4]_net_1\, 
        un25_tx_byte_cntr_a_4_axb_3_i, 
        \tx_packet_length[5]_net_1\, 
        un25_tx_byte_cntr_a_4_axb_4_i, 
        \tx_packet_length[6]_net_1\, 
        un25_tx_byte_cntr_a_4_axb_5_i, 
        \tx_packet_length[7]_net_1\, 
        un25_tx_byte_cntr_a_4_axb_6_i, 
        \tx_packet_length[8]_net_1\, N_15_i, 
        \tx_packet_length[9]_net_1\, N_13_i, 
        \tx_packet_length[10]_net_1\, 
        un25_tx_byte_cntr_a_4_axb_9_i, \un25_tx_byte_cntr_a_4[1]\, 
        un25_tx_byte_cntr_a_4_cry_0_Y, \un25_tx_byte_cntr_a_4[2]\, 
        \un25_tx_byte_cntr_a_4_i[2]\, \un25_tx_byte_cntr_a_4[3]\, 
        \un25_tx_byte_cntr_a_4_i[3]\, \un25_tx_byte_cntr_a_4[4]\, 
        \un25_tx_byte_cntr_a_4_i[4]\, \un25_tx_byte_cntr_a_4[5]\, 
        \un25_tx_byte_cntr_a_4_i[5]\, \tx_packet_length[0]_net_1\, 
        N_19_i, TX_DataEn_1_m, \tx_idle_line_s\, tx_idle_line, 
        \start_tx_FIFO_s\, \TX_STATE[3]_net_1\, \TX_STATE_69\, 
        \TX_STATE[4]_net_1\, \TX_STATE_68\, \TX_STATE[5]_net_1\, 
        \TX_STATE_67\, \TX_STATE[6]_net_1\, \TX_STATE_66\, 
        \TX_STATE[7]_net_1\, \TX_STATE_65\, \TX_STATE_64\, 
        \un1_tx_packet_length_0_sqmuxa_o\, 
        \iTX_FIFO_rd_en_ret_1_RNO\, N_589, 
        \tx_byte_cntr_cry_cy_Y[0]\, \TX_STATE[0]_net_1\, 
        \TX_STATE[2]_net_1\, TX_PreAmble_net_1, \TX_PreAmble_34\, 
        TX_DataEn_7, \TX_STATE_72\, \TX_STATE[1]_net_1\, 
        \TX_STATE_71\, \TX_STATE_70\, \PostAmble_cntr[0]_net_1\, 
        \PostAmble_cntr_s[0]\, \PostAmble_cntr[1]_net_1\, 
        \PostAmble_cntr_s[1]\, \PostAmble_cntr[2]_net_1\, 
        \PostAmble_cntr_s[2]\, \PostAmble_cntr[3]_net_1\, 
        \PostAmble_cntr_s[3]\, \PostAmble_cntr[4]_net_1\, 
        \PostAmble_cntr_s[4]\, \PostAmble_cntr[5]_net_1\, 
        \PostAmble_cntr_s[5]\, \PostAmble_cntr[6]_net_1\, 
        \PostAmble_cntr_s[6]\, \PostAmble_cntr[7]_net_1\, 
        \PostAmble_cntr_s[7]\, \PostAmble_cntr[8]_net_1\, 
        \PostAmble_cntr_s[8]\, \PostAmble_cntr[9]_net_1\, 
        \PostAmble_cntr_s[9]\, \PostAmble_cntr[10]_net_1\, 
        \PostAmble_cntr_s[10]\, \PostAmble_cntr[11]_net_1\, 
        \PostAmble_cntr_s[11]\, \txen_early_cntr[0]_net_1\, 
        \txen_early_cntr_s[0]\, \txen_early_cntr[1]_net_1\, 
        \txen_early_cntr_s[1]\, \txen_early_cntr[2]_net_1\, 
        \txen_early_cntr_s[2]\, \txen_early_cntr[3]_net_1\, 
        \txen_early_cntr_s[3]\, \txen_early_cntr[4]_net_1\, 
        \txen_early_cntr_s[4]\, \txen_early_cntr[5]_net_1\, 
        \txen_early_cntr_s[5]\, \txen_early_cntr[6]_net_1\, 
        \txen_early_cntr_s[6]\, \txen_early_cntr[7]_net_1\, 
        \txen_early_cntr_s[7]\, \txen_early_cntr[8]_net_1\, 
        \txen_early_cntr_s[8]\, \txen_early_cntr[9]_net_1\, 
        \txen_early_cntr_s[9]\, \txen_early_cntr[10]_net_1\, 
        \txen_early_cntr_s[10]\, \txen_early_cntr[11]_net_1\, 
        \txen_early_cntr_s[11]\, \tx_byte_cntr[0]_net_1\, 
        \tx_byte_cntr_s[0]\, \tx_byte_cntr[1]_net_1\, 
        \tx_byte_cntr_s[1]\, \tx_byte_cntr[2]_net_1\, 
        \tx_byte_cntr_s[2]\, \tx_byte_cntr[3]_net_1\, 
        \tx_byte_cntr_s[3]\, \tx_byte_cntr[4]_net_1\, 
        \tx_byte_cntr_s[4]\, \tx_byte_cntr[5]_net_1\, 
        \tx_byte_cntr_s[5]\, \tx_byte_cntr[6]_net_1\, 
        \tx_byte_cntr_s[6]\, \tx_byte_cntr[7]_net_1\, 
        \tx_byte_cntr_s[7]\, \tx_byte_cntr[8]_net_1\, 
        \tx_byte_cntr_s[8]\, \tx_byte_cntr[9]_net_1\, 
        \tx_byte_cntr_s[9]\, \tx_byte_cntr[10]_net_1\, 
        \tx_byte_cntr_s[10]\, \tx_byte_cntr[11]_net_1\, 
        \tx_byte_cntr_s[11]_net_1\, \PreAmble_cntr[0]_net_1\, 
        \PreAmble_cntr_s[0]\, N_329_i, \PreAmble_cntr[1]_net_1\, 
        \PreAmble_cntr_s[1]\, \PreAmble_cntr[2]_net_1\, 
        \PreAmble_cntr_s[2]\, \PreAmble_cntr[3]_net_1\, 
        \PreAmble_cntr_s[3]\, \PreAmble_cntr[4]_net_1\, 
        \PreAmble_cntr_s[4]\, \PreAmble_cntr[5]_net_1\, 
        \PreAmble_cntr_s[5]\, \PreAmble_cntr[6]_net_1\, 
        \PreAmble_cntr_s[6]\, PostAmble_cntr_cry_cy, 
        tx_state29_6_RNI9SJ61_Y, tx_state29_6, tx_state29_7, 
        tx_state29_8, \PostAmble_cntr_cry[0]\, 
        \PostAmble_cntr_cry[1]\, \PostAmble_cntr_cry[2]\, 
        \PostAmble_cntr_cry[3]\, \PostAmble_cntr_cry[4]\, 
        \PostAmble_cntr_cry[5]\, \PostAmble_cntr_cry[6]\, 
        \PostAmble_cntr_cry[7]\, \PostAmble_cntr_cry[8]\, 
        \PostAmble_cntr_cry[9]\, \PostAmble_cntr_cry[10]\, 
        txen_early_cntr_cry_cy, \TX_STATE_RNIAIGV2_Y[7]\, m15_e_6, 
        m15_e_7, m15_e_8, \txen_early_cntr_cry[0]\, 
        \txen_early_cntr_cry[1]\, \txen_early_cntr_cry[2]\, 
        \txen_early_cntr_cry[3]\, \txen_early_cntr_cry[4]\, 
        \txen_early_cntr_cry[5]\, \txen_early_cntr_cry[6]\, 
        \txen_early_cntr_cry[7]\, \txen_early_cntr_cry[8]\, 
        \txen_early_cntr_cry[9]\, \txen_early_cntr_cry[10]\, 
        tx_byte_cntr_cry_cy, \tx_byte_cntr_cry[0]_net_1\, 
        \tx_byte_cntr_cry[1]_net_1\, \tx_byte_cntr_cry[2]_net_1\, 
        \tx_byte_cntr_cry[3]_net_1\, \tx_byte_cntr_cry[4]_net_1\, 
        \tx_byte_cntr_cry[5]_net_1\, \tx_byte_cntr_cry[6]_net_1\, 
        \tx_byte_cntr_cry[7]_net_1\, \tx_byte_cntr_cry[8]_net_1\, 
        \tx_byte_cntr_cry[9]_net_1\, \tx_byte_cntr_cry[10]_net_1\, 
        PreAmble_cntr_cry_cy, \PreAmble_cntr_RNIHNV31_Y[6]\, 
        PreAmble_cntr_0_sqmuxa_0_83_i_o3_0, 
        PreAmble_cntr_0_sqmuxa_0_83_i_o3_4, 
        \PreAmble_cntr_cry[0]\, \PreAmble_cntr_cry[1]\, 
        \PreAmble_cntr_cry[2]\, \PreAmble_cntr_cry[3]\, 
        \PreAmble_cntr_cry[4]\, \PreAmble_cntr_cry[5]\, 
        un25_tx_byte_cntr_a_4_cry_0, N_81, 
        un25_tx_byte_cntr_a_4_cry_1, un25_tx_byte_cntr_a_4_cry_2, 
        un25_tx_byte_cntr_a_4_cry_3, un25_tx_byte_cntr_a_4_cry_4, 
        un25_tx_byte_cntr_a_4_cry_5, un25_tx_byte_cntr_a_4_cry_6, 
        un25_tx_byte_cntr_a_4_cry_7, un25_tx_byte_cntr_a_4_cry_8, 
        \un25_tx_byte_cntr_1_data_tmp[0]\, 
        \un25_tx_byte_cntr_1_data_tmp[1]\, 
        \un25_tx_byte_cntr_1_data_tmp[2]\, 
        \un25_tx_byte_cntr_1_data_tmp[3]\, 
        \un25_tx_byte_cntr_1_data_tmp[4]\, un25_tx_byte_cntr, 
        N_213_i, m56_i_0_0_0, un14_tx_byte_cntr_0_a2_8_a2_0_6_1, 
        un9_start_tx_fifo_s, N_1390, 
        \un1_byte_clk_en_inv_2_0_0_0_2\, 
        un14_tx_byte_cntr_0_a2_8_a2_0_5, N_957, N_1447, N_719, 
        N_80, N_1383, un14_tx_byte_cntr_0_a2_8_a2_0_6, N_1336, 
        N_1388, N_1355 : std_logic;

    for all : IdleLineDetector_0
	Use entity work.IdleLineDetector_0(DEF_ARCH);
begin 

    TX_PreAmble <= TX_PreAmble_net_1;
    un1_tx_packet_length_0_sqmuxa_o <= 
        \un1_tx_packet_length_0_sqmuxa_o\;

    iTX_FIFO_rd_en_ret_1 : SLE
      port map(D => \iTX_FIFO_rd_en_ret_1_RNO\, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \un1_tx_packet_length_0_sqmuxa_o\);
    
    \tx_packet_length_RNO[2]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => N_81, B => N_710, C => 
        \tx_packet_length[2]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => un25_tx_byte_cntr_a_4_axb_1_i);
    
    \txen_early_cntr_RNIJFKLC[2]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \txen_early_cntr[2]_net_1\, C
         => \TX_STATE_RNIAIGV2_Y[7]\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[1]\, S => \txen_early_cntr_s[2]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[2]\);
    
    \tx_byte_cntr[8]\ : SLE
      port map(D => \tx_byte_cntr_s[8]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_byte_cntr[8]_net_1\);
    
    \tx_byte_cntr[2]\ : SLE
      port map(D => \tx_byte_cntr_s[2]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_byte_cntr[2]_net_1\);
    
    \PreAmble_cntr[6]\ : SLE
      port map(D => \PreAmble_cntr_s[6]\, CLK => BIT_CLK, EN => 
        N_329_i, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PreAmble_cntr[6]_net_1\);
    
    \PreAmble_cntr_RNI4FPH8[5]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \PreAmble_cntr_RNIHNV31_Y[6]\, 
        C => \PreAmble_cntr[5]_net_1\, D => GND_net_1, FCI => 
        \PreAmble_cntr_cry[4]\, S => \PreAmble_cntr_s[5]\, Y => 
        OPEN, FCO => \PreAmble_cntr_cry[5]\);
    
    \TX_SM.un14_tx_byte_cntr_0_a2_8_a2_0_5\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \tx_byte_cntr[9]_net_1\, B => 
        \tx_byte_cntr[8]_net_1\, C => \tx_byte_cntr[7]_net_1\, D
         => \tx_byte_cntr[4]_net_1\, Y => 
        un14_tx_byte_cntr_0_a2_8_a2_0_5);
    
    \PreAmble_cntr_RNI7UJB2[0]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \PreAmble_cntr_RNIHNV31_Y[6]\, 
        C => \PreAmble_cntr[0]_net_1\, D => GND_net_1, FCI => 
        PreAmble_cntr_cry_cy, S => \PreAmble_cntr_s[0]\, Y => 
        OPEN, FCO => \PreAmble_cntr_cry[0]\);
    
    \TX_STATE[7]\ : SLE
      port map(D => \TX_STATE_65\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_STATE[7]_net_1\);
    
    \tx_packet_length_ret_0[10]\ : SLE
      port map(D => \un25_tx_byte_cntr_a_4_i[11]\, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => un2_apb3_reset_i, 
        ADn => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \un25_tx_byte_cntr_a_4[11]\);
    
    \TX_STATE_ns_8_0_.m56_i_0_0_a2\ : CFG4
      generic map(INIT => x"E000")

      port map(A => N_957, B => N_1447, C => 
        un14_tx_byte_cntr_0_a2_8_a2_0_5, D => 
        un14_tx_byte_cntr_0_a2_8_a2_0_6, Y => N_1336);
    
    \tx_byte_cntr_cry[7]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[7]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[6]_net_1\, S => \tx_byte_cntr_s[7]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[7]_net_1\);
    
    start_tx_FIFO_s : SLE
      port map(D => start_tx_FIFO, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \start_tx_FIFO_s\);
    
    \tx_packet_length[4]\ : SLE
      port map(D => un25_tx_byte_cntr_a_4_axb_3_i, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => un2_apb3_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \tx_packet_length[4]_net_1\);
    
    \tx_byte_cntr[0]\ : SLE
      port map(D => \tx_byte_cntr_s[0]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_byte_cntr[0]_net_1\);
    
    \tx_packet_length[1]\ : SLE
      port map(D => \un25_tx_byte_cntr_a_4_i_i[1]\, CLK => 
        BIT_CLK, EN => un1_byte_clk_en_inv_2_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \tx_packet_length[1]_net_1\);
    
    \txen_early_cntr_RNI5MOBM[5]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \txen_early_cntr[5]_net_1\, C
         => \TX_STATE_RNIAIGV2_Y[7]\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[4]\, S => \txen_early_cntr_s[5]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[5]\);
    
    \TX_SM.un25_tx_byte_cntr_a_4_cry_7\ : ARI1
      generic map(INIT => x"63B7F")

      port map(A => N_705, B => N_81, C => \TX_STATE[5]_net_1\, D
         => \tx_packet_length[8]_net_1\, FCI => 
        un25_tx_byte_cntr_a_4_cry_6, S => 
        \un25_tx_byte_cntr_a_4_i[8]\, Y => OPEN, FCO => 
        un25_tx_byte_cntr_a_4_cry_7);
    
    \tx_packet_length_ret_0[1]\ : SLE
      port map(D => \un25_tx_byte_cntr_a_4_i[2]\, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => un2_apb3_reset_i, 
        ADn => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \un25_tx_byte_cntr_a_4[2]\);
    
    \tx_byte_cntr_cry[4]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[4]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[3]_net_1\, S => \tx_byte_cntr_s[4]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[4]_net_1\);
    
    \PostAmble_cntr_RNIMPNEJ[10]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => tx_state29_6_RNI9SJ61_Y, C
         => \PostAmble_cntr[10]_net_1\, D => GND_net_1, FCI => 
        \PostAmble_cntr_cry[9]\, S => \PostAmble_cntr_s[10]\, Y
         => OPEN, FCO => \PostAmble_cntr_cry[10]\);
    
    TX_STATE_69 : CFG4
      generic map(INIT => x"11F0")

      port map(A => m56_i_0_0_0, B => N_1336, C => 
        \TX_STATE[3]_net_1\, D => byte_clk_en, Y => \TX_STATE_69\);
    
    \tx_packet_length_RNO[6]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => N_81, B => N_707, C => 
        \tx_packet_length[6]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => un25_tx_byte_cntr_a_4_axb_5_i);
    
    \tx_packet_length_RNO[3]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => N_81, B => N_709, C => 
        \tx_packet_length[3]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => un25_tx_byte_cntr_a_4_axb_2_i);
    
    \TX_STATE[2]\ : SLE
      port map(D => \TX_STATE_70\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_STATE[2]_net_1\);
    
    \TX_PreAmble\ : SLE
      port map(D => \TX_PreAmble_34\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        TX_PreAmble_net_1);
    
    \tx_packet_length_ret_0_RNO[10]\ : CFG1
      generic map(INIT => "01")

      port map(A => un25_tx_byte_cntr_a_4_cry_9, Y => 
        \un25_tx_byte_cntr_a_4_i[11]\);
    
    \tx_packet_length[9]\ : SLE
      port map(D => N_13_i, CLK => BIT_CLK, EN => 
        un1_byte_clk_en_inv_2_i, ALn => un2_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_packet_length[9]_net_1\);
    
    \tx_packet_length_ret_0[6]\ : SLE
      port map(D => \un25_tx_byte_cntr_a_4_i[7]\, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => un2_apb3_reset_i, 
        ADn => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \un25_tx_byte_cntr_a_4[7]\);
    
    \PreAmble_cntr_RNIH597[3]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \PreAmble_cntr[3]_net_1\, B => 
        \PreAmble_cntr[4]_net_1\, Y => 
        PreAmble_cntr_0_sqmuxa_0_83_i_o3_0);
    
    \txen_early_cntr_RNIFF8E9[1]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \txen_early_cntr[1]_net_1\, C
         => \TX_STATE_RNIAIGV2_Y[7]\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[0]\, S => \txen_early_cntr_s[1]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[1]\);
    
    \TX_STATE_ns_8_0_.m55_0_a3_0_a2_0_a2\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_589, B => \TX_STATE[6]_net_1\, Y => 
        TX_DataEn_1_m);
    
    \txen_early_cntr[5]\ : SLE
      port map(D => \txen_early_cntr_s[5]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => un2_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \txen_early_cntr[5]_net_1\);
    
    \PreAmble_cntr_RNI935A7[4]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \PreAmble_cntr_RNIHNV31_Y[6]\, 
        C => \PreAmble_cntr[4]_net_1\, D => GND_net_1, FCI => 
        \PreAmble_cntr_cry[3]\, S => \PreAmble_cntr_s[4]\, Y => 
        OPEN, FCO => \PreAmble_cntr_cry[4]\);
    
    TX_PreAmble_34 : CFG3
      generic map(INIT => x"AC")

      port map(A => \TX_STATE[6]_net_1\, B => TX_PreAmble_net_1, 
        C => byte_clk_en, Y => \TX_PreAmble_34\);
    
    \tx_packet_length_ret_0[7]\ : SLE
      port map(D => \un25_tx_byte_cntr_a_4_i[8]\, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => un2_apb3_reset_i, 
        ADn => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \un25_tx_byte_cntr_a_4[8]\);
    
    \tx_byte_cntr[6]\ : SLE
      port map(D => \tx_byte_cntr_s[6]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_byte_cntr[6]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \tx_crc_byte2_en\ : SLE
      port map(D => \TX_STATE[2]_net_1\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => tx_crc_byte2_en);
    
    \tx_packet_length_RNO[0]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => N_81, B => N_705, C => 
        \tx_packet_length[0]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => N_19_i);
    
    \tx_byte_cntr_cry[10]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[10]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[9]_net_1\, S => \tx_byte_cntr_s[10]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[10]_net_1\);
    
    \PreAmble_cntr_RNO[6]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \PreAmble_cntr_RNIHNV31_Y[6]\, 
        C => \PreAmble_cntr[6]_net_1\, D => GND_net_1, FCI => 
        \PreAmble_cntr_cry[5]\, S => \PreAmble_cntr_s[6]\, Y => 
        OPEN, FCO => OPEN);
    
    \tx_packet_length[3]\ : SLE
      port map(D => un25_tx_byte_cntr_a_4_axb_2_i, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => un2_apb3_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \tx_packet_length[3]_net_1\);
    
    \PreAmble_cntr[1]\ : SLE
      port map(D => \PreAmble_cntr_s[1]\, CLK => BIT_CLK, EN => 
        N_329_i, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PreAmble_cntr[1]_net_1\);
    
    un1_byte_clk_en_inv_2_0_0_0_2 : CFG4
      generic map(INIT => x"FFFB")

      port map(A => \TX_STATE[2]_net_1\, B => byte_clk_en, C => 
        \TX_STATE[4]_net_1\, D => \TX_STATE[3]_net_1\, Y => 
        \un1_byte_clk_en_inv_2_0_0_0_2\);
    
    \PostAmble_cntr[6]\ : SLE
      port map(D => \PostAmble_cntr_s[6]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \PostAmble_cntr[6]_net_1\);
    
    \tx_byte_cntr_s[11]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[11]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[10]_net_1\, S => 
        \tx_byte_cntr_s[11]_net_1\, Y => OPEN, FCO => OPEN);
    
    \txen_early_cntr[8]\ : SLE
      port map(D => \txen_early_cntr_s[8]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => un2_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \txen_early_cntr[8]_net_1\);
    
    \tx_byte_cntr[5]\ : SLE
      port map(D => \tx_byte_cntr_s[5]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_byte_cntr[5]_net_1\);
    
    \TX_STATE[0]\ : SLE
      port map(D => \TX_STATE_72\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_STATE[0]_net_1\);
    
    \TX_SM.TX_DataEn_7_iv\ : CFG3
      generic map(INIT => x"8F")

      port map(A => N_589, B => \TX_STATE[6]_net_1\, C => N_213_i, 
        Y => TX_DataEn_7);
    
    \PostAmble_cntr_RNI342U7[3]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => tx_state29_6_RNI9SJ61_Y, C
         => \PostAmble_cntr[3]_net_1\, D => GND_net_1, FCI => 
        \PostAmble_cntr_cry[2]\, S => \PostAmble_cntr_s[3]\, Y
         => OPEN, FCO => \PostAmble_cntr_cry[3]\);
    
    \TX_STATE_ns_8_0_.m38_i_0_0_a2_0\ : CFG4
      generic map(INIT => x"8000")

      port map(A => m15_e_7, B => m15_e_6, C => 
        \TX_STATE[7]_net_1\, D => m15_e_8, Y => N_1388);
    
    iTX_Enable : SLE
      port map(D => \TX_STATE_i_0[8]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => DRVR_EN_c);
    
    \tx_byte_cntr_cry[2]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[2]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[1]_net_1\, S => \tx_byte_cntr_s[2]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[2]_net_1\);
    
    \PreAmble_cntr[3]\ : SLE
      port map(D => \PreAmble_cntr_s[3]\, CLK => BIT_CLK, EN => 
        N_329_i, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PreAmble_cntr[3]_net_1\);
    
    \tx_packet_length_ret_0[4]\ : SLE
      port map(D => \un25_tx_byte_cntr_a_4_i[5]\, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => un2_apb3_reset_i, 
        ADn => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \un25_tx_byte_cntr_a_4[5]\);
    
    \tx_packet_length[10]\ : SLE
      port map(D => un25_tx_byte_cntr_a_4_axb_9_i, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => un2_apb3_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \tx_packet_length[10]_net_1\);
    
    \txen_early_cntr_RNIUP0C61[10]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \txen_early_cntr[10]_net_1\, 
        C => \TX_STATE_RNIAIGV2_Y[7]\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[9]\, S => \txen_early_cntr_s[10]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[10]\);
    
    \tx_byte_cntr[11]\ : SLE
      port map(D => \tx_byte_cntr_s[11]_net_1\, CLK => BIT_CLK, 
        EN => byte_clk_en, ALn => un2_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_byte_cntr[11]_net_1\);
    
    \TX_SM.un25_tx_byte_cntr_a_4_cry_4\ : ARI1
      generic map(INIT => x"637BF")

      port map(A => N_708, B => N_81, C => \TX_STATE[5]_net_1\, D
         => \tx_packet_length[5]_net_1\, FCI => 
        un25_tx_byte_cntr_a_4_cry_3, S => 
        \un25_tx_byte_cntr_a_4_i[5]\, Y => OPEN, FCO => 
        un25_tx_byte_cntr_a_4_cry_4);
    
    \tx_byte_cntr_cry_cy[0]\ : ARI1
      generic map(INIT => x"4EE00")

      port map(A => VCC_net_1, B => \TX_STATE[4]_net_1\, C => 
        \TX_STATE[5]_net_1\, D => GND_net_1, FCI => VCC_net_1, S
         => OPEN, Y => \tx_byte_cntr_cry_cy_Y[0]\, FCO => 
        tx_byte_cntr_cry_cy);
    
    \tx_packet_length[5]\ : SLE
      port map(D => un25_tx_byte_cntr_a_4_axb_4_i, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => un2_apb3_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \tx_packet_length[5]_net_1\);
    
    \tx_packet_length_ret_0[0]\ : SLE
      port map(D => un25_tx_byte_cntr_a_4_cry_0_Y, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => un2_apb3_reset_i, 
        ADn => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \un25_tx_byte_cntr_a_4[1]\);
    
    \PreAmble_cntr_RNIFOG26[3]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \PreAmble_cntr_RNIHNV31_Y[6]\, 
        C => \PreAmble_cntr[3]_net_1\, D => GND_net_1, FCI => 
        \PreAmble_cntr_cry[2]\, S => \PreAmble_cntr_s[3]\, Y => 
        OPEN, FCO => \PreAmble_cntr_cry[3]\);
    
    \txen_early_cntr_RNIOG0TF[3]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \txen_early_cntr[3]_net_1\, C
         => \TX_STATE_RNIAIGV2_Y[7]\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[2]\, S => \txen_early_cntr_s[3]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[3]\);
    
    \PostAmble_cntr_RNI6EP9B[5]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => tx_state29_6_RNI9SJ61_Y, C
         => \PostAmble_cntr[5]_net_1\, D => GND_net_1, FCI => 
        \PostAmble_cntr_cry[4]\, S => \PostAmble_cntr_s[5]\, Y
         => OPEN, FCO => \PostAmble_cntr_cry[5]\);
    
    \txen_early_cntr[9]\ : SLE
      port map(D => \txen_early_cntr_s[9]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => un2_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \txen_early_cntr[9]_net_1\);
    
    \TX_STATE_RNIAIGV2[7]\ : ARI1
      generic map(INIT => x"42AAA")

      port map(A => m15_e_8, B => \TX_STATE[7]_net_1\, C => 
        m15_e_6, D => m15_e_7, FCI => VCC_net_1, S => OPEN, Y => 
        \TX_STATE_RNIAIGV2_Y[7]\, FCO => txen_early_cntr_cry_cy);
    
    \PostAmble_cntr[11]\ : SLE
      port map(D => \PostAmble_cntr_s[11]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => un2_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \PostAmble_cntr[11]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \tx_byte_cntr[4]\ : SLE
      port map(D => \tx_byte_cntr_s[4]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_byte_cntr[4]_net_1\);
    
    \txen_early_cntr[1]\ : SLE
      port map(D => \txen_early_cntr_s[1]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => un2_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \txen_early_cntr[1]_net_1\);
    
    \tx_byte_cntr_cry[0]\ : ARI1
      generic map(INIT => x"4A800")

      port map(A => VCC_net_1, B => \tx_byte_cntr[0]_net_1\, C
         => \TX_STATE[5]_net_1\, D => \TX_STATE[4]_net_1\, FCI
         => tx_byte_cntr_cry_cy, S => \tx_byte_cntr_s[0]\, Y => 
        OPEN, FCO => \tx_byte_cntr_cry[0]_net_1\);
    
    \TX_SM.un25_tx_byte_cntr_a_4_cry_6\ : ARI1
      generic map(INIT => x"637BF")

      port map(A => N_706, B => N_81, C => \TX_STATE[5]_net_1\, D
         => \tx_packet_length[7]_net_1\, FCI => 
        un25_tx_byte_cntr_a_4_cry_5, S => 
        \un25_tx_byte_cntr_a_4_i[7]\, Y => OPEN, FCO => 
        un25_tx_byte_cntr_a_4_cry_6);
    
    \TX_STATE_ns_8_0_.m56_i_0_0_0\ : CFG2
      generic map(INIT => x"B")

      port map(A => un25_tx_byte_cntr, B => \TX_STATE[5]_net_1\, 
        Y => m56_i_0_0_0);
    
    \TX_STATE_ns_8_0_.m15_e_6\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \txen_early_cntr[9]_net_1\, B => 
        \txen_early_cntr[8]_net_1\, C => 
        \txen_early_cntr[7]_net_1\, D => 
        \txen_early_cntr[6]_net_1\, Y => m15_e_6);
    
    \txen_early_cntr_RNIBD9931[9]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \txen_early_cntr[9]_net_1\, C
         => \TX_STATE_RNIAIGV2_Y[7]\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[8]\, S => \txen_early_cntr_s[9]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[9]\);
    
    \PostAmble_cntr_RNIDSGLE[7]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => tx_state29_6_RNI9SJ61_Y, C
         => \PostAmble_cntr[7]_net_1\, D => GND_net_1, FCI => 
        \PostAmble_cntr_cry[6]\, S => \PostAmble_cntr_s[7]\, Y
         => OPEN, FCO => \PostAmble_cntr_cry[7]\);
    
    \tx_packet_length_ret_0_RNIOF324[7]\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \tx_byte_cntr[9]_net_1\, B => 
        \un25_tx_byte_cntr_a_4[8]\, C => 
        \un25_tx_byte_cntr_a_4[9]\, D => \tx_byte_cntr[8]_net_1\, 
        FCI => \un25_tx_byte_cntr_1_data_tmp[3]\, S => OPEN, Y
         => OPEN, FCO => \un25_tx_byte_cntr_1_data_tmp[4]\);
    
    \tx_packet_length[8]\ : SLE
      port map(D => N_15_i, CLK => BIT_CLK, EN => 
        un1_byte_clk_en_inv_2_i, ALn => un2_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_packet_length[8]_net_1\);
    
    \PostAmble_cntr_RNIJG686[2]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => tx_state29_6_RNI9SJ61_Y, C
         => \PostAmble_cntr[2]_net_1\, D => GND_net_1, FCI => 
        \PostAmble_cntr_cry[1]\, S => \PostAmble_cntr_s[2]\, Y
         => OPEN, FCO => \PostAmble_cntr_cry[2]\);
    
    \tx_byte_cntr_cry[1]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[1]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[0]_net_1\, S => \tx_byte_cntr_s[1]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[1]_net_1\);
    
    \TX_DataEn\ : SLE
      port map(D => TX_DataEn_7, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => TX_DataEn);
    
    \tx_byte_cntr[3]\ : SLE
      port map(D => \tx_byte_cntr_s[3]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_byte_cntr[3]_net_1\);
    
    \tx_byte_cntr[7]\ : SLE
      port map(D => \tx_byte_cntr_s[7]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_byte_cntr[7]_net_1\);
    
    \tx_packet_length_ret_0_RNI8D2S[0]\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \tx_packet_length[0]_net_1\, B => 
        \un25_tx_byte_cntr_a_4[1]\, C => \tx_byte_cntr[0]_net_1\, 
        D => \tx_byte_cntr[1]_net_1\, FCI => GND_net_1, S => OPEN, 
        Y => OPEN, FCO => \un25_tx_byte_cntr_1_data_tmp[0]\);
    
    \TX_STATE[8]\ : SLE
      port map(D => \TX_STATE_64\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_STATE[8]_net_1\);
    
    \TX_SM.un25_tx_byte_cntr_a_4_cry_8\ : ARI1
      generic map(INIT => x"63B7F")

      port map(A => N_711, B => N_81, C => \TX_STATE[5]_net_1\, D
         => \tx_packet_length[9]_net_1\, FCI => 
        un25_tx_byte_cntr_a_4_cry_7, S => 
        \un25_tx_byte_cntr_a_4_i[9]\, Y => OPEN, FCO => 
        un25_tx_byte_cntr_a_4_cry_8);
    
    \txen_early_cntr_RNIDQ4JP[6]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \txen_early_cntr[6]_net_1\, C
         => \TX_STATE_RNIAIGV2_Y[7]\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[5]\, S => \txen_early_cntr_s[6]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[6]\);
    
    \TX_SM.op_eq.tx_state29_6\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \PostAmble_cntr[9]_net_1\, B => 
        \PostAmble_cntr[8]_net_1\, C => \PostAmble_cntr[7]_net_1\, 
        D => \PostAmble_cntr[6]_net_1\, Y => tx_state29_6);
    
    \txen_early_cntr_RNO[11]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \txen_early_cntr[11]_net_1\, 
        C => \TX_STATE_RNIAIGV2_Y[7]\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[10]\, S => \txen_early_cntr_s[11]\, 
        Y => OPEN, FCO => OPEN);
    
    \txen_early_cntr_RNICGS66[0]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \txen_early_cntr[0]_net_1\, C
         => \TX_STATE_RNIAIGV2_Y[7]\, D => GND_net_1, FCI => 
        txen_early_cntr_cry_cy, S => \txen_early_cntr_s[0]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[0]\);
    
    \PreAmble_cntr_RNIU58J3[1]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \PreAmble_cntr_RNIHNV31_Y[6]\, 
        C => \PreAmble_cntr[1]_net_1\, D => GND_net_1, FCI => 
        \PreAmble_cntr_cry[0]\, S => \PreAmble_cntr_s[1]\, Y => 
        OPEN, FCO => \PreAmble_cntr_cry[1]\);
    
    \TX_SM.un25_tx_byte_cntr_a_4_cry_1\ : ARI1
      generic map(INIT => x"637BF")

      port map(A => N_710, B => N_81, C => \TX_STATE[5]_net_1\, D
         => \tx_packet_length[2]_net_1\, FCI => 
        un25_tx_byte_cntr_a_4_cry_0, S => 
        \un25_tx_byte_cntr_a_4_i[2]\, Y => OPEN, FCO => 
        un25_tx_byte_cntr_a_4_cry_1);
    
    TX_STATE_68 : CFG4
      generic map(INIT => x"CA0A")

      port map(A => \TX_STATE[4]_net_1\, B => \TX_STATE[6]_net_1\, 
        C => byte_clk_en, D => N_589, Y => \TX_STATE_68\);
    
    \tx_packet_complt\ : SLE
      port map(D => \TX_STATE[0]_net_1\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => tx_packet_complt);
    
    \txen_early_cntr[0]\ : SLE
      port map(D => \txen_early_cntr_s[0]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => un2_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \txen_early_cntr[0]_net_1\);
    
    un1_TX_STATE_7_i_a2_0_a2_0_a2_0_a2 : CFG4
      generic map(INIT => x"0001")

      port map(A => \TX_STATE[2]_net_1\, B => \TX_STATE[5]_net_1\, 
        C => \TX_STATE[4]_net_1\, D => \TX_STATE[3]_net_1\, Y => 
        N_213_i);
    
    \TX_STATE_ns_8_0_.m15_e_7\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \txen_early_cntr[11]_net_1\, B => 
        \txen_early_cntr[10]_net_1\, C => 
        \txen_early_cntr[1]_net_1\, D => 
        \txen_early_cntr[0]_net_1\, Y => m15_e_7);
    
    TX_STATE_71 : CFG4
      generic map(INIT => x"FAD8")

      port map(A => byte_clk_en, B => tx_state29_6_RNI9SJ61_Y, C
         => \TX_STATE[1]_net_1\, D => \TX_STATE[2]_net_1\, Y => 
        \TX_STATE_71\);
    
    \TX_SM.un14_tx_byte_cntr_0_a2_8_a2_0_6_1\ : CFG2
      generic map(INIT => x"1")

      port map(A => \tx_byte_cntr[3]_net_1\, B => 
        \tx_byte_cntr[6]_net_1\, Y => 
        un14_tx_byte_cntr_0_a2_8_a2_0_6_1);
    
    \PreAmble_cntr[2]\ : SLE
      port map(D => \PreAmble_cntr_s[2]\, CLK => BIT_CLK, EN => 
        N_329_i, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PreAmble_cntr[2]_net_1\);
    
    \PostAmble_cntr[8]\ : SLE
      port map(D => \PostAmble_cntr_s[8]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \PostAmble_cntr[8]_net_1\);
    
    \tx_packet_length[6]\ : SLE
      port map(D => un25_tx_byte_cntr_a_4_axb_5_i, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => un2_apb3_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \tx_packet_length[6]_net_1\);
    
    \tx_byte_cntr[10]\ : SLE
      port map(D => \tx_byte_cntr_s[10]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_byte_cntr[10]_net_1\);
    
    \TX_STATE_ns_8_0_.m15_e_8\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \txen_early_cntr[5]_net_1\, B => 
        \txen_early_cntr[4]_net_1\, C => 
        \txen_early_cntr[3]_net_1\, D => 
        \txen_early_cntr[2]_net_1\, Y => m15_e_8);
    
    un1_tx_packet_length_0_sqmuxa_0_0_0_o2 : CFG3
      generic map(INIT => x"F8")

      port map(A => \TX_STATE[5]_net_1\, B => un25_tx_byte_cntr, 
        C => \TX_STATE[4]_net_1\, Y => N_719);
    
    TX_STATE_72 : CFG3
      generic map(INIT => x"5C")

      port map(A => N_1355, B => \TX_STATE[0]_net_1\, C => 
        byte_clk_en, Y => \TX_STATE_72\);
    
    \txen_early_cntr[4]\ : SLE
      port map(D => \txen_early_cntr_s[4]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => un2_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \txen_early_cntr[4]_net_1\);
    
    \PostAmble_cntr[10]\ : SLE
      port map(D => \PostAmble_cntr_s[10]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => un2_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \PostAmble_cntr[10]_net_1\);
    
    \TX_SM.un14_tx_byte_cntr_0_a2_8_a2_0_6\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \tx_byte_cntr[11]_net_1\, B => 
        \tx_byte_cntr[10]_net_1\, C => \tx_byte_cntr[5]_net_1\, D
         => un14_tx_byte_cntr_0_a2_8_a2_0_6_1, Y => 
        un14_tx_byte_cntr_0_a2_8_a2_0_6);
    
    \PreAmble_cntr_RNIS4IE[0]\ : CFG4
      generic map(INIT => x"BFFF")

      port map(A => \PreAmble_cntr[5]_net_1\, B => 
        \PreAmble_cntr[2]_net_1\, C => \PreAmble_cntr[1]_net_1\, 
        D => \PreAmble_cntr[0]_net_1\, Y => 
        PreAmble_cntr_0_sqmuxa_0_83_i_o3_4);
    
    \tx_crc_byte1_en\ : SLE
      port map(D => \TX_STATE[3]_net_1\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => tx_crc_byte1_en);
    
    \PostAmble_cntr[5]\ : SLE
      port map(D => \PostAmble_cntr_s[5]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \PostAmble_cntr[5]_net_1\);
    
    \tx_byte_cntr_cry[5]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[5]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[4]_net_1\, S => \tx_byte_cntr_s[5]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[5]_net_1\);
    
    un1_tx_packet_length_0_sqmuxa_0_0_0_a2 : CFG3
      generic map(INIT => x"C8")

      port map(A => N_81, B => \TX_STATE[5]_net_1\, C => N_80, Y
         => N_1383);
    
    \PreAmble_cntr_RNI07741[6]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => PreAmble_cntr_0_sqmuxa_0_83_i_o3_0, B => 
        PreAmble_cntr_0_sqmuxa_0_83_i_o3_4, C => 
        \PreAmble_cntr[6]_net_1\, D => TX_FIFO_Empty, Y => N_589);
    
    \TX_SM.op_eq.tx_state29_7\ : CFG4
      generic map(INIT => x"4000")

      port map(A => \PostAmble_cntr[10]_net_1\, B => 
        \PostAmble_cntr[3]_net_1\, C => \PostAmble_cntr[1]_net_1\, 
        D => \PostAmble_cntr[0]_net_1\, Y => tx_state29_7);
    
    \PostAmble_cntr[2]\ : SLE
      port map(D => \PostAmble_cntr_s[2]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \PostAmble_cntr[2]_net_1\);
    
    \un3_i_0_0_i[1]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => N_81, B => N_711, C => 
        \tx_packet_length[1]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => \un25_tx_byte_cntr_a_4_i_i[1]\);
    
    TX_STATE_65 : CFG4
      generic map(INIT => x"EEF0")

      port map(A => N_1390, B => \TX_STATE_RNIAIGV2_Y[7]\, C => 
        \TX_STATE[7]_net_1\, D => byte_clk_en, Y => \TX_STATE_65\);
    
    \TX_SM.op_eq.tx_state29_8\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \PostAmble_cntr[11]_net_1\, B => 
        \PostAmble_cntr[5]_net_1\, C => \PostAmble_cntr[4]_net_1\, 
        D => \PostAmble_cntr[2]_net_1\, Y => tx_state29_8);
    
    \PostAmble_cntr[1]\ : SLE
      port map(D => \PostAmble_cntr_s[1]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \PostAmble_cntr[1]_net_1\);
    
    \tx_packet_length_ret_0[3]\ : SLE
      port map(D => \un25_tx_byte_cntr_a_4_i[4]\, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => un2_apb3_reset_i, 
        ADn => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \un25_tx_byte_cntr_a_4[4]\);
    
    \txen_early_cntr[2]\ : SLE
      port map(D => \txen_early_cntr_s[2]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => un2_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \txen_early_cntr[2]_net_1\);
    
    \tx_packet_length[2]\ : SLE
      port map(D => un25_tx_byte_cntr_a_4_axb_1_i, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => un2_apb3_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \tx_packet_length[2]_net_1\);
    
    \txen_early_cntr_RNIUIC4J[4]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \txen_early_cntr[4]_net_1\, C
         => \TX_STATE_RNIAIGV2_Y[7]\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[3]\, S => \txen_early_cntr_s[4]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[4]\);
    
    \tx_byte_cntr_cry[6]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[6]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[5]_net_1\, S => \tx_byte_cntr_s[6]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[6]_net_1\);
    
    \TX_STATE_ns_8_0_.m72_i_i_a2_i\ : CFG4
      generic map(INIT => x"7FFF")

      port map(A => \TX_STATE[1]_net_1\, B => tx_state29_7, C => 
        tx_state29_8, D => tx_state29_6, Y => N_1355);
    
    un1_byte_clk_en_inv_2_0_0_0_2_RNIC7MU : CFG4
      generic map(INIT => x"3331")

      port map(A => \TX_STATE[5]_net_1\, B => 
        \un1_byte_clk_en_inv_2_0_0_0_2\, C => N_80, D => N_81, Y
         => un1_byte_clk_en_inv_2_i);
    
    \txen_early_cntr[7]\ : SLE
      port map(D => \txen_early_cntr_s[7]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => un2_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \txen_early_cntr[7]_net_1\);
    
    \txen_early_cntr[3]\ : SLE
      port map(D => \txen_early_cntr_s[3]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => un2_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \txen_early_cntr[3]_net_1\);
    
    \PreAmble_cntr_RNIHNV31[6]\ : ARI1
      generic map(INIT => x"4FE00")

      port map(A => \TX_STATE[6]_net_1\, B => 
        \PreAmble_cntr[6]_net_1\, C => 
        PreAmble_cntr_0_sqmuxa_0_83_i_o3_0, D => 
        PreAmble_cntr_0_sqmuxa_0_83_i_o3_4, FCI => VCC_net_1, S
         => OPEN, Y => \PreAmble_cntr_RNIHNV31_Y[6]\, FCO => 
        PreAmble_cntr_cry_cy);
    
    \PreAmble_cntr[5]\ : SLE
      port map(D => \PreAmble_cntr_s[5]\, CLK => BIT_CLK, EN => 
        N_329_i, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PreAmble_cntr[5]_net_1\);
    
    \TX_SM.un25_tx_byte_cntr_a_4_cry_2\ : ARI1
      generic map(INIT => x"637BF")

      port map(A => N_709, B => N_81, C => \TX_STATE[5]_net_1\, D
         => \tx_packet_length[3]_net_1\, FCI => 
        un25_tx_byte_cntr_a_4_cry_1, S => 
        \un25_tx_byte_cntr_a_4_i[3]\, Y => OPEN, FCO => 
        un25_tx_byte_cntr_a_4_cry_2);
    
    \tx_packet_length_RNO[8]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => N_81, B => N_705, C => 
        \tx_packet_length[8]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => N_15_i);
    
    \PostAmble_cntr_RNO[11]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => tx_state29_6_RNI9SJ61_Y, C
         => \PostAmble_cntr[11]_net_1\, D => GND_net_1, FCI => 
        \PostAmble_cntr_cry[10]\, S => \PostAmble_cntr_s[11]\, Y
         => OPEN, FCO => OPEN);
    
    \TX_STATE_RNIC0CR[6]\ : CFG3
      generic map(INIT => x"4C")

      port map(A => TX_FIFO_Empty, B => byte_clk_en, C => 
        \TX_STATE[6]_net_1\, Y => N_329_i);
    
    \PostAmble_cntr_RNIP4LVC[6]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => tx_state29_6_RNI9SJ61_Y, C
         => \PostAmble_cntr[6]_net_1\, D => GND_net_1, FCI => 
        \PostAmble_cntr_cry[5]\, S => \PostAmble_cntr_s[6]\, Y
         => OPEN, FCO => \PostAmble_cntr_cry[6]\);
    
    TX_STATE_70 : CFG3
      generic map(INIT => x"E2")

      port map(A => \TX_STATE[2]_net_1\, B => byte_clk_en, C => 
        \TX_STATE[3]_net_1\, Y => \TX_STATE_70\);
    
    \tx_packet_length_RNO[5]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => N_81, B => N_708, C => 
        \tx_packet_length[5]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => un25_tx_byte_cntr_a_4_axb_4_i);
    
    TX_STATE_67 : CFG4
      generic map(INIT => x"EAF0")

      port map(A => N_719, B => N_1336, C => \TX_STATE[5]_net_1\, 
        D => byte_clk_en, Y => \TX_STATE_67\);
    
    \tx_packet_length_RNO[7]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => N_81, B => N_706, C => 
        \tx_packet_length[7]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => un25_tx_byte_cntr_a_4_axb_6_i);
    
    \PostAmble_cntr[9]\ : SLE
      port map(D => \PostAmble_cntr_s[9]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \PostAmble_cntr[9]_net_1\);
    
    \PostAmble_cntr_RNI4UAI4[1]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => tx_state29_6_RNI9SJ61_Y, C
         => \PostAmble_cntr[1]_net_1\, D => GND_net_1, FCI => 
        \PostAmble_cntr_cry[0]\, S => \PostAmble_cntr_s[1]\, Y
         => OPEN, FCO => \PostAmble_cntr_cry[1]\);
    
    \TX_SM.un25_tx_byte_cntr_a_4_cry_3\ : ARI1
      generic map(INIT => x"637BF")

      port map(A => N_704, B => N_81, C => \TX_STATE[5]_net_1\, D
         => \tx_packet_length[4]_net_1\, FCI => 
        un25_tx_byte_cntr_a_4_cry_2, S => 
        \un25_tx_byte_cntr_a_4_i[4]\, Y => OPEN, FCO => 
        un25_tx_byte_cntr_a_4_cry_3);
    
    \tx_packet_length_RNO[9]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => N_81, B => N_711, C => 
        \tx_packet_length[9]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => N_13_i);
    
    \PostAmble_cntr_RNIOE81I[9]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => tx_state29_6_RNI9SJ61_Y, C
         => \PostAmble_cntr[9]_net_1\, D => GND_net_1, FCI => 
        \PostAmble_cntr_cry[8]\, S => \PostAmble_cntr_s[9]\, Y
         => OPEN, FCO => \PostAmble_cntr_cry[9]\);
    
    \tx_packet_length_ret_0_RNILDS25[9]\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \tx_byte_cntr[11]_net_1\, B => 
        \un25_tx_byte_cntr_a_4[10]\, C => 
        \un25_tx_byte_cntr_a_4[11]\, D => 
        \tx_byte_cntr[10]_net_1\, FCI => 
        \un25_tx_byte_cntr_1_data_tmp[4]\, S => OPEN, Y => OPEN, 
        FCO => un25_tx_byte_cntr);
    
    \PostAmble_cntr_RNIMCFS2[0]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => tx_state29_6_RNI9SJ61_Y, C
         => \PostAmble_cntr[0]_net_1\, D => GND_net_1, FCI => 
        PostAmble_cntr_cry_cy, S => \PostAmble_cntr_s[0]\, Y => 
        OPEN, FCO => \PostAmble_cntr_cry[0]\);
    
    \tx_byte_cntr[1]\ : SLE
      port map(D => \tx_byte_cntr_s[1]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_byte_cntr[1]_net_1\);
    
    \PostAmble_cntr[4]\ : SLE
      port map(D => \PostAmble_cntr_s[4]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \PostAmble_cntr[4]_net_1\);
    
    iTX_FIFO_rd_en_ret_0 : SLE
      port map(D => N_589, CLK => BIT_CLK, EN => byte_clk_en, ALn
         => un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => TX_DataEn_1_o);
    
    \TX_STATE_ns_8_0_.m16_i_0_0_a2_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => un9_start_tx_fifo_s, B => \TX_STATE[8]_net_1\, 
        Y => N_1390);
    
    TX_STATE_64 : CFG4
      generic map(INIT => x"FC70")

      port map(A => un9_start_tx_fifo_s, B => byte_clk_en, C => 
        \TX_STATE[8]_net_1\, D => \TX_STATE[0]_net_1\, Y => 
        \TX_STATE_64\);
    
    \txen_early_cntr_RNI06T101[8]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \txen_early_cntr[8]_net_1\, C
         => \TX_STATE_RNIAIGV2_Y[7]\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[7]\, S => \txen_early_cntr_s[8]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[8]\);
    
    \PreAmble_cntr[4]\ : SLE
      port map(D => \PreAmble_cntr_s[4]\, CLK => BIT_CLK, EN => 
        N_329_i, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PreAmble_cntr[4]_net_1\);
    
    TX_STATE_66 : CFG4
      generic map(INIT => x"BAF0")

      port map(A => N_1388, B => N_589, C => \TX_STATE[6]_net_1\, 
        D => byte_clk_en, Y => \TX_STATE_66\);
    
    \PreAmble_cntr[0]\ : SLE
      port map(D => \PreAmble_cntr_s[0]\, CLK => BIT_CLK, EN => 
        N_329_i, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PreAmble_cntr[0]_net_1\);
    
    \tx_packet_length_ret_0_RNIG9IL1[1]\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \tx_byte_cntr[3]_net_1\, B => 
        \un25_tx_byte_cntr_a_4[2]\, C => 
        \un25_tx_byte_cntr_a_4[3]\, D => \tx_byte_cntr[2]_net_1\, 
        FCI => \un25_tx_byte_cntr_1_data_tmp[0]\, S => OPEN, Y
         => OPEN, FCO => \un25_tx_byte_cntr_1_data_tmp[1]\);
    
    \PostAmble_cntr[0]\ : SLE
      port map(D => \PostAmble_cntr_s[0]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \PostAmble_cntr[0]_net_1\);
    
    \TX_SM.un25_tx_byte_cntr_a_4_cry_5\ : ARI1
      generic map(INIT => x"637BF")

      port map(A => N_707, B => N_81, C => \TX_STATE[5]_net_1\, D
         => \tx_packet_length[6]_net_1\, FCI => 
        un25_tx_byte_cntr_a_4_cry_4, S => 
        \un25_tx_byte_cntr_a_4_i[6]\, Y => OPEN, FCO => 
        un25_tx_byte_cntr_a_4_cry_5);
    
    iTX_FIFO_rd_en_ret_1_RNO : CFG4
      generic map(INIT => x"EEF0")

      port map(A => N_719, B => N_1383, C => 
        \un1_tx_packet_length_0_sqmuxa_o\, D => byte_clk_en, Y
         => \iTX_FIFO_rd_en_ret_1_RNO\);
    
    \tx_crc_gen\ : SLE
      port map(D => \tx_byte_cntr_cry_cy_Y[0]\, CLK => BIT_CLK, 
        EN => byte_clk_en, ALn => un2_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => tx_crc_gen);
    
    iTX_Enable_RNO : CFG1
      generic map(INIT => "01")

      port map(A => \TX_STATE[8]_net_1\, Y => \TX_STATE_i_0[8]\);
    
    \PostAmble_cntr_RNI2LCBG[8]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => tx_state29_6_RNI9SJ61_Y, C
         => \PostAmble_cntr[8]_net_1\, D => GND_net_1, FCI => 
        \PostAmble_cntr_cry[7]\, S => \PostAmble_cntr_s[8]\, Y
         => OPEN, FCO => \PostAmble_cntr_cry[8]\);
    
    \TX_STATE[4]\ : SLE
      port map(D => \TX_STATE_68\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_STATE[4]_net_1\);
    
    \tx_packet_length_ret_0[5]\ : SLE
      port map(D => \un25_tx_byte_cntr_a_4_i[6]\, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => un2_apb3_reset_i, 
        ADn => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \un25_tx_byte_cntr_a_4[6]\);
    
    \tx_packet_length[7]\ : SLE
      port map(D => un25_tx_byte_cntr_a_4_axb_6_i, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => un2_apb3_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \tx_packet_length[7]_net_1\);
    
    \TX_STATE[5]\ : SLE
      port map(D => \TX_STATE_67\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_STATE[5]_net_1\);
    
    \tx_packet_length_RNO[4]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => N_81, B => N_704, C => 
        \tx_packet_length[4]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => un25_tx_byte_cntr_a_4_axb_3_i);
    
    \tx_packet_length_ret_0_RNIOQI83[5]\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \tx_byte_cntr[7]_net_1\, B => 
        \un25_tx_byte_cntr_a_4[6]\, C => 
        \un25_tx_byte_cntr_a_4[7]\, D => \tx_byte_cntr[6]_net_1\, 
        FCI => \un25_tx_byte_cntr_1_data_tmp[2]\, S => OPEN, Y
         => OPEN, FCO => \un25_tx_byte_cntr_1_data_tmp[3]\);
    
    \txen_early_cntr[10]\ : SLE
      port map(D => \txen_early_cntr_s[10]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => un2_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \txen_early_cntr[10]_net_1\);
    
    \TX_STATE[3]\ : SLE
      port map(D => \TX_STATE_69\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_STATE[3]_net_1\);
    
    \tx_packet_length_RNO[10]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => N_81, B => N_710, C => 
        \tx_packet_length[10]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => un25_tx_byte_cntr_a_4_axb_9_i);
    
    \tx_byte_cntr_cry[9]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[9]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[8]_net_1\, S => \tx_byte_cntr_s[9]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[9]_net_1\);
    
    \TX_SM.op_eq.tx_state29_6_RNI9SJ61\ : ARI1
      generic map(INIT => x"47F00")

      port map(A => \TX_STATE[1]_net_1\, B => tx_state29_6, C => 
        tx_state29_7, D => tx_state29_8, FCI => VCC_net_1, S => 
        OPEN, Y => tx_state29_6_RNI9SJ61_Y, FCO => 
        PostAmble_cntr_cry_cy);
    
    \PostAmble_cntr_RNIKOTJ9[4]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => tx_state29_6_RNI9SJ61_Y, C
         => \PostAmble_cntr[4]_net_1\, D => GND_net_1, FCI => 
        \PostAmble_cntr_cry[3]\, S => \PostAmble_cntr_s[4]\, Y
         => OPEN, FCO => \PostAmble_cntr_cry[4]\);
    
    \TX_SM.un14_tx_byte_cntr_0_a2_8_a2_0\ : CFG3
      generic map(INIT => x"02")

      port map(A => \tx_byte_cntr[2]_net_1\, B => 
        \tx_byte_cntr[1]_net_1\, C => \tx_byte_cntr[0]_net_1\, Y
         => N_1447);
    
    TX_IDLE_LINE_DETECTOR : IdleLineDetector_0
      port map(manches_in_dly(1) => manches_in_dly(1), 
        manches_in_dly(0) => manches_in_dly(0), idle_line5 => 
        idle_line5, CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, 
        un2_apb3_reset_i => un2_apb3_reset_i, tx_idle_line => 
        tx_idle_line);
    
    tx_idle_line_s : SLE
      port map(D => tx_idle_line, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_idle_line_s\);
    
    \tx_packet_length[0]\ : SLE
      port map(D => N_19_i, CLK => BIT_CLK, EN => 
        un1_byte_clk_en_inv_2_i, ALn => un2_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_packet_length[0]_net_1\);
    
    \TX_SM.un9_start_tx_fifo_s\ : CFG2
      generic map(INIT => x"8")

      port map(A => \start_tx_FIFO_s\, B => \tx_idle_line_s\, Y
         => un9_start_tx_fifo_s);
    
    \TX_SM.un14_tx_byte_cntr_0_a2_8_a2\ : CFG3
      generic map(INIT => x"80")

      port map(A => un14_tx_byte_cntr_0_a2_8_a2_0_6, B => N_1447, 
        C => un14_tx_byte_cntr_0_a2_8_a2_0_5, Y => N_81);
    
    \txen_early_cntr[6]\ : SLE
      port map(D => \txen_early_cntr_s[6]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => un2_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \txen_early_cntr[6]_net_1\);
    
    \PostAmble_cntr[7]\ : SLE
      port map(D => \PostAmble_cntr_s[7]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \PostAmble_cntr[7]_net_1\);
    
    \tx_packet_length_ret_0[2]\ : SLE
      port map(D => \un25_tx_byte_cntr_a_4_i[3]\, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => un2_apb3_reset_i, 
        ADn => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \un25_tx_byte_cntr_a_4[3]\);
    
    \tx_byte_cntr[9]\ : SLE
      port map(D => \tx_byte_cntr_s[9]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_byte_cntr[9]_net_1\);
    
    \tx_packet_length_ret_0[9]\ : SLE
      port map(D => \un25_tx_byte_cntr_a_4_i[10]\, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => un2_apb3_reset_i, 
        ADn => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \un25_tx_byte_cntr_a_4[10]\);
    
    \tx_byte_cntr_cry[8]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[8]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[7]_net_1\, S => \tx_byte_cntr_s[8]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[8]_net_1\);
    
    \TX_SM.un25_tx_byte_cntr_a_4_cry_9\ : ARI1
      generic map(INIT => x"63B7F")

      port map(A => N_710, B => N_81, C => \TX_STATE[5]_net_1\, D
         => \tx_packet_length[10]_net_1\, FCI => 
        un25_tx_byte_cntr_a_4_cry_8, S => 
        \un25_tx_byte_cntr_a_4_i[10]\, Y => OPEN, FCO => 
        un25_tx_byte_cntr_a_4_cry_9);
    
    \tx_byte_cntr_cry[3]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[3]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[2]_net_1\, S => \tx_byte_cntr_s[3]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[3]_net_1\);
    
    \PostAmble_cntr[3]\ : SLE
      port map(D => \PostAmble_cntr_s[3]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \PostAmble_cntr[3]_net_1\);
    
    \txen_early_cntr_RNIMVGQS[7]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \txen_early_cntr[7]_net_1\, C
         => \TX_STATE_RNIAIGV2_Y[7]\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[6]\, S => \txen_early_cntr_s[7]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[7]\);
    
    \TX_SM.un25_tx_byte_cntr_a_4_cry_0\ : ARI1
      generic map(INIT => x"637BF")

      port map(A => N_711, B => N_81, C => \TX_STATE[5]_net_1\, D
         => \tx_packet_length[1]_net_1\, FCI => GND_net_1, S => 
        OPEN, Y => un25_tx_byte_cntr_a_4_cry_0_Y, FCO => 
        un25_tx_byte_cntr_a_4_cry_0);
    
    \TX_STATE[6]\ : SLE
      port map(D => \TX_STATE_66\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_STATE[6]_net_1\);
    
    \tx_preamble_pat_en\ : SLE
      port map(D => TX_DataEn_1_m, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => tx_preamble_pat_en);
    
    \TX_STATE[1]\ : SLE
      port map(D => \TX_STATE_71\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_STATE[1]_net_1\);
    
    \TX_SM.un9_tx_byte_cntr_0_a2_0_a2\ : CFG3
      generic map(INIT => x"80")

      port map(A => un14_tx_byte_cntr_0_a2_8_a2_0_6, B => N_957, 
        C => un14_tx_byte_cntr_0_a2_8_a2_0_5, Y => N_80);
    
    \PreAmble_cntr_RNIMESQ4[2]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \PreAmble_cntr_RNIHNV31_Y[6]\, 
        C => \PreAmble_cntr[2]_net_1\, D => GND_net_1, FCI => 
        \PreAmble_cntr_cry[1]\, S => \PreAmble_cntr_s[2]\, Y => 
        OPEN, FCO => \PreAmble_cntr_cry[2]\);
    
    \TX_STATE_ns_8_0_.m56_i_0_0_a2_0\ : CFG3
      generic map(INIT => x"40")

      port map(A => \tx_byte_cntr[2]_net_1\, B => 
        \tx_byte_cntr[1]_net_1\, C => \tx_byte_cntr[0]_net_1\, Y
         => N_957);
    
    \tx_packet_length_ret_0_RNI0E2F2[3]\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \tx_byte_cntr[5]_net_1\, B => 
        \un25_tx_byte_cntr_a_4[4]\, C => 
        \un25_tx_byte_cntr_a_4[5]\, D => \tx_byte_cntr[4]_net_1\, 
        FCI => \un25_tx_byte_cntr_1_data_tmp[1]\, S => OPEN, Y
         => OPEN, FCO => \un25_tx_byte_cntr_1_data_tmp[2]\);
    
    \tx_packet_length_ret_0[8]\ : SLE
      port map(D => \un25_tx_byte_cntr_a_4_i[9]\, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => un2_apb3_reset_i, 
        ADn => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \un25_tx_byte_cntr_a_4[9]\);
    
    \txen_early_cntr[11]\ : SLE
      port map(D => \txen_early_cntr_s[11]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => un2_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \txen_early_cntr[11]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity ManchesEncoder is

    port( manches_in_dly                  : in    std_logic_vector(1 downto 0);
          start_tx_FIFO                   : in    std_logic;
          un1_tx_packet_length_0_sqmuxa_o : out   std_logic;
          TX_DataEn_1_o                   : out   std_logic;
          TX_FIFO_Empty                   : in    std_logic;
          idle_line5                      : out   std_logic;
          tx_col_detect_en                : out   std_logic;
          CommsFPGA_CCC_0_GL0             : in    std_logic;
          DRVR_EN_c                       : out   std_logic;
          internal_loopback               : in    std_logic;
          external_loopback               : in    std_logic;
          tx_packet_complt                : out   std_logic;
          un2_apb3_reset                  : in    std_logic;
          N_706                           : in    std_logic;
          N_704                           : in    std_logic;
          N_709                           : in    std_logic;
          N_708                           : in    std_logic;
          N_707                           : in    std_logic;
          N_710                           : in    std_logic;
          N_711                           : in    std_logic;
          N_705                           : in    std_logic;
          TX_PreAmble                     : out   std_logic;
          CommsFPGA_CCC_0_GL1             : in    std_logic;
          byte_clk_en                     : in    std_logic;
          BIT_CLK                         : in    std_logic;
          un2_apb3_reset_i                : in    std_logic;
          MANCH_OUT_P_c_i                 : out   std_logic;
          MANCH_OUT_P_c                   : out   std_logic
        );

end ManchesEncoder;

architecture DEF_ARCH of ManchesEncoder is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CRC16_Generator_0
    port( tx_crc_data    : out   std_logic_vector(15 downto 0);
          N_705          : in    std_logic := 'U';
          N_709          : in    std_logic := 'U';
          N_710          : in    std_logic := 'U';
          N_711          : in    std_logic := 'U';
          N_704          : in    std_logic := 'U';
          N_707          : in    std_logic := 'U';
          N_708          : in    std_logic := 'U';
          N_706          : in    std_logic := 'U';
          tx_crc_gen     : in    std_logic := 'U';
          byte_clk_en    : in    std_logic := 'U';
          BIT_CLK        : in    std_logic := 'U';
          tx_crc_reset_i : in    std_logic := 'U'
        );
  end component;

  component TX_Collision_Detector
    port( un2_apb3_reset      : in    std_logic := 'U';
          external_loopback   : in    std_logic := 'U';
          internal_loopback   : in    std_logic := 'U';
          DRVR_EN_c           : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          tx_col_detect_en    : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component TX_SM
    port( manches_in_dly                  : in    std_logic_vector(1 downto 0) := (others => 'U');
          CommsFPGA_CCC_0_GL0             : in    std_logic := 'U';
          idle_line5                      : out   std_logic;
          TX_FIFO_Empty                   : in    std_logic := 'U';
          N_705                           : in    std_logic := 'U';
          N_706                           : in    std_logic := 'U';
          N_707                           : in    std_logic := 'U';
          N_708                           : in    std_logic := 'U';
          N_704                           : in    std_logic := 'U';
          N_709                           : in    std_logic := 'U';
          N_710                           : in    std_logic := 'U';
          N_711                           : in    std_logic := 'U';
          TX_DataEn                       : out   std_logic;
          TX_PreAmble                     : out   std_logic;
          tx_crc_byte1_en                 : out   std_logic;
          tx_crc_byte2_en                 : out   std_logic;
          tx_packet_complt                : out   std_logic;
          tx_crc_gen                      : out   std_logic;
          TX_DataEn_1_o                   : out   std_logic;
          un1_tx_packet_length_0_sqmuxa_o : out   std_logic;
          start_tx_FIFO                   : in    std_logic := 'U';
          DRVR_EN_c                       : out   std_logic;
          byte_clk_en                     : in    std_logic := 'U';
          tx_preamble_pat_en              : out   std_logic;
          BIT_CLK                         : in    std_logic := 'U';
          un2_apb3_reset_i                : in    std_logic := 'U'
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal tx_crc_reset_i, \tx_crc_reset\, \MANCH_OUT_P_c\, 
        \p2s_data[5]_net_1\, VCC_net_1, \p2s_data_9[5]\, 
        GND_net_1, \p2s_data[6]_net_1\, N_403_i, 
        \p2s_data[7]_net_1\, N_402_i, \byte_clk_en_d[0]_net_1\, 
        \TX_PreAmble_d[0]_net_1\, \TX_PreAmble\, 
        \TX_PreAmble_d[1]_net_1\, \p2s_data[0]_net_1\, N_406_i, 
        \p2s_data[1]_net_1\, \p2s_data_9[1]\, \p2s_data[2]_net_1\, 
        N_405_i, \p2s_data[3]_net_1\, \p2s_data_9[3]\, 
        \p2s_data[4]_net_1\, N_404_i, \TX_DataEn_d1\, TX_DataEn, 
        MANCHESTER_OUT_5, tx_preamble_pat_en, N_455, 
        tx_crc_byte1_en, \p2s_data_9_i_0_m2_1_1[0]\, N_1417, 
        N_642, \tx_crc_data[8]\, \tx_crc_data[0]\, 
        \p2s_data_9_m2_1_0[1]\, \p2s_data_9_m2[1]\, 
        \tx_crc_data[1]\, N_44_1, \p2s_data_9_m2_1_0[2]\, 
        \p2s_data_9_m2[2]\, \tx_crc_data[2]\, 
        \p2s_data_9_m2_1_0[6]\, \p2s_data_9_m2[6]\, 
        \tx_crc_data[6]\, \p2s_data_9_m2_1_0[5]\, 
        \p2s_data_9_m2[5]\, \tx_crc_data[5]\, 
        \p2s_data_9_m2_1_0[3]\, \p2s_data_9_m2[3]\, 
        \tx_crc_data[3]\, \p2s_data_9_m2_1_0[4]\, 
        \p2s_data_9_m2[4]\, \tx_crc_data[4]\, 
        \p2s_data_9_m2_1_0[7]\, \p2s_data_9_m2[7]\, 
        \tx_crc_data[7]\, un24_tx_dataen, N_538, N_1329, 
        \un1_TX_PreAmble_d_i[0]\, tx_crc_byte2_en, 
        \tx_packet_complt\, N_1472, N_544, \tx_crc_data[9]\, 
        \tx_crc_data[11]\, \tx_crc_data[13]\, \tx_crc_data[12]\, 
        \tx_crc_data[10]\, \tx_crc_data[15]\, \tx_crc_data[14]\, 
        \DRVR_EN_c\, tx_crc_gen : std_logic;

    for all : CRC16_Generator_0
	Use entity work.CRC16_Generator_0(DEF_ARCH);
    for all : TX_Collision_Detector
	Use entity work.TX_Collision_Detector(DEF_ARCH);
    for all : TX_SM
	Use entity work.TX_SM(DEF_ARCH);
begin 

    DRVR_EN_c <= \DRVR_EN_c\;
    tx_packet_complt <= \tx_packet_complt\;
    TX_PreAmble <= \TX_PreAmble\;
    MANCH_OUT_P_c <= \MANCH_OUT_P_c\;

    \byte_clk_en_d[0]\ : SLE
      port map(D => byte_clk_en, CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \byte_clk_en_d[0]_net_1\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_m2[3]\ : CFG4
      generic map(INIT => x"EA51")

      port map(A => N_455, B => N_1417, C => N_709, D => 
        \p2s_data_9_m2_1_0[3]\, Y => \p2s_data_9_m2[3]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_0_1[3]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => N_1472, B => \tx_crc_data[11]\, C => 
        \p2s_data_9_m2[3]\, D => N_544, Y => \p2s_data_9[3]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_m2_1_0[4]\ : CFG4
      generic map(INIT => x"0C55")

      port map(A => \tx_crc_data[4]\, B => \p2s_data[3]_net_1\, C
         => N_44_1, D => N_455, Y => \p2s_data_9_m2_1_0[4]\);
    
    \TX_PreAmble_d[0]\ : SLE
      port map(D => \TX_PreAmble\, CLK => CommsFPGA_CCC_0_GL1, EN
         => VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \TX_PreAmble_d[0]_net_1\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_m2_1_0[5]\ : CFG4
      generic map(INIT => x"0C55")

      port map(A => \tx_crc_data[5]\, B => \p2s_data[4]_net_1\, C
         => N_44_1, D => N_455, Y => \p2s_data_9_m2_1_0[5]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_0_1[5]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => N_1472, B => \tx_crc_data[13]\, C => 
        \p2s_data_9_m2[5]\, D => N_544, Y => \p2s_data_9[5]\);
    
    \PARALLEL_2_SERIAL_PROC.un5_tx_dataen_i_o2_1_o2_1_o2\ : CFG4
      generic map(INIT => x"73FF")

      port map(A => tx_preamble_pat_en, B => TX_DataEn, C => 
        \TX_PreAmble_d[1]_net_1\, D => \byte_clk_en_d[0]_net_1\, 
        Y => N_455);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_m2[4]\ : CFG4
      generic map(INIT => x"EA51")

      port map(A => N_455, B => N_1417, C => N_704, D => 
        \p2s_data_9_m2_1_0[4]\, Y => \p2s_data_9_m2[4]\);
    
    \un1_TX_PreAmble_d_0_o2_0_o2_0_o2[0]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => N_1329, B => \TX_PreAmble\, C => 
        tx_preamble_pat_en, Y => \un1_TX_PreAmble_d_i[0]\);
    
    \p2s_data[0]\ : SLE
      port map(D => N_406_i, CLK => BIT_CLK, EN => VCC_net_1, ALn
         => un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \p2s_data[0]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \p2s_data[6]\ : SLE
      port map(D => N_403_i, CLK => BIT_CLK, EN => VCC_net_1, ALn
         => un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \p2s_data[6]_net_1\);
    
    \MAN_OUT_DATA_PROC.un24_tx_dataen\ : CFG2
      generic map(INIT => x"E")

      port map(A => TX_DataEn, B => \TX_DataEn_d1\, Y => 
        un24_tx_dataen);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_ss0_i_0_0_1\ : CFG4
      generic map(INIT => x"AB03")

      port map(A => \byte_clk_en_d[0]_net_1\, B => TX_DataEn, C
         => \TX_PreAmble\, D => N_1329, Y => N_44_1);
    
    tx_crc_reset_RNI5CLE : CLKINT
      port map(A => \tx_crc_reset\, Y => tx_crc_reset_i);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_i_0_0_o2[7]\ : CFG4
      generic map(INIT => x"5FDF")

      port map(A => TX_DataEn, B => N_538, C => 
        \byte_clk_en_d[0]_net_1\, D => tx_preamble_pat_en, Y => 
        N_544);
    
    TX_CRC_GEN_INST : CRC16_Generator_0
      port map(tx_crc_data(15) => \tx_crc_data[15]\, 
        tx_crc_data(14) => \tx_crc_data[14]\, tx_crc_data(13) => 
        \tx_crc_data[13]\, tx_crc_data(12) => \tx_crc_data[12]\, 
        tx_crc_data(11) => \tx_crc_data[11]\, tx_crc_data(10) => 
        \tx_crc_data[10]\, tx_crc_data(9) => \tx_crc_data[9]\, 
        tx_crc_data(8) => \tx_crc_data[8]\, tx_crc_data(7) => 
        \tx_crc_data[7]\, tx_crc_data(6) => \tx_crc_data[6]\, 
        tx_crc_data(5) => \tx_crc_data[5]\, tx_crc_data(4) => 
        \tx_crc_data[4]\, tx_crc_data(3) => \tx_crc_data[3]\, 
        tx_crc_data(2) => \tx_crc_data[2]\, tx_crc_data(1) => 
        \tx_crc_data[1]\, tx_crc_data(0) => \tx_crc_data[0]\, 
        N_705 => N_705, N_709 => N_709, N_710 => N_710, N_711 => 
        N_711, N_704 => N_704, N_707 => N_707, N_708 => N_708, 
        N_706 => N_706, tx_crc_gen => tx_crc_gen, byte_clk_en => 
        byte_clk_en, BIT_CLK => BIT_CLK, tx_crc_reset_i => 
        tx_crc_reset_i);
    
    TX_COLLISION_DETECTOR_INST : TX_Collision_Detector
      port map(un2_apb3_reset => un2_apb3_reset, 
        external_loopback => external_loopback, internal_loopback
         => internal_loopback, DRVR_EN_c => \DRVR_EN_c\, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, 
        tx_col_detect_en => tx_col_detect_en);
    
    \p2s_data[2]\ : SLE
      port map(D => N_405_i, CLK => BIT_CLK, EN => VCC_net_1, ALn
         => un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \p2s_data[2]_net_1\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_m2[7]\ : CFG4
      generic map(INIT => x"EA51")

      port map(A => N_455, B => N_1417, C => N_706, D => 
        \p2s_data_9_m2_1_0[7]\, Y => \p2s_data_9_m2[7]\);
    
    \MAN_OUT_DATA_PROC.MANCHESTER_OUT_5_u\ : CFG4
      generic map(INIT => x"5A78")

      port map(A => BIT_CLK, B => \un1_TX_PreAmble_d_i[0]\, C => 
        \p2s_data[7]_net_1\, D => un24_tx_dataen, Y => 
        MANCHESTER_OUT_5);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_ss0_i_0_a2_3\ : CFG3
      generic map(INIT => x"40")

      port map(A => tx_crc_byte2_en, B => 
        \byte_clk_en_d[0]_net_1\, C => TX_DataEn, Y => N_1417);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_i_0_m2_1_1[0]\ : CFG3
      generic map(INIT => x"27")

      port map(A => tx_crc_byte1_en, B => \tx_crc_data[8]\, C => 
        \tx_crc_data[0]\, Y => \p2s_data_9_i_0_m2_1_1[0]\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_m2_1_0[2]\ : CFG4
      generic map(INIT => x"0C55")

      port map(A => \tx_crc_data[2]\, B => \p2s_data[1]_net_1\, C
         => N_44_1, D => N_455, Y => \p2s_data_9_m2_1_0[2]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_m2_1_0[6]\ : CFG4
      generic map(INIT => x"0C55")

      port map(A => \tx_crc_data[6]\, B => \p2s_data[5]_net_1\, C
         => N_44_1, D => N_455, Y => \p2s_data_9_m2_1_0[6]\);
    
    \p2s_data_RNO[6]\ : CFG4
      generic map(INIT => x"D0DD")

      port map(A => N_1472, B => \tx_crc_data[14]\, C => 
        \p2s_data_9_m2[6]\, D => N_544, Y => N_403_i);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_m2_1_0[1]\ : CFG4
      generic map(INIT => x"0C55")

      port map(A => \tx_crc_data[1]\, B => \p2s_data[0]_net_1\, C
         => N_44_1, D => N_455, Y => \p2s_data_9_m2_1_0[1]\);
    
    \p2s_data[4]\ : SLE
      port map(D => N_404_i, CLK => BIT_CLK, EN => VCC_net_1, ALn
         => un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \p2s_data[4]_net_1\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_i_0_0_m2[0]\ : CFG4
      generic map(INIT => x"7323")

      port map(A => tx_crc_byte1_en, B => 
        \p2s_data_9_i_0_m2_1_1[0]\, C => N_1417, D => N_705, Y
         => N_642);
    
    TRANSMIT_SM : TX_SM
      port map(manches_in_dly(1) => manches_in_dly(1), 
        manches_in_dly(0) => manches_in_dly(0), 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, idle_line5
         => idle_line5, TX_FIFO_Empty => TX_FIFO_Empty, N_705 => 
        N_705, N_706 => N_706, N_707 => N_707, N_708 => N_708, 
        N_704 => N_704, N_709 => N_709, N_710 => N_710, N_711 => 
        N_711, TX_DataEn => TX_DataEn, TX_PreAmble => 
        \TX_PreAmble\, tx_crc_byte1_en => tx_crc_byte1_en, 
        tx_crc_byte2_en => tx_crc_byte2_en, tx_packet_complt => 
        \tx_packet_complt\, tx_crc_gen => tx_crc_gen, 
        TX_DataEn_1_o => TX_DataEn_1_o, 
        un1_tx_packet_length_0_sqmuxa_o => 
        un1_tx_packet_length_0_sqmuxa_o, start_tx_FIFO => 
        start_tx_FIFO, DRVR_EN_c => \DRVR_EN_c\, byte_clk_en => 
        byte_clk_en, tx_preamble_pat_en => tx_preamble_pat_en, 
        BIT_CLK => BIT_CLK, un2_apb3_reset_i => un2_apb3_reset_i);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_m2_1_0[7]\ : CFG4
      generic map(INIT => x"0C55")

      port map(A => \tx_crc_data[7]\, B => \p2s_data[6]_net_1\, C
         => N_44_1, D => N_455, Y => \p2s_data_9_m2_1_0[7]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_m2[2]\ : CFG4
      generic map(INIT => x"EA51")

      port map(A => N_455, B => N_1417, C => N_710, D => 
        \p2s_data_9_m2_1_0[2]\, Y => \p2s_data_9_m2[2]\);
    
    \p2s_data_RNO[2]\ : CFG4
      generic map(INIT => x"D0DD")

      port map(A => N_1472, B => \tx_crc_data[10]\, C => 
        \p2s_data_9_m2[2]\, D => N_544, Y => N_405_i);
    
    \p2s_data_RNO[4]\ : CFG4
      generic map(INIT => x"D0DD")

      port map(A => N_1472, B => \tx_crc_data[12]\, C => 
        \p2s_data_9_m2[4]\, D => N_544, Y => N_404_i);
    
    \p2s_data[1]\ : SLE
      port map(D => \p2s_data_9[1]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \p2s_data[1]_net_1\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_m2_1_0[3]\ : CFG4
      generic map(INIT => x"0C55")

      port map(A => \tx_crc_data[3]\, B => \p2s_data[2]_net_1\, C
         => N_44_1, D => N_455, Y => \p2s_data_9_m2_1_0[3]\);
    
    \p2s_data_RNO[0]\ : CFG3
      generic map(INIT => x"32")

      port map(A => tx_preamble_pat_en, B => N_455, C => N_642, Y
         => N_406_i);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_i_0_o2_0[7]\ : CFG2
      generic map(INIT => x"D")

      port map(A => tx_crc_byte1_en, B => 
        \TX_PreAmble_d[1]_net_1\, Y => N_538);
    
    \p2s_data[3]\ : SLE
      port map(D => \p2s_data_9[3]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \p2s_data[3]_net_1\);
    
    MANCHESTER_OUT : SLE
      port map(D => MANCHESTER_OUT_5, CLK => CommsFPGA_CCC_0_GL1, 
        EN => VCC_net_1, ALn => un2_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \MANCH_OUT_P_c\);
    
    \TX_PreAmble_d[1]\ : SLE
      port map(D => \TX_PreAmble_d[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL1, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \TX_PreAmble_d[1]_net_1\);
    
    MANCHESTER_OUT_RNI19ND : CFG1
      generic map(INIT => "01")

      port map(A => \MANCH_OUT_P_c\, Y => MANCH_OUT_P_c_i);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_m2[5]\ : CFG4
      generic map(INIT => x"EA51")

      port map(A => N_455, B => N_1417, C => N_708, D => 
        \p2s_data_9_m2_1_0[5]\, Y => \p2s_data_9_m2[5]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_ss0_i_0_a2_5\ : CFG2
      generic map(INIT => x"4")

      port map(A => tx_preamble_pat_en, B => 
        \TX_PreAmble_d[1]_net_1\, Y => N_1329);
    
    \p2s_data[5]\ : SLE
      port map(D => \p2s_data_9[5]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \p2s_data[5]_net_1\);
    
    TX_DataEn_d1 : SLE
      port map(D => TX_DataEn, CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_DataEn_d1\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_0_1[1]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => N_1472, B => \tx_crc_data[9]\, C => 
        \p2s_data_9_m2[1]\, D => N_544, Y => \p2s_data_9[1]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_i_0_a2_3[7]\ : CFG4
      generic map(INIT => x"0020")

      port map(A => TX_DataEn, B => N_538, C => 
        \byte_clk_en_d[0]_net_1\, D => tx_preamble_pat_en, Y => 
        N_1472);
    
    tx_crc_reset : CFG2
      generic map(INIT => x"1")

      port map(A => un2_apb3_reset, B => \tx_packet_complt\, Y
         => \tx_crc_reset\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_m2[1]\ : CFG4
      generic map(INIT => x"EA51")

      port map(A => N_455, B => N_1417, C => N_711, D => 
        \p2s_data_9_m2_1_0[1]\, Y => \p2s_data_9_m2[1]\);
    
    \p2s_data_RNO[7]\ : CFG4
      generic map(INIT => x"D0DD")

      port map(A => N_1472, B => \tx_crc_data[15]\, C => 
        \p2s_data_9_m2[7]\, D => N_544, Y => N_402_i);
    
    \p2s_data[7]\ : SLE
      port map(D => N_402_i, CLK => BIT_CLK, EN => VCC_net_1, ALn
         => un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \p2s_data[7]_net_1\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_m2[6]\ : CFG4
      generic map(INIT => x"EA51")

      port map(A => N_455, B => N_1417, C => N_707, D => 
        \p2s_data_9_m2_1_0[6]\, Y => \p2s_data_9_m2[6]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity IdleLineDetector_1 is

    port( idle_line5          : in    std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          un2_apb3_reset_i    : in    std_logic;
          idle_line           : out   std_logic
        );

end IdleLineDetector_1;

architecture DEF_ARCH of IdleLineDetector_1 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, N_149_i, GND_net_1, 
        \idle_line_cntr[0]_net_1\, \idle_line_cntr_s[0]\, 
        \idle_line_cntr[1]_net_1\, \idle_line_cntr_s[1]\, 
        \idle_line_cntr[2]_net_1\, \idle_line_cntr_s[2]\, 
        \idle_line_cntr[3]_net_1\, \idle_line_cntr_s[3]\, 
        \idle_line_cntr[4]_net_1\, \idle_line_cntr_s[4]\, 
        \idle_line_cntr[5]_net_1\, \idle_line_cntr_s[5]\, 
        \idle_line_cntr[6]_net_1\, \idle_line_cntr_s[6]\, 
        \idle_line_cntr[7]_net_1\, \idle_line_cntr_s[7]\, 
        \idle_line_cntr[8]_net_1\, \idle_line_cntr_s[8]\, 
        \idle_line_cntr[9]_net_1\, \idle_line_cntr_s[9]\, 
        \idle_line_cntr[10]_net_1\, \idle_line_cntr_s[10]\, 
        \idle_line_cntr[11]_net_1\, \idle_line_cntr_s[11]\, 
        \idle_line_cntr[12]_net_1\, \idle_line_cntr_s[12]\, 
        \idle_line_cntr[13]_net_1\, \idle_line_cntr_s[13]\, 
        \idle_line_cntr[14]_net_1\, \idle_line_cntr_s[14]\, 
        \idle_line_cntr[15]_net_1\, \idle_line_cntr_s[15]\, 
        idle_line_cntr_cry_cy, un5_manches_in_dly_9_RNINM8S_Y, 
        un5_manches_in_dly_9, un5_manches_in_dly_10, 
        un5_manches_in_dly_11, \idle_line_cntr_cry[0]\, 
        \idle_line_cntr_cry[1]\, \idle_line_cntr_cry[2]\, 
        \idle_line_cntr_cry[3]\, \idle_line_cntr_cry[4]\, 
        \idle_line_cntr_cry[5]\, \idle_line_cntr_cry[6]\, 
        \idle_line_cntr_cry[7]\, \idle_line_cntr_cry[8]\, 
        \idle_line_cntr_cry[9]\, \idle_line_cntr_cry[10]\, 
        \idle_line_cntr_cry[11]\, \idle_line_cntr_cry[12]\, 
        \idle_line_cntr_cry[13]\, \idle_line_cntr_cry[14]\, 
        un5_manches_in_dly_8 : std_logic;

begin 


    \idle_line\ : SLE
      port map(D => N_149_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        idle_line);
    
    \IDLE_LINE_DETECT_PROC.un5_manches_in_dly_11\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \idle_line_cntr[11]_net_1\, B => 
        \idle_line_cntr[8]_net_1\, C => \idle_line_cntr[7]_net_1\, 
        D => un5_manches_in_dly_8, Y => un5_manches_in_dly_11);
    
    \idle_line_cntr_RNILB687[6]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[6]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[5]\, S => \idle_line_cntr_s[6]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[6]\);
    
    \idle_line_cntr_RNIBRPHF[12]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[12]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[11]\, S => \idle_line_cntr_s[12]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[12]\);
    
    \idle_line_cntr_RNI24F29[8]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[8]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[7]\, S => \idle_line_cntr_s[8]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[8]\);
    
    \idle_line_cntr[4]\ : SLE
      port map(D => \idle_line_cntr_s[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[4]_net_1\);
    
    \idle_line_cntr[14]\ : SLE
      port map(D => \idle_line_cntr_s[14]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[14]_net_1\);
    
    \idle_line_cntr_RNIM0HM2[1]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[1]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[0]\, S => \idle_line_cntr_s[1]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[1]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \idle_line_cntr_RNI9689E[11]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[11]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[10]\, S => \idle_line_cntr_s[11]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[11]\);
    
    \IDLE_LINE_DETECT_PROC.un5_manches_in_dly_9\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \idle_line_cntr[10]_net_1\, B => 
        \idle_line_cntr[9]_net_1\, C => \idle_line_cntr[2]_net_1\, 
        D => \idle_line_cntr[1]_net_1\, Y => un5_manches_in_dly_9);
    
    \IDLE_LINE_DETECT_PROC.un5_manches_in_dly_10\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \idle_line_cntr[6]_net_1\, B => 
        \idle_line_cntr[5]_net_1\, C => \idle_line_cntr[4]_net_1\, 
        D => \idle_line_cntr[3]_net_1\, Y => 
        un5_manches_in_dly_10);
    
    \idle_line_cntr_RNICNTD5[4]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[4]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[3]\, S => \idle_line_cntr_s[4]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[4]\);
    
    \idle_line_cntr[9]\ : SLE
      port map(D => \idle_line_cntr_s[9]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[9]_net_1\);
    
    \idle_line_cntr[8]\ : SLE
      port map(D => \idle_line_cntr_s[8]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[8]_net_1\);
    
    \idle_line_cntr[7]\ : SLE
      port map(D => \idle_line_cntr_s[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[7]_net_1\);
    
    \idle_line_cntr[15]\ : SLE
      port map(D => \idle_line_cntr_s[15]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[15]_net_1\);
    
    \idle_line_cntr[11]\ : SLE
      port map(D => \idle_line_cntr_s[11]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[11]_net_1\);
    
    \idle_line_cntr[10]\ : SLE
      port map(D => \idle_line_cntr_s[10]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[10]_net_1\);
    
    \idle_line_cntr_RNIEHBQG[13]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[13]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[12]\, S => \idle_line_cntr_s[13]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[13]\);
    
    \idle_line_cntr[1]\ : SLE
      port map(D => \idle_line_cntr_s[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[1]_net_1\);
    
    \IDLE_LINE_DETECT_PROC.un5_manches_in_dly_8\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \idle_line_cntr[15]_net_1\, B => 
        \idle_line_cntr[14]_net_1\, C => 
        \idle_line_cntr[13]_net_1\, D => 
        \idle_line_cntr[12]_net_1\, Y => un5_manches_in_dly_8);
    
    \idle_line_cntr_RNO[15]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[15]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[14]\, S => \idle_line_cntr_s[15]\, Y
         => OPEN, FCO => OPEN);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \idle_line_cntr_RNI8IM0D[10]\ : ARI1
      generic map(INIT => x"4D800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[10]_net_1\, D => N_149_i, FCI => 
        \idle_line_cntr_cry[9]\, S => \idle_line_cntr_s[10]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[10]\);
    
    \idle_line_cntr_RNI77LJ3[2]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[2]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[1]\, S => \idle_line_cntr_s[2]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[2]\);
    
    \IDLE_LINE_DETECT_PROC.un5_manches_in_dly_9_RNINM8S\ : ARI1
      generic map(INIT => x"4007F")

      port map(A => idle_line5, B => un5_manches_in_dly_9, C => 
        un5_manches_in_dly_10, D => un5_manches_in_dly_11, FCI
         => VCC_net_1, S => OPEN, Y => 
        un5_manches_in_dly_9_RNINM8S_Y, FCO => 
        idle_line_cntr_cry_cy);
    
    \idle_line_cntr_RNI6RCP1[0]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[0]_net_1\, D => GND_net_1, FCI => 
        idle_line_cntr_cry_cy, S => \idle_line_cntr_s[0]\, Y => 
        OPEN, FCO => \idle_line_cntr_cry[0]\);
    
    \IDLE_LINE_DETECT_PROC.un5_manches_in_dly_9_RNINM8S_0\ : CFG4
      generic map(INIT => x"0800")

      port map(A => un5_manches_in_dly_10, B => 
        un5_manches_in_dly_9, C => idle_line5, D => 
        un5_manches_in_dly_11, Y => N_149_i);
    
    \idle_line_cntr_RNII8T2I[14]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[14]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[13]\, S => \idle_line_cntr_s[14]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[14]\);
    
    \idle_line_cntr[6]\ : SLE
      port map(D => \idle_line_cntr_s[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[6]_net_1\);
    
    \idle_line_cntr_RNIPEPG4[3]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[3]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[2]\, S => \idle_line_cntr_s[3]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[3]\);
    
    \idle_line_cntr[13]\ : SLE
      port map(D => \idle_line_cntr_s[13]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[13]_net_1\);
    
    \idle_line_cntr[0]\ : SLE
      port map(D => \idle_line_cntr_s[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[0]_net_1\);
    
    \idle_line_cntr_RNI012B6[5]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[5]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[4]\, S => \idle_line_cntr_s[5]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[5]\);
    
    \idle_line_cntr[12]\ : SLE
      port map(D => \idle_line_cntr_s[12]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[12]_net_1\);
    
    \idle_line_cntr[3]\ : SLE
      port map(D => \idle_line_cntr_s[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[3]_net_1\);
    
    \idle_line_cntr[5]\ : SLE
      port map(D => \idle_line_cntr_s[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[5]_net_1\);
    
    \idle_line_cntr_RNIH8SRA[9]\ : ARI1
      generic map(INIT => x"4D800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[9]_net_1\, D => N_149_i, FCI => 
        \idle_line_cntr_cry[8]\, S => \idle_line_cntr_s[9]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[9]\);
    
    \idle_line_cntr_RNIBNA58[7]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[7]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[6]\, S => \idle_line_cntr_s[7]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[7]\);
    
    \idle_line_cntr[2]\ : SLE
      port map(D => \idle_line_cntr_s[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \idle_line_cntr[2]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity ManchesDecoder_Adapter is

    port( RX_FIFO_DIN         : out   std_logic_vector(7 downto 0);
          manches_in_dly      : out   std_logic_vector(1 downto 0);
          idle_line5          : in    std_logic;
          un2_apb3_reset      : in    std_logic;
          internal_loopback   : in    std_logic;
          MANCHESTER_IN_c     : in    std_logic;
          MANCH_OUT_P_c       : in    std_logic;
          rx_packet_end_all   : in    std_logic;
          idle_line           : out   std_logic;
          irx_center_sample   : out   std_logic;
          sampler_clk1x_en    : out   std_logic;
          clk1x_enable        : in    std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          un2_apb3_reset_i    : in    std_logic
        );

end ManchesDecoder_Adapter;

architecture DEF_ARCH of ManchesDecoder_Adapter is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component IdleLineDetector_1
    port( idle_line5          : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          un2_apb3_reset_i    : in    std_logic := 'U';
          idle_line           : out   std_logic
        );
  end component;

    signal \clock_adjust\, clock_adjust_i, \manches_in_dly[0]\, 
        GND_net_1, \un1_manches_in[0]_net_1\, VCC_net_1, 
        \manches_in_dly[1]\, \decoder_Transition_d[0]_net_1\, 
        un2_rst_i, \decoder_Transition\, 
        \decoder_Transition_d[1]_net_1\, 
        \decoder_Transition_d[2]_net_1\, \RX_FIFO_DIN[0]\, 
        \iNRZ_data\, \sampler_clk1x_en\, \RX_FIFO_DIN[1]\, 
        \RX_FIFO_DIN[2]\, \RX_FIFO_DIN[3]\, \RX_FIFO_DIN[4]\, 
        \RX_FIFO_DIN[5]\, \RX_FIFO_DIN[6]\, 
        \decoder_ShiftReg[0]_net_1\, \clkdiv[3]_net_1\, 
        \manches_ShiftReg[0]_net_1\, un18_rst_i, iNRZ_data_1, 
        irx_center_sample_net_1, isampler_clk1x_en_1, 
        decoder_Transition_1, \manches_Transition\, 
        manches_Transition_1, un16_irx_center_sample, 
        un16_clk1x_enable, \clkdiv[0]_net_1\, \clkdiv_3[0]_net_1\, 
        \clkdiv[1]_net_1\, \clkdiv_3[1]_net_1\, \clkdiv[2]_net_1\, 
        \clkdiv_3[2]_net_1\, \clkdiv_3[3]_net_1\, \idle_line\, 
        \un1_iidle_line\, CO1 : std_logic;

    for all : IdleLineDetector_1
	Use entity work.IdleLineDetector_1(DEF_ARCH);
begin 

    RX_FIFO_DIN(6) <= \RX_FIFO_DIN[6]\;
    RX_FIFO_DIN(5) <= \RX_FIFO_DIN[5]\;
    RX_FIFO_DIN(4) <= \RX_FIFO_DIN[4]\;
    RX_FIFO_DIN(3) <= \RX_FIFO_DIN[3]\;
    RX_FIFO_DIN(2) <= \RX_FIFO_DIN[2]\;
    RX_FIFO_DIN(1) <= \RX_FIFO_DIN[1]\;
    RX_FIFO_DIN(0) <= \RX_FIFO_DIN[0]\;
    manches_in_dly(1) <= \manches_in_dly[1]\;
    manches_in_dly(0) <= \manches_in_dly[0]\;
    idle_line <= \idle_line\;
    irx_center_sample <= irx_center_sample_net_1;
    sampler_clk1x_en <= \sampler_clk1x_en\;

    \s2p_data[2]\ : SLE
      port map(D => \RX_FIFO_DIN[1]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => \sampler_clk1x_en\, ALn => un2_apb3_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN[2]\);
    
    \imanches_in_dly[0]\ : SLE
      port map(D => \un1_manches_in[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \manches_in_dly[0]\);
    
    \decoder_Transition_d[2]\ : SLE
      port map(D => \decoder_Transition_d[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clk1x_enable, ALn => un2_rst_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \decoder_Transition_d[2]_net_1\);
    
    \NRZ_DATA_PROC.un18_rst\ : CFG2
      generic map(INIT => x"1")

      port map(A => \idle_line\, B => un2_apb3_reset, Y => 
        un18_rst_i);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \s2p_data[4]\ : SLE
      port map(D => \RX_FIFO_DIN[3]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => \sampler_clk1x_en\, ALn => un2_apb3_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN[4]\);
    
    clock_adjust_RNIMA1A : CFG1
      generic map(INIT => "01")

      port map(A => \clock_adjust\, Y => clock_adjust_i);
    
    \TRANISTION_DETECT_SHIFTREG_PROC.un2_rst\ : CFG2
      generic map(INIT => x"1")

      port map(A => rx_packet_end_all, B => un2_apb3_reset, Y => 
        un2_rst_i);
    
    \irx_center_sample\ : SLE
      port map(D => un16_irx_center_sample, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clock_adjust_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        irx_center_sample_net_1);
    
    \clkdiv_3[2]\ : CFG3
      generic map(INIT => x"06")

      port map(A => CO1, B => \clkdiv[2]_net_1\, C => 
        \un1_iidle_line\, Y => \clkdiv_3[2]_net_1\);
    
    \s2p_data[1]\ : SLE
      port map(D => \RX_FIFO_DIN[0]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => \sampler_clk1x_en\, ALn => un2_apb3_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN[1]\);
    
    \decoder_ShiftReg[0]\ : SLE
      port map(D => \clkdiv[3]_net_1\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => clk1x_enable, ALn => un2_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \decoder_ShiftReg[0]_net_1\);
    
    \clkdiv_3[1]\ : CFG4
      generic map(INIT => x"006A")

      port map(A => \clkdiv[1]_net_1\, B => \clkdiv[0]_net_1\, C
         => clk1x_enable, D => \un1_iidle_line\, Y => 
        \clkdiv_3[1]_net_1\);
    
    \manches_ShiftReg[0]\ : SLE
      port map(D => \manches_in_dly[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clk1x_enable, ALn => un2_rst_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \manches_ShiftReg[0]_net_1\);
    
    iNRZ_data : SLE
      port map(D => iNRZ_data_1, CLK => CommsFPGA_CCC_0_GL0, EN
         => irx_center_sample_net_1, ALn => un18_rst_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \iNRZ_data\);
    
    \clkdiv[2]\ : SLE
      port map(D => \clkdiv_3[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clock_adjust_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \clkdiv[2]_net_1\);
    
    \s2p_data[3]\ : SLE
      port map(D => \RX_FIFO_DIN[2]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => \sampler_clk1x_en\, ALn => un2_apb3_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN[3]\);
    
    \decoder_Transition_d[0]\ : SLE
      port map(D => \decoder_Transition\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clk1x_enable, ALn => un2_rst_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \decoder_Transition_d[0]_net_1\);
    
    decoder_Transition : SLE
      port map(D => decoder_Transition_1, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clk1x_enable, ALn => un2_rst_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \decoder_Transition\);
    
    \clkdiv_3[3]\ : CFG4
      generic map(INIT => x"FF6A")

      port map(A => \clkdiv[3]_net_1\, B => \clkdiv[2]_net_1\, C
         => CO1, D => \un1_iidle_line\, Y => \clkdiv_3[3]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \clkdiv[1]\ : SLE
      port map(D => \clkdiv_3[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clock_adjust_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \clkdiv[1]_net_1\);
    
    \s2p_data[5]\ : SLE
      port map(D => \RX_FIFO_DIN[4]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => \sampler_clk1x_en\, ALn => un2_apb3_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN[5]\);
    
    RX_IDLE_LINE_DETECTOR : IdleLineDetector_1
      port map(idle_line5 => idle_line5, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, un2_apb3_reset_i => un2_apb3_reset_i, 
        idle_line => \idle_line\);
    
    un10_clk1x_enable : CFG2
      generic map(INIT => x"6")

      port map(A => \clkdiv[3]_net_1\, B => 
        \decoder_ShiftReg[0]_net_1\, Y => decoder_Transition_1);
    
    \RX_CENTER_SAMPLE_PROC.un16_irx_center_sample_0_a2\ : CFG3
      generic map(INIT => x"40")

      port map(A => \clkdiv[2]_net_1\, B => \clkdiv[1]_net_1\, C
         => \clkdiv[0]_net_1\, Y => un16_irx_center_sample);
    
    clock_adjust : SLE
      port map(D => un16_clk1x_enable, CLK => CommsFPGA_CCC_0_GL0, 
        EN => clk1x_enable, ALn => un2_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \clock_adjust\);
    
    \un1_manches_in[0]\ : CFG3
      generic map(INIT => x"A3")

      port map(A => MANCH_OUT_P_c, B => MANCHESTER_IN_c, C => 
        internal_loopback, Y => \un1_manches_in[0]_net_1\);
    
    \SAMPLE_CLK1X_EN_PROC.isampler_clk1x_en_1_0_a2\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \clkdiv[0]_net_1\, B => \clkdiv[3]_net_1\, C
         => \clkdiv[2]_net_1\, D => \clkdiv[1]_net_1\, Y => 
        isampler_clk1x_en_1);
    
    manches_Transition : SLE
      port map(D => manches_Transition_1, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clk1x_enable, ALn => un2_rst_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \manches_Transition\);
    
    \CLOCK_ADJUST_PROC.un16_clk1x_enable\ : CFG2
      generic map(INIT => x"8")

      port map(A => \decoder_Transition_d[2]_net_1\, B => 
        \manches_Transition\, Y => un16_clk1x_enable);
    
    \s2p_data[7]\ : SLE
      port map(D => \RX_FIFO_DIN[6]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => \sampler_clk1x_en\, ALn => un2_apb3_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RX_FIFO_DIN(7));
    
    \clkdiv[0]\ : SLE
      port map(D => \clkdiv_3[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clock_adjust_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \clkdiv[0]_net_1\);
    
    \clkdiv[3]\ : SLE
      port map(D => \clkdiv_3[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clock_adjust_i, ALn => 
        un2_apb3_reset_i, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \clkdiv[3]_net_1\);
    
    un1_iidle_line : CFG2
      generic map(INIT => x"E")

      port map(A => \idle_line\, B => rx_packet_end_all, Y => 
        \un1_iidle_line\);
    
    \clkdiv_3[0]\ : CFG3
      generic map(INIT => x"14")

      port map(A => \un1_iidle_line\, B => \clkdiv[0]_net_1\, C
         => clk1x_enable, Y => \clkdiv_3[0]_net_1\);
    
    \imanches_in_dly[1]\ : SLE
      port map(D => \manches_in_dly[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \manches_in_dly[1]\);
    
    \un1_clkdiv_1.CO1\ : CFG3
      generic map(INIT => x"80")

      port map(A => \clkdiv[0]_net_1\, B => clk1x_enable, C => 
        \clkdiv[1]_net_1\, Y => CO1);
    
    \decoder_Transition_d[1]\ : SLE
      port map(D => \decoder_Transition_d[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clk1x_enable, ALn => un2_rst_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \decoder_Transition_d[1]_net_1\);
    
    \s2p_data[0]\ : SLE
      port map(D => \iNRZ_data\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \sampler_clk1x_en\, ALn => un2_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN[0]\);
    
    \NRZ_DATA_PROC.iNRZ_data_1\ : CFG2
      generic map(INIT => x"6")

      port map(A => \clkdiv[3]_net_1\, B => \manches_in_dly[1]\, 
        Y => iNRZ_data_1);
    
    \s2p_data[6]\ : SLE
      port map(D => \RX_FIFO_DIN[5]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => \sampler_clk1x_en\, ALn => un2_apb3_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN[6]\);
    
    un4_clk1x_enable : CFG2
      generic map(INIT => x"6")

      port map(A => \manches_in_dly[1]\, B => 
        \manches_ShiftReg[0]_net_1\, Y => manches_Transition_1);
    
    isampler_clk1x_en : SLE
      port map(D => isampler_clk1x_en_1, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clock_adjust_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sampler_clk1x_en\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CRC16_Generator_1 is

    port( RX_FIFO_DIN         : in    std_logic_vector(7 downto 0);
          rx_crc_data_calc    : out   std_logic_vector(15 downto 0);
          lfsr_c_i_i_0        : in    std_logic;
          rx_crc_gen          : in    std_logic;
          sampler_clk1x_en    : in    std_logic;
          iRX_FIFO_wr_en      : in    std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          rx_crc_reset_i      : in    std_logic
        );

end CRC16_Generator_1;

architecture DEF_ARCH of CRC16_Generator_1 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \rx_crc_data_calc[13]\, GND_net_1, 
        \rx_crc_data_calc[5]\, \N_46_i\, VCC_net_1, 
        \rx_crc_data_calc[14]\, \rx_crc_data_calc[6]\, 
        \rx_crc_data_calc[15]\, \lfsr_c[15]\, 
        \rx_crc_data_calc[0]\, \lfsr_c[0]\, \rx_crc_data_calc[1]\, 
        \lfsr_c[1]\, \rx_crc_data_calc[2]\, N_79_i, 
        \rx_crc_data_calc[3]\, \lfsr_c[3]\, \rx_crc_data_calc[4]\, 
        \lfsr_c[5]\, \lfsr_c[6]\, \rx_crc_data_calc[7]\, 
        \lfsr_c[7]\, \rx_crc_data_calc[8]\, N_133_i_i, 
        \rx_crc_data_calc[9]\, N_132_i_i, \rx_crc_data_calc[10]\, 
        \rx_crc_data_calc[11]\, \rx_crc_data_calc[12]\, N_116_i
         : std_logic;

begin 

    rx_crc_data_calc(15) <= \rx_crc_data_calc[15]\;
    rx_crc_data_calc(14) <= \rx_crc_data_calc[14]\;
    rx_crc_data_calc(13) <= \rx_crc_data_calc[13]\;
    rx_crc_data_calc(12) <= \rx_crc_data_calc[12]\;
    rx_crc_data_calc(11) <= \rx_crc_data_calc[11]\;
    rx_crc_data_calc(10) <= \rx_crc_data_calc[10]\;
    rx_crc_data_calc(9) <= \rx_crc_data_calc[9]\;
    rx_crc_data_calc(8) <= \rx_crc_data_calc[8]\;
    rx_crc_data_calc(7) <= \rx_crc_data_calc[7]\;
    rx_crc_data_calc(6) <= \rx_crc_data_calc[6]\;
    rx_crc_data_calc(5) <= \rx_crc_data_calc[5]\;
    rx_crc_data_calc(4) <= \rx_crc_data_calc[4]\;
    rx_crc_data_calc(3) <= \rx_crc_data_calc[3]\;
    rx_crc_data_calc(2) <= \rx_crc_data_calc[2]\;
    rx_crc_data_calc(1) <= \rx_crc_data_calc[1]\;
    rx_crc_data_calc(0) <= \rx_crc_data_calc[0]\;

    \lfsr_q[9]\ : SLE
      port map(D => N_132_i_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \N_46_i\, ALn => rx_crc_reset_i, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_calc[9]\);
    
    \lfsr_q[6]\ : SLE
      port map(D => \lfsr_c[6]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \N_46_i\, ALn => rx_crc_reset_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rx_crc_data_calc[6]\);
    
    \lfsr_q[3]\ : SLE
      port map(D => \lfsr_c[3]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \N_46_i\, ALn => rx_crc_reset_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rx_crc_data_calc[3]\);
    
    \lfsr_q[10]\ : SLE
      port map(D => \rx_crc_data_calc[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \N_46_i\, ALn => 
        rx_crc_reset_i, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_calc[10]\);
    
    \lfsr_q[2]\ : SLE
      port map(D => N_79_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \N_46_i\, ALn => rx_crc_reset_i, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_calc[2]\);
    
    \lfsr_c_0_a2[5]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \rx_crc_data_calc[12]\, B => 
        \rx_crc_data_calc[11]\, C => RX_FIFO_DIN(4), D => 
        RX_FIFO_DIN(3), Y => \lfsr_c[5]\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \lfsr_q[1]\ : SLE
      port map(D => \lfsr_c[1]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \N_46_i\, ALn => rx_crc_reset_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rx_crc_data_calc[1]\);
    
    \lfsr_q[7]\ : SLE
      port map(D => \lfsr_c[7]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \N_46_i\, ALn => rx_crc_reset_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rx_crc_data_calc[7]\);
    
    \lfsr_c_0_a2[3]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \rx_crc_data_calc[9]\, B => 
        \rx_crc_data_calc[10]\, C => RX_FIFO_DIN(2), D => 
        RX_FIFO_DIN(1), Y => \lfsr_c[3]\);
    
    \lfsr_q[4]\ : SLE
      port map(D => lfsr_c_i_i_0, CLK => CommsFPGA_CCC_0_GL0, EN
         => \N_46_i\, ALn => rx_crc_reset_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rx_crc_data_calc[4]\);
    
    \lfsr_q[11]\ : SLE
      port map(D => \rx_crc_data_calc[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \N_46_i\, ALn => 
        rx_crc_reset_i, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_calc[11]\);
    
    \lfsr_q[5]\ : SLE
      port map(D => \lfsr_c[5]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \N_46_i\, ALn => rx_crc_reset_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rx_crc_data_calc[5]\);
    
    \lfsr_c_0_a2[1]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => N_116_i, B => \lfsr_c[7]\, C => \lfsr_c[5]\, 
        D => \lfsr_c[3]\, Y => \lfsr_c[1]\);
    
    \lfsr_q_RNO[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => N_116_i, B => \rx_crc_data_calc[1]\, Y => 
        N_132_i_i);
    
    \lfsr_q[0]\ : SLE
      port map(D => \lfsr_c[0]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \N_46_i\, ALn => rx_crc_reset_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rx_crc_data_calc[0]\);
    
    \lfsr_c_0_a2[7]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \rx_crc_data_calc[13]\, B => 
        \rx_crc_data_calc[14]\, C => RX_FIFO_DIN(6), D => 
        RX_FIFO_DIN(5), Y => \lfsr_c[7]\);
    
    \lfsr_c_0_a2[15]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \lfsr_c[0]\, B => \rx_crc_data_calc[7]\, Y
         => \lfsr_c[15]\);
    
    \lfsr_q[12]\ : SLE
      port map(D => \rx_crc_data_calc[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \N_46_i\, ALn => 
        rx_crc_reset_i, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_calc[12]\);
    
    \lfsr_c_0_a2_2_x4[2]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \rx_crc_data_calc[8]\, B => 
        \rx_crc_data_calc[9]\, C => RX_FIFO_DIN(1), D => 
        RX_FIFO_DIN(0), Y => N_79_i);
    
    \lfsr_q[14]\ : SLE
      port map(D => \rx_crc_data_calc[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \N_46_i\, ALn => 
        rx_crc_reset_i, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_calc[14]\);
    
    \lfsr_c_0_a2_i_x2[8]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => RX_FIFO_DIN(6), B => N_116_i, C => 
        \rx_crc_data_calc[0]\, D => \rx_crc_data_calc[14]\, Y => 
        N_133_i_i);
    
    \lfsr_c_0_a2[6]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \rx_crc_data_calc[13]\, B => 
        \rx_crc_data_calc[12]\, C => RX_FIFO_DIN(5), D => 
        RX_FIFO_DIN(4), Y => \lfsr_c[6]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \lfsr_c_0_a2_1_0_x2[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => RX_FIFO_DIN(7), B => \rx_crc_data_calc[15]\, 
        Y => N_116_i);
    
    \lfsr_q[8]\ : SLE
      port map(D => N_133_i_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \N_46_i\, ALn => rx_crc_reset_i, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_calc[8]\);
    
    \lfsr_q[13]\ : SLE
      port map(D => \rx_crc_data_calc[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \N_46_i\, ALn => 
        rx_crc_reset_i, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_calc[13]\);
    
    \lfsr_c_0_a2[0]\ : CFG3
      generic map(INIT => x"96")

      port map(A => \lfsr_c[1]\, B => \rx_crc_data_calc[8]\, C
         => RX_FIFO_DIN(0), Y => \lfsr_c[0]\);
    
    N_46_i : CFG3
      generic map(INIT => x"80")

      port map(A => iRX_FIFO_wr_en, B => sampler_clk1x_en, C => 
        rx_crc_gen, Y => \N_46_i\);
    
    \lfsr_q[15]\ : SLE
      port map(D => \lfsr_c[15]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \N_46_i\, ALn => rx_crc_reset_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rx_crc_data_calc[15]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity ReadFIFO_Write_SM is

    port( consumer_type2_reg  : in    std_logic_vector(9 downto 0);
          consumer_type4_reg  : in    std_logic_vector(9 downto 0);
          consumer_type3_reg  : in    std_logic_vector(9 downto 0);
          consumer_type1_reg  : in    std_logic_vector(9 downto 0);
          rx_crc_data_calc    : out   std_logic_vector(11 downto 10);
          RX_FIFO_DIN         : in    std_logic_vector(7 downto 0);
          RX_FIFO_DIN_pipe    : out   std_logic_vector(8 downto 0);
          lfsr_c_i_i_0        : in    std_logic;
          DRVR_EN_c           : in    std_logic;
          clk1x_enable        : in    std_logic;
          un2_apb3_reset      : in    std_logic;
          tx_col_detect_en    : in    std_logic;
          packet_avail        : in    std_logic;
          sampler_clk1x_en    : in    std_logic;
          idle_line           : in    std_logic;
          RX_InProcess_d1     : out   std_logic;
          rx_packet_complt    : out   std_logic;
          N_535               : out   std_logic;
          RX_EarlyTerm        : out   std_logic;
          SM_advance_i        : out   std_logic;
          rx_crc_HighByte_en  : out   std_logic;
          iRX_FIFO_wr_en      : out   std_logic;
          N_41_i              : in    std_logic;
          N_993_i             : in    std_logic;
          un2_apb3_reset_i    : in    std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          rx_CRC_error_i      : out   std_logic;
          rx_CRC_error        : out   std_logic
        );

end ReadFIFO_Write_SM;

architecture DEF_ARCH of ReadFIFO_Write_SM is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CRC16_Generator_1
    port( RX_FIFO_DIN         : in    std_logic_vector(7 downto 0) := (others => 'U');
          rx_crc_data_calc    : out   std_logic_vector(15 downto 0);
          lfsr_c_i_i_0        : in    std_logic := 'U';
          rx_crc_gen          : in    std_logic := 'U';
          sampler_clk1x_en    : in    std_logic := 'U';
          iRX_FIFO_wr_en      : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          rx_crc_reset_i      : in    std_logic := 'U'
        );
  end component;

    signal rx_crc_reset_i, \rx_crc_reset\, 
        \un65_sm_advance_i_cry_9\, \un65_sm_advance_i_i[1]\, 
        un9_rst, un9_rst_i, rx_CRC_error_net_1, 
        \bit_cntr[2]_net_1\, VCC_net_1, un16_rst_i, N_151_i_i, 
        GND_net_1, \SM_advancebit_cntr[0]_net_1\, N_174_i_i, 
        \SM_advancebit_cntr[1]_net_1\, N_338_i, 
        \SM_advancebit_cntr[2]_net_1\, N_150_i_i, 
        \un56_sm_advance_i[4]\, \un56_sm_advance_i_i[4]\, 
        un1_ReadFIFO_WR_STATE_14, \un56_sm_advance_i[3]\, 
        \un56_sm_advance_i_i[3]\, \un56_sm_advance_i[2]\, 
        \un56_sm_advance_i_i[2]\, \un56_sm_advance_i[1]\, 
        \un56_sm_advance_i_i[1]\, \un65_sm_advance_i[9]\, 
        \un65_sm_advance_i_i[9]\, \un65_sm_advance_i[8]\, 
        \un65_sm_advance_i_i[8]\, \un65_sm_advance_i[7]\, 
        \un65_sm_advance_i_i[7]\, \un65_sm_advance_i[6]\, 
        \un65_sm_advance_i_i[6]\, \un65_sm_advance_i[5]\, 
        \un65_sm_advance_i_i[5]\, \un65_sm_advance_i[4]\, 
        \un65_sm_advance_i_i[4]\, \un65_sm_advance_i[3]\, 
        \un65_sm_advance_i_i[3]\, \un65_sm_advance_i[2]\, 
        \un65_sm_advance_i_i[2]\, \un65_sm_advance_i[1]\, 
        \bit_cntr[0]_net_1\, N_1082_i, \bit_cntr[1]_net_1\, 
        N_337_i, \rx_crc_data_store[8]_net_1\, 
        \RX_FIFO_DIN_pipe[0]\, \rx_crc_data_store[9]_net_1\, 
        \RX_FIFO_DIN_pipe[1]\, \rx_crc_data_store[10]_net_1\, 
        \RX_FIFO_DIN_pipe[2]\, \rx_crc_data_store[11]_net_1\, 
        \RX_FIFO_DIN_pipe[3]\, \rx_crc_data_store[12]_net_1\, 
        \RX_FIFO_DIN_pipe[4]\, \rx_crc_data_store[13]_net_1\, 
        \RX_FIFO_DIN_pipe[5]\, \rx_crc_data_store[14]_net_1\, 
        \RX_FIFO_DIN_pipe[6]\, \rx_crc_data_store[15]_net_1\, 
        \RX_FIFO_DIN_pipe[7]\, \un56_sm_advance_i[11]\, 
        un65_sm_advance_i_cry_0_Y, \un56_sm_advance_i[10]\, 
        \un56_sm_advance_i_i[10]\, \un56_sm_advance_i[9]\, 
        \un56_sm_advance_i_i[9]\, \un56_sm_advance_i[8]\, 
        \un56_sm_advance_i_i[8]\, \un56_sm_advance_i[7]\, 
        \un56_sm_advance_i_i[7]\, \un56_sm_advance_i[6]\, 
        \un56_sm_advance_i_i[6]\, \un56_sm_advance_i[5]\, 
        \un56_sm_advance_i_i[5]\, \rx_packet_length[4]_net_1\, 
        N_43_i, \rx_packet_length[5]_net_1\, 
        un56_sm_advance_i_axb_4_i, \rx_packet_length[6]_net_1\, 
        un56_sm_advance_i_axb_5_i, \rx_packet_length[7]_net_1\, 
        un56_sm_advance_i_axb_6_i, \rx_packet_length[8]_net_1\, 
        un56_sm_advance_i_axb_7_i, \rx_packet_length[9]_net_1\, 
        un56_sm_advance_i_axb_8_i, \rx_packet_length[10]_net_1\, 
        un56_sm_advance_i_axb_9_i, \rx_crc_data_store[0]_net_1\, 
        \un1_rx_fifo_din_d3[0]_net_1\, 
        \rx_crc_data_store[1]_net_1\, 
        \un1_rx_fifo_din_d3[1]_net_1\, 
        \rx_crc_data_store[2]_net_1\, 
        \un1_rx_fifo_din_d3[2]_net_1\, 
        \rx_crc_data_store[3]_net_1\, 
        \un1_rx_fifo_din_d3[3]_net_1\, 
        \rx_crc_data_store[4]_net_1\, 
        \un1_rx_fifo_din_d3[4]_net_1\, 
        \rx_crc_data_store[5]_net_1\, 
        \un1_rx_fifo_din_d3[5]_net_1\, 
        \rx_crc_data_store[6]_net_1\, 
        \un1_rx_fifo_din_d3[6]_net_1\, 
        \rx_crc_data_store[7]_net_1\, 
        \un1_rx_fifo_din_d3[7]_net_1\, \consumer_type[0]_net_1\, 
        N_313, \un1_ReadFIFO_WR_STATE_12_0_i_i_a3_0\, 
        \consumer_type[1]_net_1\, N_1356, 
        \consumer_type[2]_net_1\, N_66_i, 
        \consumer_type[3]_net_1\, N_819_i, 
        \consumer_type[4]_net_1\, N_820_i, 
        \consumer_type[5]_net_1\, N_72_i, 
        \consumer_type[6]_net_1\, N_74_i, 
        \consumer_type[7]_net_1\, N_812_i, 
        \consumer_type[8]_net_1\, N_813_i, 
        \consumer_type[9]_net_1\, N_815_i, 
        \rx_packet_length[0]_net_1\, N_348_i, 
        \rx_packet_length[1]_net_1\, un56_sm_advance_i_axb_0_i, 
        \rx_packet_length[2]_net_1\, un56_sm_advance_i_axb_1_i, 
        \rx_packet_length[3]_net_1\, un56_sm_advance_i_axb_2_i, 
        iRX_FIFO_wr_en_net_1, un5_packet_avail, N_996_i, 
        \irx_packet_end\, N_669_i, 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0_0\, 
        \ReadFIFO_WR_STATE[3]_net_1\, rx_crc_HighByte_en_net_1, 
        N_399, \rx_crc_gen\, un1_ReadFIFO_WR_STATE_15, 
        SM_advance_i_net_1, un2_packet_avail, \rx_end_rst\, 
        N_259_i, \RX_EarlyTerm\, \ReadFIFO_WR_STATE[4]_net_1\, 
        N_21, N_20, \N_535\, N_18, N_17, N_15, N_14, N_12, N_11, 
        N_9, N_8, N_6, N_5, N_3, N_2, N_24, 
        \un65_sm_advance_i[10]\, \un65_sm_advance_i_i[10]\, N_87, 
        \rx_packet_complt_1_sqmuxa\, \RX_InProcess\, N_250_i, 
        N_23, \ReadFIFO_WR_STATE[2]_net_1\, 
        \ReadFIFO_WR_STATE[1]_net_1\, 
        \ReadFIFO_WR_STATE_ns[8]_net_1\, 
        \ReadFIFO_WR_STATE[0]_net_1\, \ReadFIFO_WR_STATE_ns[9]\, 
        \ReadFIFO_WR_STATE[9]_net_1\, N_233_i, 
        \ReadFIFO_WR_STATE[8]_net_1\, N_321, 
        \ReadFIFO_WR_STATE[7]_net_1\, \ReadFIFO_WR_STATE_202\, 
        \ReadFIFO_WR_STATE[6]_net_1\, \ReadFIFO_WR_STATE_ns[3]\, 
        \ReadFIFO_WR_STATE[5]_net_1\, \ReadFIFO_WR_STATE_ns[4]\, 
        \ReadFIFO_WR_STATE_ns[5]\, \ReadFIFO_WR_STATE_ns[6]\, 
        \rx_byte_cntr[0]_net_1\, \rx_byte_cntr_lm[0]\, N_992_i, 
        \rx_byte_cntr[1]_net_1\, \rx_byte_cntr_lm[1]\, 
        \rx_byte_cntr[2]_net_1\, \rx_byte_cntr_lm[2]\, 
        \rx_byte_cntr[3]_net_1\, \rx_byte_cntr_lm[3]\, 
        \rx_byte_cntr[4]_net_1\, \rx_byte_cntr_lm[4]\, 
        \rx_byte_cntr[5]_net_1\, \rx_byte_cntr_lm[5]\, 
        \rx_byte_cntr[6]_net_1\, \rx_byte_cntr_lm[6]\, 
        \rx_byte_cntr[7]_net_1\, \rx_byte_cntr_lm[7]\, 
        \rx_byte_cntr[8]_net_1\, \rx_byte_cntr_lm[8]\, 
        \rx_byte_cntr[9]_net_1\, \rx_byte_cntr_lm[9]\, 
        \rx_byte_cntr[10]_net_1\, \rx_byte_cntr_lm[10]\, 
        \rx_byte_cntr[11]_net_1\, \rx_byte_cntr_lm[11]\, 
        \un56_sm_advance_i_cry_0\, N_1475, N_539, 
        \un56_sm_advance_i_cry_1\, \un56_sm_advance_i_cry_2\, 
        \un56_sm_advance_i_cry_3\, \un56_sm_advance_i_cry_4\, 
        \un56_sm_advance_i_cry_5\, \un56_sm_advance_i_cry_6\, 
        \un56_sm_advance_i_cry_7\, N_572, 
        \un56_sm_advance_i_cry_8\, \un65_sm_advance_i_cry_0\, 
        \un65_sm_advance_i_cry_1\, \un65_sm_advance_i_cry_2\, 
        \un65_sm_advance_i_cry_3\, \un65_sm_advance_i_cry_4\, 
        \un65_sm_advance_i_cry_5\, \un65_sm_advance_i_cry_6\, 
        \un65_sm_advance_i_cry_7\, \un65_sm_advance_i_cry_8\, 
        un67_sm_advance_i_cry_0, un67_sm_advance_i_cry_1, 
        un67_sm_advance_i_cry_2, un67_sm_advance_i_cry_3, 
        un67_sm_advance_i_cry_4, un67_sm_advance_i_cry_5, 
        un67_sm_advance_i_cry_6, un67_sm_advance_i_cry_7, 
        un67_sm_advance_i_cry_8, un67_sm_advance_i_cry_9, 
        un67_sm_advance_i_cry_10, un67_sm_advance_i, 
        \un58_sm_advance_i_0_data_tmp[0]\, 
        \un58_sm_advance_i_0_data_tmp[1]\, 
        \un58_sm_advance_i_0_data_tmp[2]\, 
        \un58_sm_advance_i_0_data_tmp[3]\, 
        \un58_sm_advance_i_0_data_tmp[4]\, 
        \un58_sm_advance_i_0_data_tmp[5]\, 
        \un1_sampler_clk1x_en_0_data_tmp[0]\, 
        \rx_crc_data_calc[0]\, \rx_crc_data_calc[1]\, 
        \un1_sampler_clk1x_en_0_data_tmp[1]\, 
        \rx_crc_data_calc[2]\, \rx_crc_data_calc[3]\, 
        \un1_sampler_clk1x_en_0_data_tmp[2]\, 
        \rx_crc_data_calc[4]\, \rx_crc_data_calc[5]\, 
        \un1_sampler_clk1x_en_0_data_tmp[3]\, 
        \rx_crc_data_calc[6]\, \rx_crc_data_calc[7]\, 
        \un1_sampler_clk1x_en_0_data_tmp[4]\, 
        \rx_crc_data_calc[8]\, \rx_crc_data_calc[9]\, 
        \un1_sampler_clk1x_en_0_data_tmp[5]\, 
        \rx_crc_data_calc[10]\, \rx_crc_data_calc[11]\, 
        \un1_sampler_clk1x_en_0_data_tmp[6]\, 
        \rx_crc_data_calc[12]\, \rx_crc_data_calc[13]\, 
        \un1_sampler_clk1x_en_0_data_tmp[7]\, 
        \rx_crc_data_calc[14]\, \rx_crc_data_calc[15]\, 
        rx_byte_cntr_s_391_FCO, \rx_byte_cntr_cry[1]_net_1\, 
        \rx_byte_cntr_s[1]\, \rx_byte_cntr_cry[2]_net_1\, 
        \rx_byte_cntr_s[2]\, \rx_byte_cntr_cry[3]_net_1\, 
        \rx_byte_cntr_s[3]\, \rx_byte_cntr_cry[4]_net_1\, 
        \rx_byte_cntr_s[4]\, \rx_byte_cntr_cry[5]_net_1\, 
        \rx_byte_cntr_s[5]\, \rx_byte_cntr_cry[6]_net_1\, 
        \rx_byte_cntr_s[6]\, \rx_byte_cntr_cry[7]_net_1\, 
        \rx_byte_cntr_s[7]\, \rx_byte_cntr_cry[8]_net_1\, 
        \rx_byte_cntr_s[8]\, \rx_byte_cntr_cry[9]_net_1\, 
        \rx_byte_cntr_s[9]\, \rx_byte_cntr_s[11]_net_1\, 
        \rx_byte_cntr_cry[10]_net_1\, \rx_byte_cntr_s[10]\, 
        un56_sm_advance_i_s_9_395_FCO, un56_sm_advance_i_s_9_sf, 
        N_992_i_1, N_1358, N_1469, 
        \ReadFIFO_WR_STATE_ns_0_0_a2_0_0[9]_net_1\, 
        un32_sm_advance_i_7, un38_sm_advance_i_7, N_1328, 
        consumer_type_0_sqmuxa, N_1467, un38_sm_advance_i_NE_4, 
        un38_sm_advance_i_NE_3, un38_sm_advance_i_NE_1, 
        un38_sm_advance_i_NE_0, un29_sm_advance_i_NE_4, 
        un29_sm_advance_i_NE_3, un29_sm_advance_i_NE_2, 
        un29_sm_advance_i_NE_1, un29_sm_advance_i_NE_0, 
        un32_sm_advance_i_NE_4, un32_sm_advance_i_NE_3, 
        un32_sm_advance_i_NE_1, un32_sm_advance_i_NE_0, 
        un35_sm_advance_i_NE_4, un35_sm_advance_i_NE_3, 
        un35_sm_advance_i_NE_2, un35_sm_advance_i_NE_1, 
        un35_sm_advance_i_NE_0, N_1036, N_1292, 
        \ReadFIFO_WR_STATE_ns_0_0_0[5]_net_1\, 
        un38_sm_advance_i_NE_6, un32_sm_advance_i_NE_6, N_1333, 
        un29_sm_advance_i_NE_7, un32_sm_advance_i_NE_7, 
        un35_sm_advance_i_NE_7, N_1382, un39_sm_advance_i, 
        un40_sm_advance_i_1, un40_sm_advance_i_0, 
        un40_sm_advance_i : std_logic;

    for all : CRC16_Generator_1
	Use entity work.CRC16_Generator_1(DEF_ARCH);
begin 

    rx_crc_data_calc(11) <= \rx_crc_data_calc[11]\;
    rx_crc_data_calc(10) <= \rx_crc_data_calc[10]\;
    RX_FIFO_DIN_pipe(7) <= \RX_FIFO_DIN_pipe[7]\;
    RX_FIFO_DIN_pipe(6) <= \RX_FIFO_DIN_pipe[6]\;
    RX_FIFO_DIN_pipe(5) <= \RX_FIFO_DIN_pipe[5]\;
    RX_FIFO_DIN_pipe(4) <= \RX_FIFO_DIN_pipe[4]\;
    RX_FIFO_DIN_pipe(3) <= \RX_FIFO_DIN_pipe[3]\;
    RX_FIFO_DIN_pipe(2) <= \RX_FIFO_DIN_pipe[2]\;
    RX_FIFO_DIN_pipe(1) <= \RX_FIFO_DIN_pipe[1]\;
    RX_FIFO_DIN_pipe(0) <= \RX_FIFO_DIN_pipe[0]\;
    N_535 <= \N_535\;
    RX_EarlyTerm <= \RX_EarlyTerm\;
    SM_advance_i <= SM_advance_i_net_1;
    rx_crc_HighByte_en <= rx_crc_HighByte_en_net_1;
    iRX_FIFO_wr_en <= iRX_FIFO_wr_en_net_1;
    rx_CRC_error <= rx_CRC_error_net_1;

    \consumer_type_RNO[4]\ : CFG4
      generic map(INIT => x"F088")

      port map(A => RX_FIFO_DIN(2), B => consumer_type_0_sqmuxa, 
        C => \consumer_type[4]_net_1\, D => 
        \ReadFIFO_WR_STATE[8]_net_1\, Y => N_820_i);
    
    ReadFIFO_WR_STATE_202 : CFG3
      generic map(INIT => x"CA")

      port map(A => \ReadFIFO_WR_STATE[7]_net_1\, B => 
        \ReadFIFO_WR_STATE[8]_net_1\, C => \N_535\, Y => 
        \ReadFIFO_WR_STATE_202\);
    
    un56_sm_advance_i_cry_8 : ARI1
      generic map(INIT => x"6FF35")

      port map(A => N_1475, B => RX_FIFO_DIN(1), C => 
        \rx_packet_length[9]_net_1\, D => N_572, FCI => 
        \un56_sm_advance_i_cry_7\, S => \un56_sm_advance_i_i[3]\, 
        Y => OPEN, FCO => \un56_sm_advance_i_cry_8\);
    
    \rx_packet_length[5]\ : SLE
      port map(D => un56_sm_advance_i_axb_4_i, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \rx_packet_length[5]_net_1\);
    
    \ReadFIFO_WR_SM.un32_sm_advance_i_NE_7\ : CFG3
      generic map(INIT => x"FE")

      port map(A => un32_sm_advance_i_NE_4, B => 
        un32_sm_advance_i_NE_1, C => un32_sm_advance_i_NE_0, Y
         => un32_sm_advance_i_NE_7);
    
    \ReadFIFO_WR_SM.un35_sm_advance_i_NE_4\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type3_reg(1), B => 
        consumer_type3_reg(0), C => \consumer_type[1]_net_1\, D
         => \consumer_type[0]_net_1\, Y => un35_sm_advance_i_NE_4);
    
    \rx_packet_length_ret[4]\ : SLE
      port map(D => \un56_sm_advance_i_i[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => GND_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \un56_sm_advance_i[7]\);
    
    \ReadFIFO_WR_SM.consumer_type_12_i_i[1]\ : CFG4
      generic map(INIT => x"AA0C")

      port map(A => RX_FIFO_DIN(7), B => \consumer_type[1]_net_1\, 
        C => N_1467, D => N_1292, Y => N_1356);
    
    rx_crc_LowByte_en : SLE
      port map(D => \ReadFIFO_WR_STATE[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0_0\, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => RX_FIFO_DIN_pipe(8));
    
    \ReadFIFO_WR_SM.un58_sm_advance_i_0_I_27\ : ARI1
      generic map(INIT => x"68241")

      port map(A => \un56_sm_advance_i[4]\, B => 
        \rx_byte_cntr[8]_net_1\, C => \rx_byte_cntr[9]_net_1\, D
         => \un56_sm_advance_i[3]\, FCI => 
        \un58_sm_advance_i_0_data_tmp[3]\, S => OPEN, Y => OPEN, 
        FCO => \un58_sm_advance_i_0_data_tmp[4]\);
    
    un56_sm_advance_i_cry_6 : ARI1
      generic map(INIT => x"6FF35")

      port map(A => N_1475, B => RX_FIFO_DIN(7), C => 
        \rx_packet_length[7]_net_1\, D => N_539, FCI => 
        \un56_sm_advance_i_cry_5\, S => \un56_sm_advance_i_i[5]\, 
        Y => OPEN, FCO => \un56_sm_advance_i_cry_6\);
    
    \rx_byte_cntr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rx_byte_cntr[10]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \rx_byte_cntr_cry[9]_net_1\, S => \rx_byte_cntr_s[10]\, Y
         => OPEN, FCO => \rx_byte_cntr_cry[10]_net_1\);
    
    \rx_packet_length_ret[0]\ : SLE
      port map(D => un65_sm_advance_i_cry_0_Y, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => GND_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \un56_sm_advance_i[11]\);
    
    \rx_byte_cntr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rx_byte_cntr[9]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \rx_byte_cntr_cry[8]_net_1\, S => \rx_byte_cntr_s[9]\, Y
         => OPEN, FCO => \rx_byte_cntr_cry[9]_net_1\);
    
    un1_ReadFIFO_WR_STATE_12_0_i_i_a3_0_o2 : CFG3
      generic map(INIT => x"DF")

      port map(A => sampler_clk1x_en, B => 
        \ReadFIFO_WR_STATE[6]_net_1\, C => SM_advance_i_net_1, Y
         => N_572);
    
    \SM_advancebit_cntr_RNO[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => N_996_i, B => \SM_advancebit_cntr[0]_net_1\, 
        Y => N_174_i_i);
    
    \rx_packet_length[10]\ : SLE
      port map(D => un56_sm_advance_i_axb_9_i, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \rx_packet_length[10]_net_1\);
    
    un1_iRX_EarlyTerm_1_sqmuxa_1_0_0 : CFG4
      generic map(INIT => x"CECC")

      port map(A => N_1333, B => \N_535\, C => 
        \ReadFIFO_WR_STATE[8]_net_1\, D => N_1475, Y => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0_0\);
    
    \rx_byte_cntr[11]\ : SLE
      port map(D => \rx_byte_cntr_lm[11]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_992_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_byte_cntr[11]_net_1\);
    
    \ReadFIFO_WR_SM.un58_sm_advance_i_0_I_33\ : ARI1
      generic map(INIT => x"68241")

      port map(A => \un56_sm_advance_i[8]\, B => 
        \rx_byte_cntr[4]_net_1\, C => \rx_byte_cntr[5]_net_1\, D
         => \un56_sm_advance_i[7]\, FCI => 
        \un58_sm_advance_i_0_data_tmp[1]\, S => OPEN, Y => OPEN, 
        FCO => \un58_sm_advance_i_0_data_tmp[2]\);
    
    ReadFIFO_WR_STATE_1_sqmuxa_1_i_i_a3_0_a2 : CFG2
      generic map(INIT => x"4")

      port map(A => \un58_sm_advance_i_0_data_tmp[5]\, B => 
        \ReadFIFO_WR_STATE[5]_net_1\, Y => N_399);
    
    \ReadFIFO_WR_STATE[4]\ : SLE
      port map(D => \ReadFIFO_WR_STATE_ns[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \ReadFIFO_WR_STATE[4]_net_1\);
    
    \ReadFIFO_WR_SM.un29_sm_advance_i_NE_2\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type1_reg(7), B => 
        consumer_type1_reg(6), C => \consumer_type[7]_net_1\, D
         => \consumer_type[6]_net_1\, Y => un29_sm_advance_i_NE_2);
    
    un1_ReadFIFO_WR_STATE_15_0_0_0 : CFG4
      generic map(INIT => x"FFEF")

      port map(A => \ReadFIFO_WR_STATE[9]_net_1\, B => 
        \ReadFIFO_WR_STATE[8]_net_1\, C => N_1475, D => N_1036, Y
         => un1_ReadFIFO_WR_STATE_15);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_6\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[6]_net_1\, B => 
        \un65_sm_advance_i[6]\, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_5, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_6);
    
    rx_end_rst : SLE
      port map(D => N_259_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0_0\, ALn => 
        un2_apb3_reset_i, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rx_end_rst\);
    
    \rx_packet_length_ret[5]\ : SLE
      port map(D => \un56_sm_advance_i_i[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => GND_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \un56_sm_advance_i[6]\);
    
    \rx_fifo_din_d3[2]\ : SLE
      port map(D => N_9, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \N_535\, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RX_FIFO_DIN_pipe[2]\);
    
    \SM_advancebit_cntr[0]\ : SLE
      port map(D => N_174_i_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => un9_rst_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SM_advancebit_cntr[0]_net_1\);
    
    \rx_byte_cntr_lm_0[1]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \ReadFIFO_WR_STATE[1]_net_1\, B => 
        \ReadFIFO_WR_STATE[2]_net_1\, C => N_1358, D => 
        \rx_byte_cntr_s[1]\, Y => \rx_byte_cntr_lm[1]\);
    
    \iRX_FIFO_wr_en\ : SLE
      port map(D => un5_packet_avail, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_996_i, ALn => un16_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        iRX_FIFO_wr_en_net_1);
    
    \rx_packet_length[8]\ : SLE
      port map(D => un56_sm_advance_i_axb_7_i, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \rx_packet_length[8]_net_1\);
    
    \ReadFIFO_WR_STATE_ns[8]\ : CFG4
      generic map(INIT => x"E222")

      port map(A => \ReadFIFO_WR_STATE[1]_net_1\, B => 
        sampler_clk1x_en, C => SM_advance_i_net_1, D => 
        \ReadFIFO_WR_STATE[2]_net_1\, Y => 
        \ReadFIFO_WR_STATE_ns[8]_net_1\);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_1\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[1]_net_1\, B => 
        \un56_sm_advance_i[11]\, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_0, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_1);
    
    \rx_packet_length_ret[2]\ : SLE
      port map(D => \un56_sm_advance_i_i[9]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => GND_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \un56_sm_advance_i[9]\);
    
    \consumer_type[4]\ : SLE
      port map(D => N_820_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_ReadFIFO_WR_STATE_12_0_i_i_a3_0\, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type[4]_net_1\);
    
    \rx_byte_cntr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rx_byte_cntr[8]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \rx_byte_cntr_cry[7]_net_1\, S => \rx_byte_cntr_s[8]\, Y
         => OPEN, FCO => \rx_byte_cntr_cry[8]_net_1\);
    
    \consumer_type_RNO[7]\ : CFG4
      generic map(INIT => x"F088")

      port map(A => RX_FIFO_DIN(5), B => consumer_type_0_sqmuxa, 
        C => \consumer_type[7]_net_1\, D => 
        \ReadFIFO_WR_STATE[8]_net_1\, Y => N_812_i);
    
    \rx_packet_length_ret_1[6]\ : SLE
      port map(D => \un65_sm_advance_i_i[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => GND_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \un65_sm_advance_i[3]\);
    
    \rx_fifo_din_d1[0]\ : SLE
      port map(D => RX_FIFO_DIN(0), CLK => CommsFPGA_CCC_0_GL0, 
        EN => \N_535\, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => N_2);
    
    \rx_byte_cntr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rx_byte_cntr[3]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \rx_byte_cntr_cry[2]_net_1\, S => \rx_byte_cntr_s[3]\, Y
         => OPEN, FCO => \rx_byte_cntr_cry[3]_net_1\);
    
    \ReadFIFO_WR_SM.un38_sm_advance_i_NE_0\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type4_reg(3), B => 
        consumer_type4_reg(2), C => \consumer_type[3]_net_1\, D
         => \consumer_type[2]_net_1\, Y => un38_sm_advance_i_NE_0);
    
    \rx_crc_data_store[1]\ : SLE
      port map(D => \un1_rx_fifo_din_d3[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_41_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[1]_net_1\);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_11\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[11]_net_1\, B => 
        \un65_sm_advance_i[1]\, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_10, S => OPEN, Y => OPEN, 
        FCO => un67_sm_advance_i);
    
    \ReadFIFO_WRITE_PROC.un16_rst\ : CFG2
      generic map(INIT => x"1")

      port map(A => un9_rst, B => \irx_packet_end\, Y => 
        un16_rst_i);
    
    \ReadFIFO_WR_SM.un38_sm_advance_i_7\ : CFG2
      generic map(INIT => x"6")

      port map(A => \consumer_type[7]_net_1\, B => 
        consumer_type4_reg(7), Y => un38_sm_advance_i_7);
    
    consumer_type_0_sqmuxa_0_a3_0_a3_0_a2 : CFG3
      generic map(INIT => x"80")

      port map(A => \ReadFIFO_WR_STATE[9]_net_1\, B => \N_535\, C
         => packet_avail, Y => consumer_type_0_sqmuxa);
    
    un56_sm_advance_i_s_10 : CFG2
      generic map(INIT => x"4")

      port map(A => \un56_sm_advance_i_cry_8\, B => 
        un56_sm_advance_i_s_9_sf, Y => \un56_sm_advance_i_i[1]\);
    
    \rx_byte_cntr_lm_0[0]\ : CFG4
      generic map(INIT => x"0004")

      port map(A => \ReadFIFO_WR_STATE[1]_net_1\, B => N_1358, C
         => \rx_byte_cntr[0]_net_1\, D => 
        \ReadFIFO_WR_STATE[2]_net_1\, Y => \rx_byte_cntr_lm[0]\);
    
    \ReadFIFO_WR_SM.un58_sm_advance_i_0_I_9\ : ARI1
      generic map(INIT => x"68241")

      port map(A => \un56_sm_advance_i[2]\, B => 
        \rx_byte_cntr[10]_net_1\, C => \rx_byte_cntr[11]_net_1\, 
        D => \un56_sm_advance_i[1]\, FCI => 
        \un58_sm_advance_i_0_data_tmp[4]\, S => OPEN, Y => OPEN, 
        FCO => \un58_sm_advance_i_0_data_tmp[5]\);
    
    \un1_rx_fifo_din_d3[4]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \RX_FIFO_DIN_pipe[4]\, B => 
        rx_crc_HighByte_en_net_1, Y => 
        \un1_rx_fifo_din_d3[4]_net_1\);
    
    \rx_byte_cntr_lm_0[6]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \ReadFIFO_WR_STATE[1]_net_1\, B => 
        \ReadFIFO_WR_STATE[2]_net_1\, C => N_1358, D => 
        \rx_byte_cntr_s[6]\, Y => \rx_byte_cntr_lm[6]\);
    
    \rx_fifo_din_d3[4]\ : SLE
      port map(D => N_15, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \N_535\, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RX_FIFO_DIN_pipe[4]\);
    
    \consumer_type[7]\ : SLE
      port map(D => N_812_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_ReadFIFO_WR_STATE_12_0_i_i_a3_0\, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type[7]_net_1\);
    
    \ReadFIFO_WR_STATE_RNO[9]\ : CFG4
      generic map(INIT => x"0EEE")

      port map(A => \ReadFIFO_WR_STATE[9]_net_1\, B => idle_line, 
        C => N_1328, D => N_1358, Y => N_233_i);
    
    RX_InProcess_RNO : CFG2
      generic map(INIT => x"7")

      port map(A => N_1475, B => N_1469, Y => N_250_i);
    
    un65_sm_advance_i_cry_2 : ARI1
      generic map(INIT => x"6FF35")

      port map(A => N_1475, B => RX_FIFO_DIN(3), C => 
        \rx_packet_length[3]_net_1\, D => N_539, FCI => 
        \un65_sm_advance_i_cry_1\, S => \un65_sm_advance_i_i[9]\, 
        Y => OPEN, FCO => \un65_sm_advance_i_cry_2\);
    
    un56_sm_advance_i_s_9_395 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \un56_sm_advance_i_cry_8\, C
         => GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => 
        OPEN, Y => OPEN, FCO => un56_sm_advance_i_s_9_395_FCO);
    
    \rx_fifo_din_d1[5]\ : SLE
      port map(D => RX_FIFO_DIN(5), CLK => CommsFPGA_CCC_0_GL0, 
        EN => \N_535\, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => N_17);
    
    \ReadFIFO_WR_SM.un1_sampler_clk1x_en_0_I_45\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \rx_crc_data_store[9]_net_1\, B => 
        \rx_crc_data_calc[8]\, C => \rx_crc_data_calc[9]\, D => 
        \rx_crc_data_store[8]_net_1\, FCI => 
        \un1_sampler_clk1x_en_0_data_tmp[3]\, S => OPEN, Y => 
        OPEN, FCO => \un1_sampler_clk1x_en_0_data_tmp[4]\);
    
    \rx_crc_data_store[12]\ : SLE
      port map(D => \RX_FIFO_DIN_pipe[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_993_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[12]_net_1\);
    
    \ReadFIFO_WR_STATE_ns_0_0_0[6]\ : CFG4
      generic map(INIT => x"7340")

      port map(A => \un58_sm_advance_i_0_data_tmp[5]\, B => 
        \N_535\, C => \ReadFIFO_WR_STATE[5]_net_1\, D => 
        \ReadFIFO_WR_STATE[3]_net_1\, Y => 
        \ReadFIFO_WR_STATE_ns[6]\);
    
    \rx_crc_HighByte_en\ : SLE
      port map(D => N_399, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0_0\, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        rx_crc_HighByte_en_net_1);
    
    \rx_byte_cntr_lm_0[5]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \ReadFIFO_WR_STATE[1]_net_1\, B => 
        \ReadFIFO_WR_STATE[2]_net_1\, C => N_1358, D => 
        \rx_byte_cntr_s[5]\, Y => \rx_byte_cntr_lm[5]\);
    
    \ReadFIFO_WR_SM.un29_sm_advance_i_NE_7\ : CFG3
      generic map(INIT => x"FE")

      port map(A => un29_sm_advance_i_NE_4, B => 
        un29_sm_advance_i_NE_1, C => un29_sm_advance_i_NE_0, Y
         => un29_sm_advance_i_NE_7);
    
    un56_sm_advance_i_cry_1 : ARI1
      generic map(INIT => x"6FF35")

      port map(A => N_1475, B => RX_FIFO_DIN(2), C => 
        \rx_packet_length[2]_net_1\, D => N_539, FCI => 
        \un56_sm_advance_i_cry_0\, S => \un56_sm_advance_i_i[10]\, 
        Y => OPEN, FCO => \un56_sm_advance_i_cry_1\);
    
    \rx_CRC_error\ : SLE
      port map(D => N_87, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0_0\, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rx_CRC_error_net_1);
    
    \rx_crc_data_store[8]\ : SLE
      port map(D => \RX_FIFO_DIN_pipe[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_993_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[8]_net_1\);
    
    \ReadFIFO_WR_STATE_RNI1PDR[6]\ : CFG4
      generic map(INIT => x"04FF")

      port map(A => \ReadFIFO_WR_STATE[2]_net_1\, B => N_1469, C
         => \ReadFIFO_WR_STATE[6]_net_1\, D => SM_advance_i_net_1, 
        Y => N_992_i_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    un56_sm_advance_i_s_10_RNO : CFG4
      generic map(INIT => x"F5F3")

      port map(A => \rx_packet_length[10]_net_1\, B => 
        RX_FIFO_DIN(2), C => N_1475, D => N_572, Y => 
        un56_sm_advance_i_s_9_sf);
    
    \rx_fifo_din_d1[2]\ : SLE
      port map(D => RX_FIFO_DIN(2), CLK => CommsFPGA_CCC_0_GL0, 
        EN => \N_535\, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => N_8);
    
    \consumer_type[6]\ : SLE
      port map(D => N_74_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_ReadFIFO_WR_STATE_12_0_i_i_a3_0\, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type[6]_net_1\);
    
    \ReadFIFO_WR_STATE_ns_0_0[9]\ : CFG4
      generic map(INIT => x"4F44")

      port map(A => idle_line, B => \ReadFIFO_WR_STATE[0]_net_1\, 
        C => \un1_sampler_clk1x_en_0_data_tmp[7]\, D => 
        \ReadFIFO_WR_STATE_ns_0_0_a2_0_0[9]_net_1\, Y => 
        \ReadFIFO_WR_STATE_ns[9]\);
    
    \rx_crc_data_store[5]\ : SLE
      port map(D => \un1_rx_fifo_din_d3[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_41_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[5]_net_1\);
    
    \ReadFIFO_WR_SM.un1_sampler_clk1x_en_0_I_9\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \rx_crc_data_store[3]_net_1\, B => 
        \rx_crc_data_calc[2]\, C => \rx_crc_data_calc[3]\, D => 
        \rx_crc_data_store[2]_net_1\, FCI => 
        \un1_sampler_clk1x_en_0_data_tmp[0]\, S => OPEN, Y => 
        OPEN, FCO => \un1_sampler_clk1x_en_0_data_tmp[1]\);
    
    \rx_packet_length[6]\ : SLE
      port map(D => un56_sm_advance_i_axb_5_i, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \rx_packet_length[6]_net_1\);
    
    \ReadFIFO_WR_STATE[2]\ : SLE
      port map(D => \ReadFIFO_WR_STATE[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \N_535\, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \ReadFIFO_WR_STATE[2]_net_1\);
    
    \consumer_type_RNO[2]\ : CFG4
      generic map(INIT => x"F088")

      port map(A => RX_FIFO_DIN(0), B => consumer_type_0_sqmuxa, 
        C => \consumer_type[2]_net_1\, D => 
        \ReadFIFO_WR_STATE[8]_net_1\, Y => N_66_i);
    
    \rx_byte_cntr[1]\ : SLE
      port map(D => \rx_byte_cntr_lm[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_992_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_byte_cntr[1]_net_1\);
    
    rx_byte_cntr_s_391 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rx_byte_cntr[0]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => 
        OPEN, Y => OPEN, FCO => rx_byte_cntr_s_391_FCO);
    
    un56_sm_advance_i_cry_4 : ARI1
      generic map(INIT => x"6FF35")

      port map(A => N_1475, B => RX_FIFO_DIN(5), C => 
        \rx_packet_length[5]_net_1\, D => N_539, FCI => 
        \un56_sm_advance_i_cry_3\, S => \un56_sm_advance_i_i[7]\, 
        Y => OPEN, FCO => \un56_sm_advance_i_cry_4\);
    
    \ReadFIFO_WR_SM.un58_sm_advance_i_0_I_1\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \un56_sm_advance_i[11]\, B => 
        \rx_byte_cntr[0]_net_1\, C => \rx_byte_cntr[1]_net_1\, D
         => \rx_packet_length[0]_net_1\, FCI => GND_net_1, S => 
        OPEN, Y => OPEN, FCO => \un58_sm_advance_i_0_data_tmp[0]\);
    
    \ReadFIFO_WR_STATE_ns_0_0_0_o2[4]\ : CFG3
      generic map(INIT => x"7F")

      port map(A => \ReadFIFO_WR_STATE[6]_net_1\, B => 
        SM_advance_i_net_1, C => sampler_clk1x_en, Y => N_539);
    
    \ReadFIFO_WR_SM.un38_sm_advance_i_NE_1\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type4_reg(5), B => 
        consumer_type4_reg(4), C => \consumer_type[5]_net_1\, D
         => \consumer_type[4]_net_1\, Y => un38_sm_advance_i_NE_1);
    
    un65_sm_advance_i_cry_6 : ARI1
      generic map(INIT => x"6FF35")

      port map(A => N_1475, B => RX_FIFO_DIN(7), C => 
        \rx_packet_length[7]_net_1\, D => N_539, FCI => 
        \un65_sm_advance_i_cry_5\, S => \un65_sm_advance_i_i[5]\, 
        Y => OPEN, FCO => \un65_sm_advance_i_cry_6\);
    
    \rx_byte_cntr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rx_byte_cntr[7]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \rx_byte_cntr_cry[6]_net_1\, S => \rx_byte_cntr_s[7]\, Y
         => OPEN, FCO => \rx_byte_cntr_cry[7]_net_1\);
    
    \rx_packet_complt\ : SLE
      port map(D => \rx_packet_complt_1_sqmuxa\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0_0\, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rx_packet_complt);
    
    iRX_EarlyTerm : SLE
      port map(D => \ReadFIFO_WR_STATE[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0_0\, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RX_EarlyTerm\);
    
    \ReadFIFO_WR_SM.un58_sm_advance_i_0_I_21\ : ARI1
      generic map(INIT => x"68241")

      port map(A => \un56_sm_advance_i[6]\, B => 
        \rx_byte_cntr[6]_net_1\, C => \rx_byte_cntr[7]_net_1\, D
         => \un56_sm_advance_i[5]\, FCI => 
        \un58_sm_advance_i_0_data_tmp[2]\, S => OPEN, Y => OPEN, 
        FCO => \un58_sm_advance_i_0_data_tmp[3]\);
    
    \rx_packet_length_ret[8]\ : SLE
      port map(D => \un56_sm_advance_i_i[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => GND_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \un56_sm_advance_i[3]\);
    
    \ReadFIFO_WR_SM.un38_sm_advance_i_NE_4\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type4_reg(1), B => 
        consumer_type4_reg(0), C => \consumer_type[1]_net_1\, D
         => \consumer_type[0]_net_1\, Y => un38_sm_advance_i_NE_4);
    
    un65_sm_advance_i_cry_3 : ARI1
      generic map(INIT => x"6FF35")

      port map(A => N_1475, B => RX_FIFO_DIN(4), C => 
        \rx_packet_length[4]_net_1\, D => N_539, FCI => 
        \un65_sm_advance_i_cry_2\, S => \un65_sm_advance_i_i[8]\, 
        Y => OPEN, FCO => \un65_sm_advance_i_cry_3\);
    
    \ReadFIFO_WR_SM.un1_sampler_clk1x_en_0_I_21\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \rx_crc_data_store[15]_net_1\, B => 
        \rx_crc_data_calc[14]\, C => \rx_crc_data_calc[15]\, D
         => \rx_crc_data_store[14]_net_1\, FCI => 
        \un1_sampler_clk1x_en_0_data_tmp[6]\, S => OPEN, Y => 
        OPEN, FCO => \un1_sampler_clk1x_en_0_data_tmp[7]\);
    
    \bit_cntr[2]\ : SLE
      port map(D => N_151_i_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => un16_rst_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \bit_cntr[2]_net_1\);
    
    \rx_packet_length_ret_1[0]\ : SLE
      port map(D => \un65_sm_advance_i_i[9]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => GND_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \un65_sm_advance_i[9]\);
    
    \bit_cntr[0]\ : SLE
      port map(D => N_1082_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => un16_rst_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \bit_cntr[0]_net_1\);
    
    \ReadFIFO_WR_SM.un29_sm_advance_i_NE_4\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type1_reg(1), B => 
        consumer_type1_reg(0), C => \consumer_type[1]_net_1\, D
         => \consumer_type[0]_net_1\, Y => un29_sm_advance_i_NE_4);
    
    un56_sm_advance_i_cry_3 : ARI1
      generic map(INIT => x"6FF35")

      port map(A => N_1475, B => RX_FIFO_DIN(4), C => 
        \rx_packet_length[4]_net_1\, D => N_539, FCI => 
        \un56_sm_advance_i_cry_2\, S => \un56_sm_advance_i_i[8]\, 
        Y => OPEN, FCO => \un56_sm_advance_i_cry_3\);
    
    \rx_byte_cntr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rx_byte_cntr[4]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \rx_byte_cntr_cry[3]_net_1\, S => \rx_byte_cntr_s[4]\, Y
         => OPEN, FCO => \rx_byte_cntr_cry[4]_net_1\);
    
    \rx_packet_length_ret[1]\ : SLE
      port map(D => \un56_sm_advance_i_i[10]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => GND_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \un56_sm_advance_i[10]\);
    
    \ReadFIFO_WR_SM.un32_sm_advance_i_7\ : CFG2
      generic map(INIT => x"6")

      port map(A => \consumer_type[7]_net_1\, B => 
        consumer_type2_reg(7), Y => un32_sm_advance_i_7);
    
    \rx_packet_length_ret_1[3]\ : SLE
      port map(D => \un65_sm_advance_i_i[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => GND_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \un65_sm_advance_i[6]\);
    
    \rx_packet_length_ret[9]\ : SLE
      port map(D => \un56_sm_advance_i_i[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => GND_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \un56_sm_advance_i[2]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \ReadFIFO_WR_STATE[7]\ : SLE
      port map(D => \ReadFIFO_WR_STATE_202\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \ReadFIFO_WR_STATE[7]_net_1\);
    
    \ReadFIFO_WR_SM.un40_sm_advance_i\ : CFG4
      generic map(INIT => x"E000")

      port map(A => un32_sm_advance_i_NE_6, B => 
        un32_sm_advance_i_NE_7, C => un40_sm_advance_i_1, D => 
        un40_sm_advance_i_0, Y => un40_sm_advance_i);
    
    \rx_fifo_din_d2[6]\ : SLE
      port map(D => N_20, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \N_535\, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        N_21);
    
    \ReadFIFO_WR_SM.un32_sm_advance_i_NE_6\ : CFG4
      generic map(INIT => x"FFF6")

      port map(A => \consumer_type[6]_net_1\, B => 
        consumer_type2_reg(6), C => un32_sm_advance_i_NE_3, D => 
        un32_sm_advance_i_7, Y => un32_sm_advance_i_NE_6);
    
    \ReadFIFO_WR_SM.un38_sm_advance_i_NE_6\ : CFG4
      generic map(INIT => x"FFF6")

      port map(A => \consumer_type[6]_net_1\, B => 
        consumer_type4_reg(6), C => un38_sm_advance_i_NE_3, D => 
        un38_sm_advance_i_7, Y => un38_sm_advance_i_NE_6);
    
    \rx_packet_length[2]\ : SLE
      port map(D => un56_sm_advance_i_axb_1_i, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \rx_packet_length[2]_net_1\);
    
    \rx_byte_cntr_lm_0[9]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \ReadFIFO_WR_STATE[1]_net_1\, B => 
        \ReadFIFO_WR_STATE[2]_net_1\, C => N_1358, D => 
        \rx_byte_cntr_s[9]\, Y => \rx_byte_cntr_lm[9]\);
    
    \rx_fifo_din_d2[0]\ : SLE
      port map(D => N_2, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \N_535\, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        N_3);
    
    \rx_packet_length_ret_1[8]\ : SLE
      port map(D => \un65_sm_advance_i_i[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => GND_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \un65_sm_advance_i[1]\);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_8\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[8]_net_1\, B => 
        \un65_sm_advance_i[4]\, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_7, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_8);
    
    \ReadFIFO_WR_SM.consumer_type_12_i_i_a2_1[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \N_535\, B => \ReadFIFO_WR_STATE[8]_net_1\, Y
         => N_1292);
    
    \SM_advancebit_cntr[1]\ : SLE
      port map(D => N_338_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => un9_rst_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SM_advancebit_cntr[1]_net_1\);
    
    \rx_packet_length_ret[3]\ : SLE
      port map(D => \un56_sm_advance_i_i[8]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => GND_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \un56_sm_advance_i[8]\);
    
    \bit_cntr[1]\ : SLE
      port map(D => N_337_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => un16_rst_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \bit_cntr[1]_net_1\);
    
    \rx_byte_cntr[9]\ : SLE
      port map(D => \rx_byte_cntr_lm[9]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_992_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_byte_cntr[9]_net_1\);
    
    \consumer_type_RNO[6]\ : CFG4
      generic map(INIT => x"F088")

      port map(A => RX_FIFO_DIN(4), B => consumer_type_0_sqmuxa, 
        C => \consumer_type[6]_net_1\, D => 
        \ReadFIFO_WR_STATE[8]_net_1\, Y => N_74_i);
    
    \un1_rx_fifo_din_d3[1]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \RX_FIFO_DIN_pipe[1]\, B => 
        rx_crc_HighByte_en_net_1, Y => 
        \un1_rx_fifo_din_d3[1]_net_1\);
    
    \rx_crc_data_store[13]\ : SLE
      port map(D => \RX_FIFO_DIN_pipe[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_993_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[13]_net_1\);
    
    \rx_crc_data_store[0]\ : SLE
      port map(D => \un1_rx_fifo_din_d3[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_41_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[0]_net_1\);
    
    \rx_byte_cntr_s[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rx_byte_cntr[11]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \rx_byte_cntr_cry[10]_net_1\, S => 
        \rx_byte_cntr_s[11]_net_1\, Y => OPEN, FCO => OPEN);
    
    \rx_byte_cntr_lm_0[10]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \ReadFIFO_WR_STATE[1]_net_1\, B => 
        \ReadFIFO_WR_STATE[2]_net_1\, C => N_1358, D => 
        \rx_byte_cntr_s[10]\, Y => \rx_byte_cntr_lm[10]\);
    
    \ReadFIFO_WR_SM.un38_sm_advance_i_NE\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => un38_sm_advance_i_NE_0, B => 
        un38_sm_advance_i_NE_6, C => un38_sm_advance_i_NE_4, D
         => un38_sm_advance_i_NE_1, Y => un39_sm_advance_i);
    
    \ReadFIFO_WR_SM.un1_sampler_clk1x_en_0_I_15\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \rx_crc_data_store[5]_net_1\, B => 
        \rx_crc_data_calc[4]\, C => \rx_crc_data_calc[5]\, D => 
        \rx_crc_data_store[4]_net_1\, FCI => 
        \un1_sampler_clk1x_en_0_data_tmp[1]\, S => OPEN, Y => 
        OPEN, FCO => \un1_sampler_clk1x_en_0_data_tmp[2]\);
    
    \ReadFIFO_WR_SM.un35_sm_advance_i_NE_0\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type3_reg(3), B => 
        consumer_type3_reg(2), C => \consumer_type[3]_net_1\, D
         => \consumer_type[2]_net_1\, Y => un35_sm_advance_i_NE_0);
    
    \rx_packet_length_ret_1[5]\ : SLE
      port map(D => \un65_sm_advance_i_i[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => GND_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \un65_sm_advance_i[4]\);
    
    \consumer_type[1]\ : SLE
      port map(D => N_1356, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_ReadFIFO_WR_STATE_12_0_i_i_a3_0\, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type[1]_net_1\);
    
    \ReadFIFO_WR_SM.consumer_type_12_i_i[0]\ : CFG4
      generic map(INIT => x"AA0C")

      port map(A => RX_FIFO_DIN(6), B => \consumer_type[0]_net_1\, 
        C => N_1467, D => N_1292, Y => N_313);
    
    \bit_cntr_RNO[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => N_996_i, B => \bit_cntr[0]_net_1\, Y => 
        N_1082_i);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_4\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[4]_net_1\, B => 
        \un65_sm_advance_i[8]\, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_3, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_4);
    
    \rx_fifo_din_d1[4]\ : SLE
      port map(D => RX_FIFO_DIN(4), CLK => CommsFPGA_CCC_0_GL0, 
        EN => \N_535\, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => N_14);
    
    \rx_packet_length_13_i_0_i[1]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => \rx_packet_length[1]_net_1\, B => 
        RX_FIFO_DIN(1), C => N_1475, D => N_539, Y => 
        un56_sm_advance_i_axb_0_i);
    
    \rx_byte_cntr_lm_0[11]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \ReadFIFO_WR_STATE[1]_net_1\, B => 
        \ReadFIFO_WR_STATE[2]_net_1\, C => N_1358, D => 
        \rx_byte_cntr_s[11]_net_1\, Y => \rx_byte_cntr_lm[11]\);
    
    \rx_byte_cntr_lm_0[7]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \ReadFIFO_WR_STATE[1]_net_1\, B => 
        \ReadFIFO_WR_STATE[2]_net_1\, C => N_1358, D => 
        \rx_byte_cntr_s[7]\, Y => \rx_byte_cntr_lm[7]\);
    
    \rx_fifo_din_d2[1]\ : SLE
      port map(D => N_5, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \N_535\, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        N_6);
    
    \rx_packet_length_RNO[10]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => \rx_packet_length[10]_net_1\, B => 
        RX_FIFO_DIN(2), C => N_1475, D => N_572, Y => 
        un56_sm_advance_i_axb_9_i);
    
    \rx_byte_cntr_lm_0[3]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \ReadFIFO_WR_STATE[1]_net_1\, B => 
        \ReadFIFO_WR_STATE[2]_net_1\, C => N_1358, D => 
        \rx_byte_cntr_s[3]\, Y => \rx_byte_cntr_lm[3]\);
    
    \un1_rx_fifo_din_d3[7]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \RX_FIFO_DIN_pipe[7]\, B => 
        rx_crc_HighByte_en_net_1, Y => 
        \un1_rx_fifo_din_d3[7]_net_1\);
    
    \rx_packet_length_RNO[8]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => \rx_packet_length[8]_net_1\, B => 
        RX_FIFO_DIN(0), C => N_1475, D => N_572, Y => 
        un56_sm_advance_i_axb_7_i);
    
    \ReadFIFO_WR_STATE[0]\ : SLE
      port map(D => \ReadFIFO_WR_STATE_ns[9]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \ReadFIFO_WR_STATE[0]_net_1\);
    
    \ReadFIFO_WR_STATE[6]\ : SLE
      port map(D => \ReadFIFO_WR_STATE_ns[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \ReadFIFO_WR_STATE[6]_net_1\);
    
    \rx_fifo_din_d2[5]\ : SLE
      port map(D => N_17, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \N_535\, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        N_18);
    
    \rx_fifo_din_d1[3]\ : SLE
      port map(D => RX_FIFO_DIN(3), CLK => CommsFPGA_CCC_0_GL0, 
        EN => \N_535\, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => N_11);
    
    \un1_rx_fifo_din_d3[0]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \RX_FIFO_DIN_pipe[0]\, B => 
        rx_crc_HighByte_en_net_1, Y => 
        \un1_rx_fifo_din_d3[0]_net_1\);
    
    un1_ReadFIFO_WR_STATE_14_0_0_1 : CFG4
      generic map(INIT => x"CE0A")

      port map(A => N_1333, B => \N_535\, C => 
        \ReadFIFO_WR_STATE[8]_net_1\, D => N_1469, Y => 
        un1_ReadFIFO_WR_STATE_14);
    
    \rx_byte_cntr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rx_byte_cntr[2]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \rx_byte_cntr_cry[1]_net_1\, S => \rx_byte_cntr_s[2]\, Y
         => OPEN, FCO => \rx_byte_cntr_cry[2]_net_1\);
    
    \ReadFIFO_WR_SM.un40_sm_advance_i_1\ : CFG4
      generic map(INIT => x"F0E0")

      port map(A => un35_sm_advance_i_NE_2, B => 
        un35_sm_advance_i_NE_3, C => un39_sm_advance_i, D => 
        un35_sm_advance_i_NE_7, Y => un40_sm_advance_i_1);
    
    \ReadFIFO_WRITE_PROC.un16_rst_0_RNIS9M7\ : CFG1
      generic map(INIT => "01")

      port map(A => un9_rst, Y => un9_rst_i);
    
    \ReadFIFO_WR_STATE_ns_0_0[3]\ : CFG4
      generic map(INIT => x"7520")

      port map(A => \N_535\, B => un40_sm_advance_i, C => 
        \ReadFIFO_WR_STATE[7]_net_1\, D => 
        \ReadFIFO_WR_STATE[6]_net_1\, Y => 
        \ReadFIFO_WR_STATE_ns[3]\);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_9\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[9]_net_1\, B => 
        \un65_sm_advance_i[3]\, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_8, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_9);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_7\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[7]_net_1\, B => 
        \un65_sm_advance_i[5]\, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_6, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_7);
    
    \rx_packet_length_RNO[5]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => \rx_packet_length[5]_net_1\, B => 
        RX_FIFO_DIN(5), C => N_1475, D => N_539, Y => 
        un56_sm_advance_i_axb_4_i);
    
    \consumer_type_RNO[5]\ : CFG4
      generic map(INIT => x"F088")

      port map(A => RX_FIFO_DIN(3), B => consumer_type_0_sqmuxa, 
        C => \consumer_type[5]_net_1\, D => 
        \ReadFIFO_WR_STATE[8]_net_1\, Y => N_72_i);
    
    un1_ReadFIFO_WR_STATE_12_0_i_i_a3_0 : CFG4
      generic map(INIT => x"CDCC")

      port map(A => N_572, B => N_1382, C => 
        \ReadFIFO_WR_STATE[7]_net_1\, D => N_1469, Y => 
        \un1_ReadFIFO_WR_STATE_12_0_i_i_a3_0\);
    
    \rx_packet_length_RNO[7]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => \rx_packet_length[7]_net_1\, B => 
        RX_FIFO_DIN(7), C => N_1475, D => N_539, Y => 
        un56_sm_advance_i_axb_6_i);
    
    \rx_byte_cntr[8]\ : SLE
      port map(D => \rx_byte_cntr_lm[8]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_992_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_byte_cntr[8]_net_1\);
    
    \rx_byte_cntr[2]\ : SLE
      port map(D => \rx_byte_cntr_lm[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_992_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_byte_cntr[2]_net_1\);
    
    \ReadFIFO_WR_SM.un32_sm_advance_i_NE_1\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type2_reg(5), B => 
        consumer_type2_reg(4), C => \consumer_type[5]_net_1\, D
         => \consumer_type[4]_net_1\, Y => un32_sm_advance_i_NE_1);
    
    \rx_packet_length_RNO[9]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => \rx_packet_length[9]_net_1\, B => 
        RX_FIFO_DIN(1), C => N_1475, D => N_572, Y => 
        un56_sm_advance_i_axb_8_i);
    
    \ReadFIFO_WR_SM.un35_sm_advance_i_NE_7\ : CFG3
      generic map(INIT => x"FE")

      port map(A => un35_sm_advance_i_NE_4, B => 
        un35_sm_advance_i_NE_1, C => un35_sm_advance_i_NE_0, Y
         => un35_sm_advance_i_NE_7);
    
    \rx_packet_length[7]\ : SLE
      port map(D => un56_sm_advance_i_axb_6_i, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \rx_packet_length[7]_net_1\);
    
    un1_ReadFIFO_WR_STATE_15_0_0_0_o3_i_a2 : CFG2
      generic map(INIT => x"1")

      port map(A => \ReadFIFO_WR_STATE[6]_net_1\, B => 
        \ReadFIFO_WR_STATE[7]_net_1\, Y => N_1475);
    
    un56_sm_advance_i_cry_0 : ARI1
      generic map(INIT => x"6AEBF")

      port map(A => RX_FIFO_DIN(1), B => N_1475, C => N_539, D
         => \rx_packet_length[1]_net_1\, FCI => GND_net_1, S => 
        OPEN, Y => OPEN, FCO => \un56_sm_advance_i_cry_0\);
    
    \rx_byte_cntr_lm_0[2]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \ReadFIFO_WR_STATE[1]_net_1\, B => 
        \ReadFIFO_WR_STATE[2]_net_1\, C => N_1358, D => 
        \rx_byte_cntr_s[2]\, Y => \rx_byte_cntr_lm[2]\);
    
    rx_end_rst_0_sqmuxa_i_o3_0_0_a2 : CFG2
      generic map(INIT => x"1")

      port map(A => \ReadFIFO_WR_STATE[4]_net_1\, B => 
        \ReadFIFO_WR_STATE[0]_net_1\, Y => N_1328);
    
    \ReadFIFO_WR_SM.un58_sm_advance_i_0_I_15\ : ARI1
      generic map(INIT => x"68241")

      port map(A => \un56_sm_advance_i[10]\, B => 
        \rx_byte_cntr[2]_net_1\, C => \rx_byte_cntr[3]_net_1\, D
         => \un56_sm_advance_i[9]\, FCI => 
        \un58_sm_advance_i_0_data_tmp[0]\, S => OPEN, Y => OPEN, 
        FCO => \un58_sm_advance_i_0_data_tmp[1]\);
    
    RX_InProcess : SLE
      port map(D => N_250_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0_0\, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RX_InProcess\);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_3\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[3]_net_1\, B => 
        \un65_sm_advance_i[9]\, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_2, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_3);
    
    un1_ReadFIFO_WR_STATE_12_0_i_i_a3_0_a2_0 : CFG2
      generic map(INIT => x"8")

      port map(A => N_1333, B => N_1475, Y => N_1382);
    
    \rx_fifo_din_d1[1]\ : SLE
      port map(D => RX_FIFO_DIN(1), CLK => CommsFPGA_CCC_0_GL0, 
        EN => \N_535\, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => N_5);
    
    \ReadFIFO_WR_SM.un38_sm_advance_i_NE_3\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type4_reg(9), B => 
        consumer_type4_reg(8), C => \consumer_type[9]_net_1\, D
         => \consumer_type[8]_net_1\, Y => un38_sm_advance_i_NE_3);
    
    \ReadFIFO_WR_SM.un32_sm_advance_i_NE_0\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type2_reg(3), B => 
        consumer_type2_reg(2), C => \consumer_type[3]_net_1\, D
         => \consumer_type[2]_net_1\, Y => un32_sm_advance_i_NE_0);
    
    un56_sm_advance_i_s_9 : ARI1
      generic map(INIT => x"4FF35")

      port map(A => N_1475, B => RX_FIFO_DIN(2), C => 
        \rx_packet_length[10]_net_1\, D => N_572, FCI => 
        un56_sm_advance_i_s_9_395_FCO, S => 
        \un56_sm_advance_i_i[2]\, Y => OPEN, FCO => OPEN);
    
    \rx_fifo_din_d3[5]\ : SLE
      port map(D => N_18, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \N_535\, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RX_FIFO_DIN_pipe[5]\);
    
    rx_crc_reset : CFG2
      generic map(INIT => x"1")

      port map(A => \rx_end_rst\, B => un2_apb3_reset, Y => 
        \rx_crc_reset\);
    
    \rx_fifo_din_d2[2]\ : SLE
      port map(D => N_8, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \N_535\, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        N_9);
    
    \rx_byte_cntr[0]\ : SLE
      port map(D => \rx_byte_cntr_lm[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_992_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_byte_cntr[0]_net_1\);
    
    \bit_cntr_RNO[2]\ : CFG4
      generic map(INIT => x"78F0")

      port map(A => \bit_cntr[0]_net_1\, B => N_996_i, C => 
        \bit_cntr[2]_net_1\, D => \bit_cntr[1]_net_1\, Y => 
        N_151_i_i);
    
    un1_ReadFIFO_WR_STATE_12_0_i_i_a3_0_a2_1 : CFG2
      generic map(INIT => x"1")

      port map(A => \ReadFIFO_WR_STATE[3]_net_1\, B => 
        \ReadFIFO_WR_STATE[5]_net_1\, Y => N_1469);
    
    \rx_packet_length[0]\ : SLE
      port map(D => N_348_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        un1_ReadFIFO_WR_STATE_14, ALn => un2_apb3_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_packet_length[0]_net_1\);
    
    \ReadFIFO_WR_SM.un29_sm_advance_i_NE_3\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type1_reg(9), B => 
        consumer_type1_reg(8), C => \consumer_type[9]_net_1\, D
         => \consumer_type[8]_net_1\, Y => un29_sm_advance_i_NE_3);
    
    \un1_rx_fifo_din_d3[2]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \RX_FIFO_DIN_pipe[2]\, B => 
        rx_crc_HighByte_en_net_1, Y => 
        \un1_rx_fifo_din_d3[2]_net_1\);
    
    \rx_packet_length_RNO[4]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => \rx_packet_length[4]_net_1\, B => 
        RX_FIFO_DIN(4), C => N_1475, D => N_539, Y => N_43_i);
    
    \rx_crc_data_store[11]\ : SLE
      port map(D => \RX_FIFO_DIN_pipe[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_993_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[11]_net_1\);
    
    \rx_byte_cntr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rx_byte_cntr[1]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        rx_byte_cntr_s_391_FCO, S => \rx_byte_cntr_s[1]\, Y => 
        OPEN, FCO => \rx_byte_cntr_cry[1]_net_1\);
    
    \bit_cntr_RNO[1]\ : CFG3
      generic map(INIT => x"78")

      port map(A => \bit_cntr[0]_net_1\, B => N_996_i, C => 
        \bit_cntr[1]_net_1\, Y => N_337_i);
    
    rx_end_rst_RNO : CFG3
      generic map(INIT => x"E0")

      port map(A => \ReadFIFO_WR_STATE[0]_net_1\, B => 
        \ReadFIFO_WR_STATE[4]_net_1\, C => idle_line, Y => 
        N_259_i);
    
    \ReadFIFO_WR_STATE_ns_0_0_0[4]\ : CFG4
      generic map(INIT => x"8FAF")

      port map(A => \ReadFIFO_WR_STATE[5]_net_1\, B => 
        \un58_sm_advance_i_0_data_tmp[5]\, C => N_539, D => 
        \N_535\, Y => \ReadFIFO_WR_STATE_ns[4]\);
    
    un1_ReadFIFO_WR_STATE_12_0_i_i_a3_0_a2_2 : CFG4
      generic map(INIT => x"3010")

      port map(A => \ReadFIFO_WR_STATE[1]_net_1\, B => 
        \ReadFIFO_WR_STATE[2]_net_1\, C => N_1469, D => 
        sampler_clk1x_en, Y => N_1333);
    
    \rx_crc_data_store[10]\ : SLE
      port map(D => \RX_FIFO_DIN_pipe[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_993_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[10]_net_1\);
    
    \consumer_type_RNO[9]\ : CFG4
      generic map(INIT => x"F088")

      port map(A => RX_FIFO_DIN(7), B => consumer_type_0_sqmuxa, 
        C => \consumer_type[9]_net_1\, D => 
        \ReadFIFO_WR_STATE[8]_net_1\, Y => N_815_i);
    
    \rx_packet_length_ret[7]\ : SLE
      port map(D => \un56_sm_advance_i_i[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => GND_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \un56_sm_advance_i[4]\);
    
    \rx_byte_cntr_lm_0[4]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \ReadFIFO_WR_STATE[1]_net_1\, B => 
        \ReadFIFO_WR_STATE[2]_net_1\, C => N_1358, D => 
        \rx_byte_cntr_s[4]\, Y => \rx_byte_cntr_lm[4]\);
    
    \consumer_type_RNO[8]\ : CFG4
      generic map(INIT => x"F088")

      port map(A => RX_FIFO_DIN(6), B => consumer_type_0_sqmuxa, 
        C => \consumer_type[8]_net_1\, D => 
        \ReadFIFO_WR_STATE[8]_net_1\, Y => N_813_i);
    
    \rx_byte_cntr[10]\ : SLE
      port map(D => \rx_byte_cntr_lm[10]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_992_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_byte_cntr[10]_net_1\);
    
    un65_sm_advance_i_cry_9 : ARI1
      generic map(INIT => x"6FF35")

      port map(A => N_1475, B => RX_FIFO_DIN(2), C => 
        \rx_packet_length[10]_net_1\, D => N_572, FCI => 
        \un65_sm_advance_i_cry_8\, S => \un65_sm_advance_i_i[2]\, 
        Y => OPEN, FCO => \un65_sm_advance_i_cry_9\);
    
    \rx_packet_length_ret_1[2]\ : SLE
      port map(D => \un65_sm_advance_i_i[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => GND_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \un65_sm_advance_i[7]\);
    
    \ReadFIFO_WRITE_PROC.un5_packet_avail_0_a3_0_a3\ : CFG3
      generic map(INIT => x"80")

      port map(A => \bit_cntr[2]_net_1\, B => \bit_cntr[1]_net_1\, 
        C => \bit_cntr[0]_net_1\, Y => un5_packet_avail);
    
    \SM_advancebit_cntr_RNO[2]\ : CFG4
      generic map(INIT => x"78F0")

      port map(A => \SM_advancebit_cntr[0]_net_1\, B => N_996_i, 
        C => \SM_advancebit_cntr[2]_net_1\, D => 
        \SM_advancebit_cntr[1]_net_1\, Y => N_150_i_i);
    
    \rx_crc_data_store[7]\ : SLE
      port map(D => \un1_rx_fifo_din_d3[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_41_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[7]_net_1\);
    
    un56_sm_advance_i_cry_5 : ARI1
      generic map(INIT => x"6FF35")

      port map(A => N_1475, B => RX_FIFO_DIN(6), C => 
        \rx_packet_length[6]_net_1\, D => N_539, FCI => 
        \un56_sm_advance_i_cry_4\, S => \un56_sm_advance_i_i[6]\, 
        Y => OPEN, FCO => \un56_sm_advance_i_cry_5\);
    
    \rx_fifo_din_d1[7]\ : SLE
      port map(D => RX_FIFO_DIN(7), CLK => CommsFPGA_CCC_0_GL0, 
        EN => \N_535\, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => N_23);
    
    \rx_byte_cntr[6]\ : SLE
      port map(D => \rx_byte_cntr_lm[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_992_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_byte_cntr[6]_net_1\);
    
    \consumer_type_RNO[3]\ : CFG4
      generic map(INIT => x"F088")

      port map(A => RX_FIFO_DIN(1), B => consumer_type_0_sqmuxa, 
        C => \consumer_type[3]_net_1\, D => 
        \ReadFIFO_WR_STATE[8]_net_1\, Y => N_819_i);
    
    \ReadFIFO_WR_SM.un35_sm_advance_i_NE_1\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type3_reg(5), B => 
        consumer_type3_reg(4), C => \consumer_type[5]_net_1\, D
         => \consumer_type[4]_net_1\, Y => un35_sm_advance_i_NE_1);
    
    \ReadFIFO_WR_SM.un1_sampler_clk1x_en_0_I_39\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \rx_crc_data_store[13]_net_1\, B => 
        \rx_crc_data_calc[12]\, C => \rx_crc_data_calc[13]\, D
         => \rx_crc_data_store[12]_net_1\, FCI => 
        \un1_sampler_clk1x_en_0_data_tmp[5]\, S => OPEN, Y => 
        OPEN, FCO => \un1_sampler_clk1x_en_0_data_tmp[6]\);
    
    \rx_packet_length_ret_1[4]\ : SLE
      port map(D => \un65_sm_advance_i_i[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => GND_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \un65_sm_advance_i[5]\);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_10\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[10]_net_1\, B => 
        \un65_sm_advance_i[2]\, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_9, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_10);
    
    \ReadFIFO_WR_SM.consumer_type_12_i_i_a2_2[1]\ : CFG2
      generic map(INIT => x"1")

      port map(A => consumer_type_0_sqmuxa, B => 
        \ReadFIFO_WR_STATE[8]_net_1\, Y => N_1467);
    
    \ReadFIFO_WR_STATE[3]\ : SLE
      port map(D => \ReadFIFO_WR_STATE_ns[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \ReadFIFO_WR_STATE[3]_net_1\);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_5\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[5]_net_1\, B => 
        \un65_sm_advance_i[7]\, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_4, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_5);
    
    \ReadFIFO_WRITE_PROC.un16_rst_0\ : CFG3
      generic map(INIT => x"EF")

      port map(A => \RX_EarlyTerm\, B => un2_apb3_reset, C => 
        clk1x_enable, Y => un9_rst);
    
    \ReadFIFO_WR_STATE[1]\ : SLE
      port map(D => \ReadFIFO_WR_STATE_ns[8]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \ReadFIFO_WR_STATE[1]_net_1\);
    
    \ReadFIFO_WR_SM.un29_sm_advance_i_NE_0\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type1_reg(3), B => 
        consumer_type1_reg(2), C => \consumer_type[3]_net_1\, D
         => \consumer_type[2]_net_1\, Y => un29_sm_advance_i_NE_0);
    
    un56_sm_advance_i_cry_7 : ARI1
      generic map(INIT => x"6FF35")

      port map(A => N_1475, B => RX_FIFO_DIN(0), C => 
        \rx_packet_length[8]_net_1\, D => N_572, FCI => 
        \un56_sm_advance_i_cry_6\, S => \un56_sm_advance_i_i[4]\, 
        Y => OPEN, FCO => \un56_sm_advance_i_cry_7\);
    
    \ReadFIFO_WR_STATE[8]\ : SLE
      port map(D => N_321, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ReadFIFO_WR_STATE[8]_net_1\);
    
    \rx_crc_data_store[9]\ : SLE
      port map(D => \RX_FIFO_DIN_pipe[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_993_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[9]_net_1\);
    
    un65_sm_advance_i_cry_4 : ARI1
      generic map(INIT => x"6FF35")

      port map(A => N_1475, B => RX_FIFO_DIN(5), C => 
        \rx_packet_length[5]_net_1\, D => N_539, FCI => 
        \un65_sm_advance_i_cry_3\, S => \un65_sm_advance_i_i[7]\, 
        Y => OPEN, FCO => \un65_sm_advance_i_cry_4\);
    
    \un1_rx_fifo_din_d3[6]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \RX_FIFO_DIN_pipe[6]\, B => 
        rx_crc_HighByte_en_net_1, Y => 
        \un1_rx_fifo_din_d3[6]_net_1\);
    
    \rx_crc_data_store[4]\ : SLE
      port map(D => \un1_rx_fifo_din_d3[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_41_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[4]_net_1\);
    
    \rx_byte_cntr[5]\ : SLE
      port map(D => \rx_byte_cntr_lm[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_992_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_byte_cntr[5]_net_1\);
    
    \rx_fifo_din_d2[7]\ : SLE
      port map(D => N_23, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \N_535\, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        N_24);
    
    \ReadFIFO_WR_SM.un35_sm_advance_i_NE_3\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type3_reg(9), B => 
        consumer_type3_reg(8), C => \consumer_type[9]_net_1\, D
         => \consumer_type[8]_net_1\, Y => un35_sm_advance_i_NE_3);
    
    \un1_rx_fifo_din_d3[3]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \RX_FIFO_DIN_pipe[3]\, B => 
        rx_crc_HighByte_en_net_1, Y => 
        \un1_rx_fifo_din_d3[3]_net_1\);
    
    rx_packet_complt_1_sqmuxa : CFG3
      generic map(INIT => x"20")

      port map(A => idle_line, B => tx_col_detect_en, C => 
        \ReadFIFO_WR_STATE[0]_net_1\, Y => 
        \rx_packet_complt_1_sqmuxa\);
    
    \ReadFIFO_WR_SM.un32_sm_advance_i_NE_4\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type2_reg(1), B => 
        consumer_type2_reg(0), C => \consumer_type[1]_net_1\, D
         => \consumer_type[0]_net_1\, Y => un32_sm_advance_i_NE_4);
    
    \rx_packet_length_ret[10]\ : SLE
      port map(D => \un56_sm_advance_i_i[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => GND_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \un56_sm_advance_i[1]\);
    
    un22_sm_advance_i_0_o2_i_o3_i_i2_0_o2_i_o2 : CFG2
      generic map(INIT => x"8")

      port map(A => sampler_clk1x_en, B => SM_advance_i_net_1, Y
         => \N_535\);
    
    \rx_fifo_din_d3[1]\ : SLE
      port map(D => N_6, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \N_535\, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RX_FIFO_DIN_pipe[1]\);
    
    un65_sm_advance_i_cry_0 : ARI1
      generic map(INIT => x"6FF35")

      port map(A => N_1475, B => RX_FIFO_DIN(1), C => 
        \rx_packet_length[1]_net_1\, D => N_539, FCI => GND_net_1, 
        S => OPEN, Y => un65_sm_advance_i_cry_0_Y, FCO => 
        \un65_sm_advance_i_cry_0\);
    
    \rx_crc_data_store[2]\ : SLE
      port map(D => \un1_rx_fifo_din_d3[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_41_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[2]_net_1\);
    
    \ReadFIFO_WR_SM.un29_sm_advance_i_NE_1\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type1_reg(5), B => 
        consumer_type1_reg(4), C => \consumer_type[5]_net_1\, D
         => \consumer_type[4]_net_1\, Y => un29_sm_advance_i_NE_1);
    
    \rx_packet_length_RNO[2]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => \rx_packet_length[2]_net_1\, B => 
        RX_FIFO_DIN(2), C => N_1475, D => N_539, Y => 
        un56_sm_advance_i_axb_1_i);
    
    \rx_packet_length_ret_1[1]\ : SLE
      port map(D => \un65_sm_advance_i_i[8]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => GND_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \un65_sm_advance_i[8]\);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_2\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[2]_net_1\, B => 
        \un65_sm_advance_i[10]\, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_1, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_2);
    
    \rx_packet_length_ret_1[7]\ : SLE
      port map(D => \un65_sm_advance_i_i[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => GND_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \un65_sm_advance_i[2]\);
    
    \rx_packet_length[4]\ : SLE
      port map(D => N_43_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        un1_ReadFIFO_WR_STATE_14, ALn => un2_apb3_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_packet_length[4]_net_1\);
    
    un65_sm_advance_i_cry_5 : ARI1
      generic map(INIT => x"6FF35")

      port map(A => N_1475, B => RX_FIFO_DIN(6), C => 
        \rx_packet_length[6]_net_1\, D => N_539, FCI => 
        \un65_sm_advance_i_cry_4\, S => \un65_sm_advance_i_i[6]\, 
        Y => OPEN, FCO => \un65_sm_advance_i_cry_5\);
    
    \rx_packet_length[1]\ : SLE
      port map(D => un56_sm_advance_i_axb_0_i, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \rx_packet_length[1]_net_1\);
    
    \rx_byte_cntr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rx_byte_cntr[5]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \rx_byte_cntr_cry[4]_net_1\, S => \rx_byte_cntr_s[5]\, Y
         => OPEN, FCO => \rx_byte_cntr_cry[5]_net_1\);
    
    N_219_i_0_o3_i_o2 : CFG2
      generic map(INIT => x"8")

      port map(A => sampler_clk1x_en, B => packet_avail, Y => 
        N_996_i);
    
    \rx_fifo_din_d2[4]\ : SLE
      port map(D => N_14, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \N_535\, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        N_15);
    
    rx_crc_reset_RNI34TD : CLKINT
      port map(A => \rx_crc_reset\, Y => rx_crc_reset_i);
    
    \ReadFIFO_WR_SM.un1_sampler_clk1x_en_0_I_21_RNIQOK8\ : CFG2
      generic map(INIT => x"8")

      port map(A => \un1_sampler_clk1x_en_0_data_tmp[7]\, B => 
        \ReadFIFO_WR_STATE[1]_net_1\, Y => N_87);
    
    \rx_fifo_din_d2[3]\ : SLE
      port map(D => N_11, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \N_535\, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        N_12);
    
    un65_sm_advance_i_cry_7 : ARI1
      generic map(INIT => x"6FF35")

      port map(A => N_1475, B => RX_FIFO_DIN(0), C => 
        \rx_packet_length[8]_net_1\, D => N_572, FCI => 
        \un65_sm_advance_i_cry_6\, S => \un65_sm_advance_i_i[4]\, 
        Y => OPEN, FCO => \un65_sm_advance_i_cry_7\);
    
    \consumer_type[5]\ : SLE
      port map(D => N_72_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_ReadFIFO_WR_STATE_12_0_i_i_a3_0\, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type[5]_net_1\);
    
    \rx_crc_data_store[14]\ : SLE
      port map(D => \RX_FIFO_DIN_pipe[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_993_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[14]_net_1\);
    
    \ReadFIFO_WR_STATE_ns_0_0[5]\ : CFG4
      generic map(INIT => x"FF80")

      port map(A => \N_535\, B => \ReadFIFO_WR_STATE[7]_net_1\, C
         => un40_sm_advance_i, D => 
        \ReadFIFO_WR_STATE_ns_0_0_0[5]_net_1\, Y => 
        \ReadFIFO_WR_STATE_ns[5]\);
    
    \un1_rx_fifo_din_d3[5]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \RX_FIFO_DIN_pipe[5]\, B => 
        rx_crc_HighByte_en_net_1, Y => 
        \un1_rx_fifo_din_d3[5]_net_1\);
    
    \ReadFIFO_WR_STATE[9]\ : SLE
      port map(D => N_233_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ReadFIFO_WR_STATE[9]_net_1\);
    
    \rx_byte_cntr[4]\ : SLE
      port map(D => \rx_byte_cntr_lm[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_992_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_byte_cntr[4]_net_1\);
    
    \SM_advancebit_cntr[2]\ : SLE
      port map(D => N_150_i_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => un9_rst_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SM_advancebit_cntr[2]_net_1\);
    
    irx_packet_end_RNO : CFG3
      generic map(INIT => x"FE")

      port map(A => \ReadFIFO_WR_STATE[1]_net_1\, B => 
        \ReadFIFO_WR_STATE[0]_net_1\, C => 
        \ReadFIFO_WR_STATE[2]_net_1\, Y => N_669_i);
    
    un1_ReadFIFO_WR_STATE_15_0_0_0_a3 : CFG3
      generic map(INIT => x"20")

      port map(A => \ReadFIFO_WR_STATE[5]_net_1\, B => 
        un67_sm_advance_i, C => \un58_sm_advance_i_0_data_tmp[5]\, 
        Y => N_1036);
    
    \consumer_type[0]\ : SLE
      port map(D => N_313, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_ReadFIFO_WR_STATE_12_0_i_i_a3_0\, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type[0]_net_1\);
    
    RX_CRC_GEN_INST : CRC16_Generator_1
      port map(RX_FIFO_DIN(7) => RX_FIFO_DIN(7), RX_FIFO_DIN(6)
         => RX_FIFO_DIN(6), RX_FIFO_DIN(5) => RX_FIFO_DIN(5), 
        RX_FIFO_DIN(4) => RX_FIFO_DIN(4), RX_FIFO_DIN(3) => 
        RX_FIFO_DIN(3), RX_FIFO_DIN(2) => RX_FIFO_DIN(2), 
        RX_FIFO_DIN(1) => RX_FIFO_DIN(1), RX_FIFO_DIN(0) => 
        RX_FIFO_DIN(0), rx_crc_data_calc(15) => 
        \rx_crc_data_calc[15]\, rx_crc_data_calc(14) => 
        \rx_crc_data_calc[14]\, rx_crc_data_calc(13) => 
        \rx_crc_data_calc[13]\, rx_crc_data_calc(12) => 
        \rx_crc_data_calc[12]\, rx_crc_data_calc(11) => 
        \rx_crc_data_calc[11]\, rx_crc_data_calc(10) => 
        \rx_crc_data_calc[10]\, rx_crc_data_calc(9) => 
        \rx_crc_data_calc[9]\, rx_crc_data_calc(8) => 
        \rx_crc_data_calc[8]\, rx_crc_data_calc(7) => 
        \rx_crc_data_calc[7]\, rx_crc_data_calc(6) => 
        \rx_crc_data_calc[6]\, rx_crc_data_calc(5) => 
        \rx_crc_data_calc[5]\, rx_crc_data_calc(4) => 
        \rx_crc_data_calc[4]\, rx_crc_data_calc(3) => 
        \rx_crc_data_calc[3]\, rx_crc_data_calc(2) => 
        \rx_crc_data_calc[2]\, rx_crc_data_calc(1) => 
        \rx_crc_data_calc[1]\, rx_crc_data_calc(0) => 
        \rx_crc_data_calc[0]\, lfsr_c_i_i_0 => lfsr_c_i_i_0, 
        rx_crc_gen => \rx_crc_gen\, sampler_clk1x_en => 
        sampler_clk1x_en, iRX_FIFO_wr_en => iRX_FIFO_wr_en_net_1, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, 
        rx_crc_reset_i => rx_crc_reset_i);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_0\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[0]_net_1\, B => 
        \rx_packet_length[0]_net_1\, C => GND_net_1, D => 
        GND_net_1, FCI => GND_net_1, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_0);
    
    \rx_fifo_din_d3[7]\ : SLE
      port map(D => N_24, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \N_535\, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RX_FIFO_DIN_pipe[7]\);
    
    un56_sm_advance_i_cry_2 : ARI1
      generic map(INIT => x"6FF35")

      port map(A => N_1475, B => RX_FIFO_DIN(3), C => 
        \rx_packet_length[3]_net_1\, D => N_539, FCI => 
        \un56_sm_advance_i_cry_1\, S => \un56_sm_advance_i_i[9]\, 
        Y => OPEN, FCO => \un56_sm_advance_i_cry_2\);
    
    \rx_packet_length[9]\ : SLE
      port map(D => un56_sm_advance_i_axb_8_i, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \rx_packet_length[9]_net_1\);
    
    \rx_byte_cntr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rx_byte_cntr[6]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \rx_byte_cntr_cry[5]_net_1\, S => \rx_byte_cntr_s[6]\, Y
         => OPEN, FCO => \rx_byte_cntr_cry[6]_net_1\);
    
    rx_packet_length_ret_0 : SLE
      port map(D => \un65_sm_advance_i_i[10]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \un65_sm_advance_i[10]\);
    
    \rx_fifo_din_d3[6]\ : SLE
      port map(D => N_21, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \N_535\, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RX_FIFO_DIN_pipe[6]\);
    
    \consumer_type[9]\ : SLE
      port map(D => N_815_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_ReadFIFO_WR_STATE_12_0_i_i_a3_0\, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type[9]_net_1\);
    
    \ReadFIFO_WR_SM.un1_sampler_clk1x_en_0_I_33\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \rx_crc_data_store[11]_net_1\, B => 
        \rx_crc_data_calc[10]\, C => \rx_crc_data_calc[11]\, D
         => \rx_crc_data_store[10]_net_1\, FCI => 
        \un1_sampler_clk1x_en_0_data_tmp[4]\, S => OPEN, Y => 
        OPEN, FCO => \un1_sampler_clk1x_en_0_data_tmp[5]\);
    
    \rx_crc_data_store[6]\ : SLE
      port map(D => \un1_rx_fifo_din_d3[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_41_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[6]_net_1\);
    
    \rx_packet_length_ret_1_RNO[8]\ : CFG1
      generic map(INIT => "01")

      port map(A => \un65_sm_advance_i_cry_9\, Y => 
        \un65_sm_advance_i_i[1]\);
    
    \SM_advance_i\ : SLE
      port map(D => un2_packet_avail, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_996_i, ALn => un9_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        SM_advance_i_net_1);
    
    un65_sm_advance_i_cry_8 : ARI1
      generic map(INIT => x"6FF35")

      port map(A => N_1475, B => RX_FIFO_DIN(1), C => 
        \rx_packet_length[9]_net_1\, D => N_572, FCI => 
        \un65_sm_advance_i_cry_7\, S => \un65_sm_advance_i_i[3]\, 
        Y => OPEN, FCO => \un65_sm_advance_i_cry_8\);
    
    \ReadFIFO_WR_STATE_ns_0_0_0[5]\ : CFG4
      generic map(INIT => x"F222")

      port map(A => \ReadFIFO_WR_STATE[4]_net_1\, B => idle_line, 
        C => sampler_clk1x_en, D => N_87, Y => 
        \ReadFIFO_WR_STATE_ns_0_0_0[5]_net_1\);
    
    \consumer_type[3]\ : SLE
      port map(D => N_819_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_ReadFIFO_WR_STATE_12_0_i_i_a3_0\, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type[3]_net_1\);
    
    \rx_byte_cntr[3]\ : SLE
      port map(D => \rx_byte_cntr_lm[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_992_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_byte_cntr[3]_net_1\);
    
    \rx_crc_data_store[3]\ : SLE
      port map(D => \un1_rx_fifo_din_d3[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_41_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[3]_net_1\);
    
    \rx_byte_cntr[7]\ : SLE
      port map(D => \rx_byte_cntr_lm[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_992_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_byte_cntr[7]_net_1\);
    
    \rx_packet_length_RNO[6]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => \rx_packet_length[6]_net_1\, B => 
        RX_FIFO_DIN(6), C => N_1475, D => N_539, Y => 
        un56_sm_advance_i_axb_5_i);
    
    \RX_InProcess_d1\ : SLE
      port map(D => \RX_InProcess\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => un2_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RX_InProcess_d1);
    
    \ReadFIFO_WR_STATE_ns_i_0_0_o2_RNIPT5I1[0]\ : CFG4
      generic map(INIT => x"F733")

      port map(A => N_992_i_1, B => N_1358, C => 
        \ReadFIFO_WR_STATE[1]_net_1\, D => sampler_clk1x_en, Y
         => N_992_i);
    
    \consumer_type[8]\ : SLE
      port map(D => N_813_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_ReadFIFO_WR_STATE_12_0_i_i_a3_0\, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type[8]_net_1\);
    
    \rx_packet_length_RNO[3]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => \rx_packet_length[3]_net_1\, B => 
        RX_FIFO_DIN(3), C => N_1475, D => N_539, Y => 
        un56_sm_advance_i_axb_2_i);
    
    \rx_packet_length[3]\ : SLE
      port map(D => un56_sm_advance_i_axb_2_i, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \rx_packet_length[3]_net_1\);
    
    \SM_advancebit_cntr_RNO[1]\ : CFG3
      generic map(INIT => x"78")

      port map(A => \SM_advancebit_cntr[0]_net_1\, B => N_996_i, 
        C => \SM_advancebit_cntr[1]_net_1\, Y => N_338_i);
    
    \rx_packet_length_ret[6]\ : SLE
      port map(D => \un56_sm_advance_i_i[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => un2_apb3_reset_i, ADn => GND_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \un56_sm_advance_i[5]\);
    
    irx_packet_end : SLE
      port map(D => N_669_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0_0\, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \irx_packet_end\);
    
    rx_crc_gen : SLE
      port map(D => un1_ReadFIFO_WR_STATE_15, CLK => 
        CommsFPGA_CCC_0_GL0, EN => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0_0\, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rx_crc_gen\);
    
    \rx_fifo_din_d1[6]\ : SLE
      port map(D => RX_FIFO_DIN(6), CLK => CommsFPGA_CCC_0_GL0, 
        EN => \N_535\, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => N_20);
    
    \rx_fifo_din_d3[3]\ : SLE
      port map(D => N_12, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \N_535\, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RX_FIFO_DIN_pipe[3]\);
    
    \rx_fifo_din_d3[0]\ : SLE
      port map(D => N_3, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \N_535\, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RX_FIFO_DIN_pipe[0]\);
    
    \ReadFIFO_WR_STATE[5]\ : SLE
      port map(D => \ReadFIFO_WR_STATE_ns[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \ReadFIFO_WR_STATE[5]_net_1\);
    
    \ReadFIFO_WR_SM.un1_sampler_clk1x_en_0_I_1\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \rx_crc_data_store[1]_net_1\, B => 
        \rx_crc_data_calc[0]\, C => \rx_crc_data_calc[1]\, D => 
        \rx_crc_data_store[0]_net_1\, FCI => GND_net_1, S => OPEN, 
        Y => OPEN, FCO => \un1_sampler_clk1x_en_0_data_tmp[0]\);
    
    un65_sm_advance_i_cry_1 : ARI1
      generic map(INIT => x"400CA")

      port map(A => N_1475, B => RX_FIFO_DIN(2), C => 
        \rx_packet_length[2]_net_1\, D => N_539, FCI => 
        \un65_sm_advance_i_cry_0\, S => \un65_sm_advance_i_i[10]\, 
        Y => OPEN, FCO => \un65_sm_advance_i_cry_1\);
    
    \ReadFIFO_WR_STATE_ns_i_0_0_o2[0]\ : CFG3
      generic map(INIT => x"D5")

      port map(A => \ReadFIFO_WR_STATE[9]_net_1\, B => \N_535\, C
         => packet_avail, Y => N_1358);
    
    \ReadFIFO_WR_SM.un1_sampler_clk1x_en_0_I_27\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \rx_crc_data_store[7]_net_1\, B => 
        \rx_crc_data_calc[6]\, C => \rx_crc_data_calc[7]\, D => 
        \rx_crc_data_store[6]_net_1\, FCI => 
        \un1_sampler_clk1x_en_0_data_tmp[2]\, S => OPEN, Y => 
        OPEN, FCO => \un1_sampler_clk1x_en_0_data_tmp[3]\);
    
    \consumer_type[2]\ : SLE
      port map(D => N_66_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_ReadFIFO_WR_STATE_12_0_i_i_a3_0\, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type[2]_net_1\);
    
    \rx_crc_data_store[15]\ : SLE
      port map(D => \RX_FIFO_DIN_pipe[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_993_i, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[15]_net_1\);
    
    rx_CRC_error_RNIASV4 : CFG1
      generic map(INIT => "01")

      port map(A => rx_CRC_error_net_1, Y => rx_CRC_error_i);
    
    \ReadFIFO_WR_SM.un32_sm_advance_i_NE_3\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type2_reg(9), B => 
        consumer_type2_reg(8), C => \consumer_type[9]_net_1\, D
         => \consumer_type[8]_net_1\, Y => un32_sm_advance_i_NE_3);
    
    \rx_packet_length_RNO[0]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => \rx_packet_length[0]_net_1\, B => 
        RX_FIFO_DIN(0), C => N_1475, D => N_539, Y => N_348_i);
    
    \ReadFIFO_WR_STATE_ns_0_0_a2_0_0[9]\ : CFG2
      generic map(INIT => x"8")

      port map(A => sampler_clk1x_en, B => 
        \ReadFIFO_WR_STATE[1]_net_1\, Y => 
        \ReadFIFO_WR_STATE_ns_0_0_a2_0_0[9]_net_1\);
    
    \ReadFIFO_WR_STATE_ns_0_i_i[1]\ : CFG3
      generic map(INIT => x"AE")

      port map(A => consumer_type_0_sqmuxa, B => 
        \ReadFIFO_WR_STATE[8]_net_1\, C => \N_535\, Y => N_321);
    
    \ReadFIFO_WR_SM.un40_sm_advance_i_0\ : CFG4
      generic map(INIT => x"3332")

      port map(A => un29_sm_advance_i_NE_3, B => DRVR_EN_c, C => 
        un29_sm_advance_i_NE_7, D => un29_sm_advance_i_NE_2, Y
         => un40_sm_advance_i_0);
    
    \ReadFIFO_WR_SM.un35_sm_advance_i_NE_2\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type3_reg(7), B => 
        consumer_type3_reg(6), C => \consumer_type[7]_net_1\, D
         => \consumer_type[6]_net_1\, Y => un35_sm_advance_i_NE_2);
    
    \SM_ADVANCE_PROC.un2_packet_avail_0_a3_0_a3\ : CFG3
      generic map(INIT => x"80")

      port map(A => \SM_advancebit_cntr[2]_net_1\, B => 
        \SM_advancebit_cntr[1]_net_1\, C => 
        \SM_advancebit_cntr[0]_net_1\, Y => un2_packet_avail);
    
    \rx_byte_cntr_lm_0[8]\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \ReadFIFO_WR_STATE[1]_net_1\, B => 
        \ReadFIFO_WR_STATE[2]_net_1\, C => N_1358, D => 
        \rx_byte_cntr_s[8]\, Y => \rx_byte_cntr_lm[8]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity AFE_RX_SM is

    port( RX_FIFO_DIN         : in    std_logic_vector(7 downto 0);
          manches_in_dly      : in    std_logic_vector(1 downto 0);
          irx_center_sample   : in    std_logic;
          idle_line           : in    std_logic;
          RX_EarlyTerm        : in    std_logic;
          un2_apb3_reset      : in    std_logic;
          clk1x_enable        : out   std_logic;
          packet_avail        : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          un2_apb3_reset_i    : in    std_logic;
          rx_packet_end_all   : out   std_logic
        );

end AFE_RX_SM;

architecture DEF_ARCH of AFE_RX_SM is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \rx_packet_end_all\, VCC_net_1, irx_packet_end_all_5, 
        GND_net_1, \packet_avail_6_0_i_i\, clk1x_enable_1, 
        \start_bit_mask\, start_bit_cntre, \start_bit_maskce\, 
        \RX_EarlyTerm_s\, \RX_EarlyTerm_s_0\, 
        \AFE_RX_STATE[4]_net_1\, N_77_i, \AFE_RX_STATE[3]_net_1\, 
        \AFE_RX_STATE_ns[1]\, \AFE_RX_STATE[2]_net_1\, 
        \AFE_RX_STATE_ns[2]_net_1\, \AFE_RX_STATE[1]_net_1\, 
        \AFE_RX_STATE_ns_i_a3_i[3]_net_1\, 
        \start_bit_cntr[0]_net_1\, \start_bit_cntr_s[0]\, 
        \start_bit_cntr[1]_net_1\, \start_bit_cntr_s[1]\, 
        \start_bit_cntr[2]_net_1\, \start_bit_cntr_s[2]\, 
        \start_bit_cntr[3]_net_1\, \start_bit_cntr_s[3]\, 
        \start_bit_cntr[4]_net_1\, \start_bit_cntr_s[4]\, 
        \start_bit_cntr[5]_net_1\, \start_bit_cntr_s[5]\, 
        \start_bit_cntr[6]_net_1\, \start_bit_cntr_s[6]\, 
        \start_bit_cntr[7]_net_1\, \start_bit_cntr_s[7]_net_1\, 
        start_bit_cntr_cry_cy, N_1058_i, 
        \start_bit_cntr_cry[0]_net_1\, 
        \start_bit_cntr_cry[1]_net_1\, 
        \start_bit_cntr_cry[2]_net_1\, 
        \start_bit_cntr_cry[3]_net_1\, 
        \start_bit_cntr_cry[4]_net_1\, 
        \start_bit_cntr_cry[5]_net_1\, 
        \start_bit_cntr_cry[6]_net_1\, 
        \packet_avail_6_0_i_i_a2_0_0\, 
        \packet_avail_6_0_i_i_a2_0_7\, 
        \packet_avail_6_0_i_i_a2_0_6\, un2_sample_5, un2_sample_4, 
        N_1374 : std_logic;

begin 

    rx_packet_end_all <= \rx_packet_end_all\;

    \start_bit_cntr[2]\ : SLE
      port map(D => \start_bit_cntr_s[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => start_bit_cntre, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \start_bit_cntr[2]_net_1\);
    
    RX_EarlyTerm_s_0 : CFG2
      generic map(INIT => x"4")

      port map(A => un2_apb3_reset, B => RX_EarlyTerm, Y => 
        \RX_EarlyTerm_s_0\);
    
    \START_BIT_COUNTER_PROC.un5_reset_i_a3\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \AFE_RX_STATE[4]_net_1\, B => un2_apb3_reset, 
        C => \rx_packet_end_all\, Y => N_1058_i);
    
    \AFE_RX_STATE[3]\ : SLE
      port map(D => \AFE_RX_STATE_ns[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \AFE_RX_STATE[3]_net_1\);
    
    \AFE_RX_STATE_ns[2]\ : CFG4
      generic map(INIT => x"00CE")

      port map(A => \AFE_RX_STATE[2]_net_1\, B => 
        \AFE_RX_STATE[3]_net_1\, C => N_1374, D => idle_line, Y
         => \AFE_RX_STATE_ns[2]_net_1\);
    
    \start_bit_cntr[5]\ : SLE
      port map(D => \start_bit_cntr_s[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => start_bit_cntre, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \start_bit_cntr[5]_net_1\);
    
    packet_avail_6_0_i_i_a2_0_6 : CFG4
      generic map(INIT => x"0010")

      port map(A => idle_line, B => RX_FIFO_DIN(5), C => 
        RX_FIFO_DIN(4), D => RX_FIFO_DIN(3), Y => 
        \packet_avail_6_0_i_i_a2_0_6\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \start_bit_cntr_cry_cy[0]\ : ARI1
      generic map(INIT => x"45500")

      port map(A => VCC_net_1, B => N_1058_i, C => GND_net_1, D
         => GND_net_1, FCI => VCC_net_1, S => OPEN, Y => OPEN, 
        FCO => start_bit_cntr_cry_cy);
    
    packet_avail_6_0_i_i_a2_0 : CFG4
      generic map(INIT => x"0800")

      port map(A => \packet_avail_6_0_i_i_a2_0_6\, B => 
        \packet_avail_6_0_i_i_a2_0_7\, C => RX_FIFO_DIN(1), D => 
        \packet_avail_6_0_i_i_a2_0_0\, Y => N_1374);
    
    start_bit_maskce : CFG2
      generic map(INIT => x"E")

      port map(A => N_1058_i, B => irx_center_sample, Y => 
        \start_bit_maskce\);
    
    \start_bit_cntr[3]\ : SLE
      port map(D => \start_bit_cntr_s[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => start_bit_cntre, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \start_bit_cntr[3]_net_1\);
    
    \start_bit_cntr_cry[5]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => N_1058_i, C => 
        \start_bit_cntr[5]_net_1\, D => GND_net_1, FCI => 
        \start_bit_cntr_cry[4]_net_1\, S => \start_bit_cntr_s[5]\, 
        Y => OPEN, FCO => \start_bit_cntr_cry[5]_net_1\);
    
    \AFE_RX_STATE_ns_a3[1]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \AFE_RX_STATE[4]_net_1\, B => 
        manches_in_dly(0), C => manches_in_dly(1), Y => 
        \AFE_RX_STATE_ns[1]\);
    
    \start_bit_cntr_cry[0]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => N_1058_i, C => 
        \start_bit_cntr[0]_net_1\, D => GND_net_1, FCI => 
        start_bit_cntr_cry_cy, S => \start_bit_cntr_s[0]\, Y => 
        OPEN, FCO => \start_bit_cntr_cry[0]_net_1\);
    
    \AFE_RX_STATE[1]\ : SLE
      port map(D => \AFE_RX_STATE_ns_i_a3_i[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \AFE_RX_STATE[1]_net_1\);
    
    clk1x_enable_1_0 : CFG4
      generic map(INIT => x"0F1F")

      port map(A => \AFE_RX_STATE[2]_net_1\, B => 
        \AFE_RX_STATE[3]_net_1\, C => N_77_i, D => 
        \AFE_RX_STATE[4]_net_1\, Y => clk1x_enable_1);
    
    \AFE_RX_STATE[4]\ : SLE
      port map(D => N_77_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \AFE_RX_STATE[4]_net_1\);
    
    packet_avail_6_0_i_i_a2_0_7 : CFG4
      generic map(INIT => x"8000")

      port map(A => RX_FIFO_DIN(6), B => RX_FIFO_DIN(7), C => 
        RX_FIFO_DIN(2), D => RX_FIFO_DIN(0), Y => 
        \packet_avail_6_0_i_i_a2_0_7\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \start_bit_cntr[0]\ : SLE
      port map(D => \start_bit_cntr_s[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => start_bit_cntre, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \start_bit_cntr[0]_net_1\);
    
    RX_EarlyTerm_s : SLE
      port map(D => \RX_EarlyTerm_s_0\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RX_EarlyTerm_s\);
    
    \start_bit_cntr[1]\ : SLE
      port map(D => \start_bit_cntr_s[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => start_bit_cntre, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \start_bit_cntr[1]_net_1\);
    
    packet_avail_6_0_i_i_a2_0_0 : CFG2
      generic map(INIT => x"2")

      port map(A => \AFE_RX_STATE[2]_net_1\, B => 
        \start_bit_mask\, Y => \packet_avail_6_0_i_i_a2_0_0\);
    
    \start_bit_cntr[4]\ : SLE
      port map(D => \start_bit_cntr_s[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => start_bit_cntre, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \start_bit_cntr[4]_net_1\);
    
    \AFE_RX_SM.irx_packet_end_all_5_0_a3_0_a3\ : CFG3
      generic map(INIT => x"10")

      port map(A => \AFE_RX_STATE[1]_net_1\, B => 
        \AFE_RX_STATE[4]_net_1\, C => idle_line, Y => 
        irx_packet_end_all_5);
    
    \start_bit_cntr_s[7]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => N_1058_i, C => 
        \start_bit_cntr[7]_net_1\, D => GND_net_1, FCI => 
        \start_bit_cntr_cry[6]_net_1\, S => 
        \start_bit_cntr_s[7]_net_1\, Y => OPEN, FCO => OPEN);
    
    start_bit_mask_1 : CFG4
      generic map(INIT => x"FF2A")

      port map(A => irx_center_sample, B => un2_sample_5, C => 
        un2_sample_4, D => N_1058_i, Y => start_bit_cntre);
    
    \START_BIT_COUNTER_PROC.un2_sample_5\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \start_bit_cntr[4]_net_1\, B => 
        \start_bit_cntr[3]_net_1\, C => \start_bit_cntr[1]_net_1\, 
        D => \start_bit_cntr[0]_net_1\, Y => un2_sample_5);
    
    \start_bit_cntr_cry[6]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => N_1058_i, C => 
        \start_bit_cntr[6]_net_1\, D => GND_net_1, FCI => 
        \start_bit_cntr_cry[5]_net_1\, S => \start_bit_cntr_s[6]\, 
        Y => OPEN, FCO => \start_bit_cntr_cry[6]_net_1\);
    
    \start_bit_cntr[6]\ : SLE
      port map(D => \start_bit_cntr_s[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => start_bit_cntre, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \start_bit_cntr[6]_net_1\);
    
    \AFE_RX_STATE_ns_i_o3[0]\ : CFG3
      generic map(INIT => x"54")

      port map(A => \AFE_RX_STATE_ns[1]\, B => 
        \AFE_RX_STATE[4]_net_1\, C => idle_line, Y => N_77_i);
    
    \packet_avail\ : SLE
      port map(D => \packet_avail_6_0_i_i\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => packet_avail);
    
    irx_packet_end_all : SLE
      port map(D => irx_packet_end_all_5, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rx_packet_end_all\);
    
    \start_bit_cntr_cry[3]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => N_1058_i, C => 
        \start_bit_cntr[3]_net_1\, D => GND_net_1, FCI => 
        \start_bit_cntr_cry[2]_net_1\, S => \start_bit_cntr_s[3]\, 
        Y => OPEN, FCO => \start_bit_cntr_cry[3]_net_1\);
    
    \AFE_RX_STATE[2]\ : SLE
      port map(D => \AFE_RX_STATE_ns[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \AFE_RX_STATE[2]_net_1\);
    
    \start_bit_cntr_cry[2]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => N_1058_i, C => 
        \start_bit_cntr[2]_net_1\, D => GND_net_1, FCI => 
        \start_bit_cntr_cry[1]_net_1\, S => \start_bit_cntr_s[2]\, 
        Y => OPEN, FCO => \start_bit_cntr_cry[2]_net_1\);
    
    \start_bit_cntr[7]\ : SLE
      port map(D => \start_bit_cntr_s[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => start_bit_cntre, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \start_bit_cntr[7]_net_1\);
    
    start_bit_mask : SLE
      port map(D => start_bit_cntre, CLK => CommsFPGA_CCC_0_GL0, 
        EN => \start_bit_maskce\, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \start_bit_mask\);
    
    packet_avail_6_0_i_i : CFG4
      generic map(INIT => x"FAF2")

      port map(A => \AFE_RX_STATE[1]_net_1\, B => 
        \RX_EarlyTerm_s\, C => N_1374, D => idle_line, Y => 
        \packet_avail_6_0_i_i\);
    
    \start_bit_cntr_cry[4]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => N_1058_i, C => 
        \start_bit_cntr[4]_net_1\, D => GND_net_1, FCI => 
        \start_bit_cntr_cry[3]_net_1\, S => \start_bit_cntr_s[4]\, 
        Y => OPEN, FCO => \start_bit_cntr_cry[4]_net_1\);
    
    \start_bit_cntr_cry[1]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => N_1058_i, C => 
        \start_bit_cntr[1]_net_1\, D => GND_net_1, FCI => 
        \start_bit_cntr_cry[0]_net_1\, S => \start_bit_cntr_s[1]\, 
        Y => OPEN, FCO => \start_bit_cntr_cry[1]_net_1\);
    
    \AFE_RX_STATE_ns_i_a3_i[3]\ : CFG4
      generic map(INIT => x"F0F2")

      port map(A => \AFE_RX_STATE[1]_net_1\, B => 
        \RX_EarlyTerm_s\, C => N_1374, D => idle_line, Y => 
        \AFE_RX_STATE_ns_i_a3_i[3]_net_1\);
    
    \clk1x_enable\ : SLE
      port map(D => clk1x_enable_1, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => un2_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => clk1x_enable);
    
    \START_BIT_COUNTER_PROC.un2_sample_4\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \start_bit_cntr[7]_net_1\, B => 
        \start_bit_cntr[6]_net_1\, C => \start_bit_cntr[5]_net_1\, 
        D => \start_bit_cntr[2]_net_1\, Y => un2_sample_4);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity ManchesDecoder is

    port( RX_FIFO_DIN_pipe    : out   std_logic_vector(8 downto 0);
          rx_crc_data_calc    : out   std_logic_vector(11 downto 10);
          consumer_type1_reg  : in    std_logic_vector(9 downto 0);
          consumer_type3_reg  : in    std_logic_vector(9 downto 0);
          consumer_type4_reg  : in    std_logic_vector(9 downto 0);
          consumer_type2_reg  : in    std_logic_vector(9 downto 0);
          manches_in_dly      : out   std_logic_vector(1 downto 0);
          RX_FIFO_DIN         : out   std_logic_vector(3 downto 2);
          lfsr_c_i_i_0        : in    std_logic;
          rx_CRC_error        : out   std_logic;
          rx_CRC_error_i      : out   std_logic;
          N_993_i             : in    std_logic;
          N_41_i              : in    std_logic;
          iRX_FIFO_wr_en      : out   std_logic;
          rx_crc_HighByte_en  : out   std_logic;
          SM_advance_i        : out   std_logic;
          N_535               : out   std_logic;
          rx_packet_complt    : out   std_logic;
          RX_InProcess_d1     : out   std_logic;
          tx_col_detect_en    : in    std_logic;
          DRVR_EN_c           : in    std_logic;
          RX_EarlyTerm        : out   std_logic;
          un2_apb3_reset_i    : in    std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          sampler_clk1x_en    : out   std_logic;
          MANCH_OUT_P_c       : in    std_logic;
          MANCHESTER_IN_c     : in    std_logic;
          internal_loopback   : in    std_logic;
          un2_apb3_reset      : in    std_logic;
          idle_line5          : in    std_logic
        );

end ManchesDecoder;

architecture DEF_ARCH of ManchesDecoder is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component ManchesDecoder_Adapter
    port( RX_FIFO_DIN         : out   std_logic_vector(7 downto 0);
          manches_in_dly      : out   std_logic_vector(1 downto 0);
          idle_line5          : in    std_logic := 'U';
          un2_apb3_reset      : in    std_logic := 'U';
          internal_loopback   : in    std_logic := 'U';
          MANCHESTER_IN_c     : in    std_logic := 'U';
          MANCH_OUT_P_c       : in    std_logic := 'U';
          rx_packet_end_all   : in    std_logic := 'U';
          idle_line           : out   std_logic;
          irx_center_sample   : out   std_logic;
          sampler_clk1x_en    : out   std_logic;
          clk1x_enable        : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          un2_apb3_reset_i    : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component ReadFIFO_Write_SM
    port( consumer_type2_reg  : in    std_logic_vector(9 downto 0) := (others => 'U');
          consumer_type4_reg  : in    std_logic_vector(9 downto 0) := (others => 'U');
          consumer_type3_reg  : in    std_logic_vector(9 downto 0) := (others => 'U');
          consumer_type1_reg  : in    std_logic_vector(9 downto 0) := (others => 'U');
          rx_crc_data_calc    : out   std_logic_vector(11 downto 10);
          RX_FIFO_DIN         : in    std_logic_vector(7 downto 0) := (others => 'U');
          RX_FIFO_DIN_pipe    : out   std_logic_vector(8 downto 0);
          lfsr_c_i_i_0        : in    std_logic := 'U';
          DRVR_EN_c           : in    std_logic := 'U';
          clk1x_enable        : in    std_logic := 'U';
          un2_apb3_reset      : in    std_logic := 'U';
          tx_col_detect_en    : in    std_logic := 'U';
          packet_avail        : in    std_logic := 'U';
          sampler_clk1x_en    : in    std_logic := 'U';
          idle_line           : in    std_logic := 'U';
          RX_InProcess_d1     : out   std_logic;
          rx_packet_complt    : out   std_logic;
          N_535               : out   std_logic;
          RX_EarlyTerm        : out   std_logic;
          SM_advance_i        : out   std_logic;
          rx_crc_HighByte_en  : out   std_logic;
          iRX_FIFO_wr_en      : out   std_logic;
          N_41_i              : in    std_logic := 'U';
          N_993_i             : in    std_logic := 'U';
          un2_apb3_reset_i    : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          rx_CRC_error_i      : out   std_logic;
          rx_CRC_error        : out   std_logic
        );
  end component;

  component AFE_RX_SM
    port( RX_FIFO_DIN         : in    std_logic_vector(7 downto 0) := (others => 'U');
          manches_in_dly      : in    std_logic_vector(1 downto 0) := (others => 'U');
          irx_center_sample   : in    std_logic := 'U';
          idle_line           : in    std_logic := 'U';
          RX_EarlyTerm        : in    std_logic := 'U';
          un2_apb3_reset      : in    std_logic := 'U';
          clk1x_enable        : out   std_logic;
          packet_avail        : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          un2_apb3_reset_i    : in    std_logic := 'U';
          rx_packet_end_all   : out   std_logic
        );
  end component;

    signal \RX_FIFO_DIN[0]\, \RX_FIFO_DIN[1]\, \RX_FIFO_DIN[2]\, 
        \RX_FIFO_DIN[3]\, \RX_FIFO_DIN[4]\, \RX_FIFO_DIN[5]\, 
        \RX_FIFO_DIN[6]\, \RX_FIFO_DIN[7]\, \manches_in_dly[0]\, 
        \manches_in_dly[1]\, rx_packet_end_all, idle_line, 
        irx_center_sample, \sampler_clk1x_en\, clk1x_enable, 
        \RX_EarlyTerm\, packet_avail, GND_net_1, VCC_net_1
         : std_logic;

    for all : ManchesDecoder_Adapter
	Use entity work.ManchesDecoder_Adapter(DEF_ARCH);
    for all : ReadFIFO_Write_SM
	Use entity work.ReadFIFO_Write_SM(DEF_ARCH);
    for all : AFE_RX_SM
	Use entity work.AFE_RX_SM(DEF_ARCH);
begin 

    manches_in_dly(1) <= \manches_in_dly[1]\;
    manches_in_dly(0) <= \manches_in_dly[0]\;
    RX_FIFO_DIN(3) <= \RX_FIFO_DIN[3]\;
    RX_FIFO_DIN(2) <= \RX_FIFO_DIN[2]\;
    RX_EarlyTerm <= \RX_EarlyTerm\;
    sampler_clk1x_en <= \sampler_clk1x_en\;

    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    MANCHESTER_DECODER_ADAPTER_INST : ManchesDecoder_Adapter
      port map(RX_FIFO_DIN(7) => \RX_FIFO_DIN[7]\, RX_FIFO_DIN(6)
         => \RX_FIFO_DIN[6]\, RX_FIFO_DIN(5) => \RX_FIFO_DIN[5]\, 
        RX_FIFO_DIN(4) => \RX_FIFO_DIN[4]\, RX_FIFO_DIN(3) => 
        \RX_FIFO_DIN[3]\, RX_FIFO_DIN(2) => \RX_FIFO_DIN[2]\, 
        RX_FIFO_DIN(1) => \RX_FIFO_DIN[1]\, RX_FIFO_DIN(0) => 
        \RX_FIFO_DIN[0]\, manches_in_dly(1) => 
        \manches_in_dly[1]\, manches_in_dly(0) => 
        \manches_in_dly[0]\, idle_line5 => idle_line5, 
        un2_apb3_reset => un2_apb3_reset, internal_loopback => 
        internal_loopback, MANCHESTER_IN_c => MANCHESTER_IN_c, 
        MANCH_OUT_P_c => MANCH_OUT_P_c, rx_packet_end_all => 
        rx_packet_end_all, idle_line => idle_line, 
        irx_center_sample => irx_center_sample, sampler_clk1x_en
         => \sampler_clk1x_en\, clk1x_enable => clk1x_enable, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, 
        un2_apb3_reset_i => un2_apb3_reset_i);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    ReadFIFO_Write_SM_PROC : ReadFIFO_Write_SM
      port map(consumer_type2_reg(9) => consumer_type2_reg(9), 
        consumer_type2_reg(8) => consumer_type2_reg(8), 
        consumer_type2_reg(7) => consumer_type2_reg(7), 
        consumer_type2_reg(6) => consumer_type2_reg(6), 
        consumer_type2_reg(5) => consumer_type2_reg(5), 
        consumer_type2_reg(4) => consumer_type2_reg(4), 
        consumer_type2_reg(3) => consumer_type2_reg(3), 
        consumer_type2_reg(2) => consumer_type2_reg(2), 
        consumer_type2_reg(1) => consumer_type2_reg(1), 
        consumer_type2_reg(0) => consumer_type2_reg(0), 
        consumer_type4_reg(9) => consumer_type4_reg(9), 
        consumer_type4_reg(8) => consumer_type4_reg(8), 
        consumer_type4_reg(7) => consumer_type4_reg(7), 
        consumer_type4_reg(6) => consumer_type4_reg(6), 
        consumer_type4_reg(5) => consumer_type4_reg(5), 
        consumer_type4_reg(4) => consumer_type4_reg(4), 
        consumer_type4_reg(3) => consumer_type4_reg(3), 
        consumer_type4_reg(2) => consumer_type4_reg(2), 
        consumer_type4_reg(1) => consumer_type4_reg(1), 
        consumer_type4_reg(0) => consumer_type4_reg(0), 
        consumer_type3_reg(9) => consumer_type3_reg(9), 
        consumer_type3_reg(8) => consumer_type3_reg(8), 
        consumer_type3_reg(7) => consumer_type3_reg(7), 
        consumer_type3_reg(6) => consumer_type3_reg(6), 
        consumer_type3_reg(5) => consumer_type3_reg(5), 
        consumer_type3_reg(4) => consumer_type3_reg(4), 
        consumer_type3_reg(3) => consumer_type3_reg(3), 
        consumer_type3_reg(2) => consumer_type3_reg(2), 
        consumer_type3_reg(1) => consumer_type3_reg(1), 
        consumer_type3_reg(0) => consumer_type3_reg(0), 
        consumer_type1_reg(9) => consumer_type1_reg(9), 
        consumer_type1_reg(8) => consumer_type1_reg(8), 
        consumer_type1_reg(7) => consumer_type1_reg(7), 
        consumer_type1_reg(6) => consumer_type1_reg(6), 
        consumer_type1_reg(5) => consumer_type1_reg(5), 
        consumer_type1_reg(4) => consumer_type1_reg(4), 
        consumer_type1_reg(3) => consumer_type1_reg(3), 
        consumer_type1_reg(2) => consumer_type1_reg(2), 
        consumer_type1_reg(1) => consumer_type1_reg(1), 
        consumer_type1_reg(0) => consumer_type1_reg(0), 
        rx_crc_data_calc(11) => rx_crc_data_calc(11), 
        rx_crc_data_calc(10) => rx_crc_data_calc(10), 
        RX_FIFO_DIN(7) => \RX_FIFO_DIN[7]\, RX_FIFO_DIN(6) => 
        \RX_FIFO_DIN[6]\, RX_FIFO_DIN(5) => \RX_FIFO_DIN[5]\, 
        RX_FIFO_DIN(4) => \RX_FIFO_DIN[4]\, RX_FIFO_DIN(3) => 
        \RX_FIFO_DIN[3]\, RX_FIFO_DIN(2) => \RX_FIFO_DIN[2]\, 
        RX_FIFO_DIN(1) => \RX_FIFO_DIN[1]\, RX_FIFO_DIN(0) => 
        \RX_FIFO_DIN[0]\, RX_FIFO_DIN_pipe(8) => 
        RX_FIFO_DIN_pipe(8), RX_FIFO_DIN_pipe(7) => 
        RX_FIFO_DIN_pipe(7), RX_FIFO_DIN_pipe(6) => 
        RX_FIFO_DIN_pipe(6), RX_FIFO_DIN_pipe(5) => 
        RX_FIFO_DIN_pipe(5), RX_FIFO_DIN_pipe(4) => 
        RX_FIFO_DIN_pipe(4), RX_FIFO_DIN_pipe(3) => 
        RX_FIFO_DIN_pipe(3), RX_FIFO_DIN_pipe(2) => 
        RX_FIFO_DIN_pipe(2), RX_FIFO_DIN_pipe(1) => 
        RX_FIFO_DIN_pipe(1), RX_FIFO_DIN_pipe(0) => 
        RX_FIFO_DIN_pipe(0), lfsr_c_i_i_0 => lfsr_c_i_i_0, 
        DRVR_EN_c => DRVR_EN_c, clk1x_enable => clk1x_enable, 
        un2_apb3_reset => un2_apb3_reset, tx_col_detect_en => 
        tx_col_detect_en, packet_avail => packet_avail, 
        sampler_clk1x_en => \sampler_clk1x_en\, idle_line => 
        idle_line, RX_InProcess_d1 => RX_InProcess_d1, 
        rx_packet_complt => rx_packet_complt, N_535 => N_535, 
        RX_EarlyTerm => \RX_EarlyTerm\, SM_advance_i => 
        SM_advance_i, rx_crc_HighByte_en => rx_crc_HighByte_en, 
        iRX_FIFO_wr_en => iRX_FIFO_wr_en, N_41_i => N_41_i, 
        N_993_i => N_993_i, un2_apb3_reset_i => un2_apb3_reset_i, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, 
        rx_CRC_error_i => rx_CRC_error_i, rx_CRC_error => 
        rx_CRC_error);
    
    AFE_RX_STATE_MACHINE : AFE_RX_SM
      port map(RX_FIFO_DIN(7) => \RX_FIFO_DIN[7]\, RX_FIFO_DIN(6)
         => \RX_FIFO_DIN[6]\, RX_FIFO_DIN(5) => \RX_FIFO_DIN[5]\, 
        RX_FIFO_DIN(4) => \RX_FIFO_DIN[4]\, RX_FIFO_DIN(3) => 
        \RX_FIFO_DIN[3]\, RX_FIFO_DIN(2) => \RX_FIFO_DIN[2]\, 
        RX_FIFO_DIN(1) => \RX_FIFO_DIN[1]\, RX_FIFO_DIN(0) => 
        \RX_FIFO_DIN[0]\, manches_in_dly(1) => 
        \manches_in_dly[1]\, manches_in_dly(0) => 
        \manches_in_dly[0]\, irx_center_sample => 
        irx_center_sample, idle_line => idle_line, RX_EarlyTerm
         => \RX_EarlyTerm\, un2_apb3_reset => un2_apb3_reset, 
        clk1x_enable => clk1x_enable, packet_avail => 
        packet_avail, CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, 
        un2_apb3_reset_i => un2_apb3_reset_i, rx_packet_end_all
         => rx_packet_end_all);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_2Kx8_FIFO_2Kx8_0_LSRAM_top is

    port( fifo_MEMWADDR                : in    std_logic_vector(10 downto 0);
          CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0);
          fifo_MEMRADDR                : in    std_logic_vector(10 downto 0);
          RDATA_int                    : out   std_logic_vector(7 downto 0);
          fifo_MEMWE                   : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic;
          N_744_i                      : in    std_logic;
          BIT_CLK                      : in    std_logic
        );

end FIFO_2Kx8_FIFO_2Kx8_0_LSRAM_top;

architecture DEF_ARCH of FIFO_2Kx8_FIFO_2Kx8_0_LSRAM_top is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component RAM1K18
    generic (MEMORYFILE:string := "");

    port( A_DOUT        : out   std_logic_vector(17 downto 0);
          B_DOUT        : out   std_logic_vector(17 downto 0);
          BUSY          : out   std_logic;
          A_CLK         : in    std_logic := 'U';
          A_DOUT_CLK    : in    std_logic := 'U';
          A_ARST_N      : in    std_logic := 'U';
          A_DOUT_EN     : in    std_logic := 'U';
          A_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_DOUT_ARST_N : in    std_logic := 'U';
          A_DOUT_SRST_N : in    std_logic := 'U';
          A_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          A_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          A_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          B_CLK         : in    std_logic := 'U';
          B_DOUT_CLK    : in    std_logic := 'U';
          B_ARST_N      : in    std_logic := 'U';
          B_DOUT_EN     : in    std_logic := 'U';
          B_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_DOUT_ARST_N : in    std_logic := 'U';
          B_DOUT_SRST_N : in    std_logic := 'U';
          B_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          B_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          B_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          A_EN          : in    std_logic := 'U';
          A_DOUT_LAT    : in    std_logic := 'U';
          A_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_WMODE       : in    std_logic := 'U';
          B_EN          : in    std_logic := 'U';
          B_DOUT_LAT    : in    std_logic := 'U';
          B_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_WMODE       : in    std_logic := 'U';
          SII_LOCK      : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;
    signal nc24, nc1, nc8, nc13, nc16, nc19, nc25, nc20, nc27, 
        nc9, nc22, nc28, nc14, nc5, nc21, nc15, nc3, nc10, nc7, 
        nc17, nc4, nc12, nc2, nc23, nc18, nc26, nc6, nc11
         : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    FIFO_2Kx8_FIFO_2Kx8_0_LSRAM_top_R0C0 : RAM1K18
      port map(A_DOUT(17) => nc24, A_DOUT(16) => nc1, A_DOUT(15)
         => nc8, A_DOUT(14) => nc13, A_DOUT(13) => nc16, 
        A_DOUT(12) => nc19, A_DOUT(11) => nc25, A_DOUT(10) => 
        nc20, A_DOUT(9) => nc27, A_DOUT(8) => nc9, A_DOUT(7) => 
        RDATA_int(7), A_DOUT(6) => RDATA_int(6), A_DOUT(5) => 
        RDATA_int(5), A_DOUT(4) => RDATA_int(4), A_DOUT(3) => 
        RDATA_int(3), A_DOUT(2) => RDATA_int(2), A_DOUT(1) => 
        RDATA_int(1), A_DOUT(0) => RDATA_int(0), B_DOUT(17) => 
        nc22, B_DOUT(16) => nc28, B_DOUT(15) => nc14, B_DOUT(14)
         => nc5, B_DOUT(13) => nc21, B_DOUT(12) => nc15, 
        B_DOUT(11) => nc3, B_DOUT(10) => nc10, B_DOUT(9) => nc7, 
        B_DOUT(8) => nc17, B_DOUT(7) => nc4, B_DOUT(6) => nc12, 
        B_DOUT(5) => nc2, B_DOUT(4) => nc23, B_DOUT(3) => nc18, 
        B_DOUT(2) => nc26, B_DOUT(1) => nc6, B_DOUT(0) => nc11, 
        BUSY => OPEN, A_CLK => BIT_CLK, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_744_i, A_BLK(1) => VCC_net_1, A_BLK(0) => VCC_net_1, 
        A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => VCC_net_1, 
        A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, A_DIN(15)
         => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13) => 
        GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => GND_net_1, 
        A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, A_DIN(8)
         => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6) => 
        GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => GND_net_1, 
        A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, A_DIN(1)
         => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13) => 
        fifo_MEMRADDR(10), A_ADDR(12) => fifo_MEMRADDR(9), 
        A_ADDR(11) => fifo_MEMRADDR(8), A_ADDR(10) => 
        fifo_MEMRADDR(7), A_ADDR(9) => fifo_MEMRADDR(6), 
        A_ADDR(8) => fifo_MEMRADDR(5), A_ADDR(7) => 
        fifo_MEMRADDR(4), A_ADDR(6) => fifo_MEMRADDR(3), 
        A_ADDR(5) => fifo_MEMRADDR(2), A_ADDR(4) => 
        fifo_MEMRADDR(1), A_ADDR(3) => fifo_MEMRADDR(0), 
        A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, A_ADDR(0)
         => GND_net_1, A_WEN(1) => GND_net_1, A_WEN(0) => 
        GND_net_1, B_CLK => m2s010_som_sb_0_CCC_71MHz, B_DOUT_CLK
         => VCC_net_1, B_ARST_N => VCC_net_1, B_DOUT_EN => 
        VCC_net_1, B_BLK(2) => fifo_MEMWE, B_BLK(1) => VCC_net_1, 
        B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => GND_net_1, 
        B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => GND_net_1, 
        B_DIN(16) => GND_net_1, B_DIN(15) => GND_net_1, B_DIN(14)
         => GND_net_1, B_DIN(13) => GND_net_1, B_DIN(12) => 
        GND_net_1, B_DIN(11) => GND_net_1, B_DIN(10) => GND_net_1, 
        B_DIN(9) => GND_net_1, B_DIN(8) => GND_net_1, B_DIN(7)
         => CoreAPB3_0_APBmslave0_PWDATA(7), B_DIN(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), B_DIN(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), B_DIN(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), B_DIN(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), B_DIN(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), B_DIN(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), B_DIN(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), B_ADDR(13) => 
        fifo_MEMWADDR(10), B_ADDR(12) => fifo_MEMWADDR(9), 
        B_ADDR(11) => fifo_MEMWADDR(8), B_ADDR(10) => 
        fifo_MEMWADDR(7), B_ADDR(9) => fifo_MEMWADDR(6), 
        B_ADDR(8) => fifo_MEMWADDR(5), B_ADDR(7) => 
        fifo_MEMWADDR(4), B_ADDR(6) => fifo_MEMWADDR(3), 
        B_ADDR(5) => fifo_MEMWADDR(2), B_ADDR(4) => 
        fifo_MEMWADDR(1), B_ADDR(3) => fifo_MEMWADDR(0), 
        B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, B_ADDR(0)
         => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0) => 
        VCC_net_1, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_2Kx8_FIFO_2Kx8_0_ram_wrapper is

    port( RDATA_int                    : out   std_logic_vector(7 downto 0);
          fifo_MEMRADDR                : in    std_logic_vector(10 downto 0);
          CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0);
          fifo_MEMWADDR                : in    std_logic_vector(10 downto 0);
          BIT_CLK                      : in    std_logic;
          N_744_i                      : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic;
          fifo_MEMWE                   : in    std_logic
        );

end FIFO_2Kx8_FIFO_2Kx8_0_ram_wrapper;

architecture DEF_ARCH of FIFO_2Kx8_FIFO_2Kx8_0_ram_wrapper is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component FIFO_2Kx8_FIFO_2Kx8_0_LSRAM_top
    port( fifo_MEMWADDR                : in    std_logic_vector(10 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0) := (others => 'U');
          fifo_MEMRADDR                : in    std_logic_vector(10 downto 0) := (others => 'U');
          RDATA_int                    : out   std_logic_vector(7 downto 0);
          fifo_MEMWE                   : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic := 'U';
          N_744_i                      : in    std_logic := 'U';
          BIT_CLK                      : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : FIFO_2Kx8_FIFO_2Kx8_0_LSRAM_top
	Use entity work.FIFO_2Kx8_FIFO_2Kx8_0_LSRAM_top(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    L1_asyncnonpipe : FIFO_2Kx8_FIFO_2Kx8_0_LSRAM_top
      port map(fifo_MEMWADDR(10) => fifo_MEMWADDR(10), 
        fifo_MEMWADDR(9) => fifo_MEMWADDR(9), fifo_MEMWADDR(8)
         => fifo_MEMWADDR(8), fifo_MEMWADDR(7) => 
        fifo_MEMWADDR(7), fifo_MEMWADDR(6) => fifo_MEMWADDR(6), 
        fifo_MEMWADDR(5) => fifo_MEMWADDR(5), fifo_MEMWADDR(4)
         => fifo_MEMWADDR(4), fifo_MEMWADDR(3) => 
        fifo_MEMWADDR(3), fifo_MEMWADDR(2) => fifo_MEMWADDR(2), 
        fifo_MEMWADDR(1) => fifo_MEMWADDR(1), fifo_MEMWADDR(0)
         => fifo_MEMWADDR(0), CoreAPB3_0_APBmslave0_PWDATA(7) => 
        CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), fifo_MEMRADDR(10) => 
        fifo_MEMRADDR(10), fifo_MEMRADDR(9) => fifo_MEMRADDR(9), 
        fifo_MEMRADDR(8) => fifo_MEMRADDR(8), fifo_MEMRADDR(7)
         => fifo_MEMRADDR(7), fifo_MEMRADDR(6) => 
        fifo_MEMRADDR(6), fifo_MEMRADDR(5) => fifo_MEMRADDR(5), 
        fifo_MEMRADDR(4) => fifo_MEMRADDR(4), fifo_MEMRADDR(3)
         => fifo_MEMRADDR(3), fifo_MEMRADDR(2) => 
        fifo_MEMRADDR(2), fifo_MEMRADDR(1) => fifo_MEMRADDR(1), 
        fifo_MEMRADDR(0) => fifo_MEMRADDR(0), RDATA_int(7) => 
        RDATA_int(7), RDATA_int(6) => RDATA_int(6), RDATA_int(5)
         => RDATA_int(5), RDATA_int(4) => RDATA_int(4), 
        RDATA_int(3) => RDATA_int(3), RDATA_int(2) => 
        RDATA_int(2), RDATA_int(1) => RDATA_int(1), RDATA_int(0)
         => RDATA_int(0), fifo_MEMWE => fifo_MEMWE, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz, 
        N_744_i => N_744_i, BIT_CLK => BIT_CLK);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv_0 is

    port( wptr_bin_sync  : inout std_logic_vector(11 downto 0) := (others => 'Z');
          wptr_gray_sync : in    std_logic_vector(10 downto 0);
          bin_N_4_0_i    : out   std_logic
        );

end FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv_0;

architecture DEF_ARCH of 
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv_0 is 

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \bin_m3_0_3\, \bin_m3_0_2\, GND_net_1, VCC_net_1
         : std_logic;

begin 


    \bin_out_xhdl1_i_o2_RNIS01B2[10]\ : CFG3
      generic map(INIT => x"69")

      port map(A => \bin_m3_0_2\, B => \bin_m3_0_3\, C => 
        wptr_bin_sync(10), Y => bin_N_4_0_i);
    
    \bin_out_xhdl1_0_a2[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => wptr_bin_sync(2), B => wptr_gray_sync(1), Y
         => wptr_bin_sync(1));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \bin_out_xhdl1_0_a2[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => wptr_bin_sync(6), B => wptr_gray_sync(5), Y
         => wptr_bin_sync(5));
    
    \bin_out_xhdl1_0_a2[2]\ : CFG4
      generic map(INIT => x"9669")

      port map(A => \bin_m3_0_3\, B => wptr_bin_sync(10), C => 
        wptr_gray_sync(2), D => \bin_m3_0_2\, Y => 
        wptr_bin_sync(2));
    
    \bin_out_xhdl1_0_a2[0]\ : CFG3
      generic map(INIT => x"96")

      port map(A => wptr_gray_sync(1), B => wptr_bin_sync(2), C
         => wptr_gray_sync(0), Y => wptr_bin_sync(0));
    
    \bin_out_xhdl1_i_o2[9]\ : CFG3
      generic map(INIT => x"96")

      port map(A => wptr_gray_sync(9), B => wptr_bin_sync(11), C
         => wptr_gray_sync(10), Y => wptr_bin_sync(9));
    
    \bin_out_xhdl1_i_o2[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => wptr_bin_sync(11), B => wptr_gray_sync(10), Y
         => wptr_bin_sync(10));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \bin_out_xhdl1_0_a2[6]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(6), B => wptr_gray_sync(7), C
         => wptr_gray_sync(8), D => wptr_bin_sync(9), Y => 
        wptr_bin_sync(6));
    
    \bin_out_xhdl1_0_a2[4]\ : CFG3
      generic map(INIT => x"96")

      port map(A => wptr_gray_sync(4), B => wptr_gray_sync(5), C
         => wptr_bin_sync(6), Y => wptr_bin_sync(4));
    
    bin_m3_0_2 : CFG3
      generic map(INIT => x"96")

      port map(A => wptr_gray_sync(3), B => wptr_gray_sync(4), C
         => wptr_gray_sync(5), Y => \bin_m3_0_2\);
    
    \bin_out_xhdl1_0_a2[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => wptr_bin_sync(9), B => wptr_gray_sync(8), Y
         => wptr_bin_sync(8));
    
    bin_m3_0_3 : CFG4
      generic map(INIT => x"9669")

      port map(A => wptr_gray_sync(7), B => wptr_gray_sync(8), C
         => wptr_gray_sync(9), D => wptr_gray_sync(6), Y => 
        \bin_m3_0_3\);
    
    \bin_out_xhdl1_0_a2[7]\ : CFG3
      generic map(INIT => x"96")

      port map(A => wptr_gray_sync(8), B => wptr_bin_sync(9), C
         => wptr_gray_sync(7), Y => wptr_bin_sync(7));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_1 is

    port( wptr_gray       : in    std_logic_vector(11 downto 0);
          wptr_gray_sync  : out   std_logic_vector(10 downto 0);
          wptr_bin_sync_0 : out   std_logic;
          BIT_CLK         : in    std_logic;
          itx_fifo_rst_i  : in    std_logic
        );

end FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_1;

architecture DEF_ARCH of 
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_1 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \sync_int[10]_net_1\, VCC_net_1, GND_net_1, 
        \sync_int[11]_net_1\, \sync_int[0]_net_1\, 
        \sync_int[1]_net_1\, \sync_int[2]_net_1\, 
        \sync_int[3]_net_1\, \sync_int[4]_net_1\, 
        \sync_int[5]_net_1\, \sync_int[6]_net_1\, 
        \sync_int[7]_net_1\, \sync_int[8]_net_1\, 
        \sync_int[9]_net_1\ : std_logic;

begin 


    \sync_int[9]\ : SLE
      port map(D => wptr_gray(9), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[9]_net_1\);
    
    \sync_int[4]\ : SLE
      port map(D => wptr_gray(4), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[4]_net_1\);
    
    \sync_out_xhdl1[10]\ : SLE
      port map(D => \sync_int[10]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(10));
    
    \sync_int[1]\ : SLE
      port map(D => wptr_gray(1), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[1]_net_1\);
    
    \sync_int[11]\ : SLE
      port map(D => wptr_gray(11), CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[11]_net_1\);
    
    \sync_out_xhdl1[6]\ : SLE
      port map(D => \sync_int[6]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(6));
    
    \sync_out_xhdl1[3]\ : SLE
      port map(D => \sync_int[3]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(3));
    
    \sync_int[6]\ : SLE
      port map(D => wptr_gray(6), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[6]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \sync_out_xhdl1[11]\ : SLE
      port map(D => \sync_int[11]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_bin_sync_0);
    
    \sync_int[3]\ : SLE
      port map(D => wptr_gray(3), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[3]_net_1\);
    
    \sync_out_xhdl1[4]\ : SLE
      port map(D => \sync_int[4]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(4));
    
    \sync_int[0]\ : SLE
      port map(D => wptr_gray(0), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[0]_net_1\);
    
    \sync_out_xhdl1[1]\ : SLE
      port map(D => \sync_int[1]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(1));
    
    \sync_int[5]\ : SLE
      port map(D => wptr_gray(5), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[5]_net_1\);
    
    \sync_int[2]\ : SLE
      port map(D => wptr_gray(2), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[2]_net_1\);
    
    \sync_out_xhdl1[9]\ : SLE
      port map(D => \sync_int[9]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(9));
    
    \sync_out_xhdl1[2]\ : SLE
      port map(D => \sync_int[2]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(2));
    
    \sync_int[8]\ : SLE
      port map(D => wptr_gray(8), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[8]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sync_out_xhdl1[7]\ : SLE
      port map(D => \sync_int[7]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(7));
    
    \sync_out_xhdl1[5]\ : SLE
      port map(D => \sync_int[5]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(5));
    
    \sync_out_xhdl1[0]\ : SLE
      port map(D => \sync_int[0]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(0));
    
    \sync_out_xhdl1[8]\ : SLE
      port map(D => \sync_int[8]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(8));
    
    \sync_int[7]\ : SLE
      port map(D => wptr_gray(7), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[7]_net_1\);
    
    \sync_int[10]\ : SLE
      port map(D => wptr_gray(10), CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_0 is

    port( rptr_gray                 : in    std_logic_vector(11 downto 0);
          rptr_gray_sync            : out   std_logic_vector(10 downto 0);
          rptr_bin_sync_0           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          itx_fifo_rst_i            : in    std_logic
        );

end FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_0;

architecture DEF_ARCH of 
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_0 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \sync_int[4]_net_1\, GND_net_1, 
        \sync_int[5]_net_1\, \sync_int[6]_net_1\, 
        \sync_int[7]_net_1\, \sync_int[8]_net_1\, 
        \sync_int[9]_net_1\, \sync_int[10]_net_1\, 
        \sync_int[11]_net_1\, \sync_int[1]_net_1\, 
        \sync_int[2]_net_1\, \sync_int[3]_net_1\, 
        \sync_int[0]_net_1\ : std_logic;

begin 


    \sync_int[9]\ : SLE
      port map(D => rptr_gray(9), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[9]_net_1\);
    
    \sync_int[4]\ : SLE
      port map(D => rptr_gray(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[4]_net_1\);
    
    \sync_out_xhdl1[10]\ : SLE
      port map(D => \sync_int[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(10));
    
    \sync_int[1]\ : SLE
      port map(D => rptr_gray(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[1]_net_1\);
    
    \sync_int[11]\ : SLE
      port map(D => rptr_gray(11), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[11]_net_1\);
    
    \sync_out_xhdl1[6]\ : SLE
      port map(D => \sync_int[6]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(6));
    
    \sync_out_xhdl1[3]\ : SLE
      port map(D => \sync_int[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(3));
    
    \sync_int[6]\ : SLE
      port map(D => rptr_gray(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[6]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \sync_out_xhdl1[11]\ : SLE
      port map(D => \sync_int[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_bin_sync_0);
    
    \sync_int[3]\ : SLE
      port map(D => rptr_gray(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[3]_net_1\);
    
    \sync_out_xhdl1[4]\ : SLE
      port map(D => \sync_int[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(4));
    
    \sync_int[0]\ : SLE
      port map(D => rptr_gray(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[0]_net_1\);
    
    \sync_out_xhdl1[1]\ : SLE
      port map(D => \sync_int[1]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(1));
    
    \sync_int[5]\ : SLE
      port map(D => rptr_gray(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[5]_net_1\);
    
    \sync_int[2]\ : SLE
      port map(D => rptr_gray(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[2]_net_1\);
    
    \sync_out_xhdl1[9]\ : SLE
      port map(D => \sync_int[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(9));
    
    \sync_out_xhdl1[2]\ : SLE
      port map(D => \sync_int[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(2));
    
    \sync_int[8]\ : SLE
      port map(D => rptr_gray(8), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[8]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sync_out_xhdl1[7]\ : SLE
      port map(D => \sync_int[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(7));
    
    \sync_out_xhdl1[5]\ : SLE
      port map(D => \sync_int[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(5));
    
    \sync_out_xhdl1[0]\ : SLE
      port map(D => \sync_int[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(0));
    
    \sync_out_xhdl1[8]\ : SLE
      port map(D => \sync_int[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(8));
    
    \sync_int[7]\ : SLE
      port map(D => rptr_gray(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[7]_net_1\);
    
    \sync_int[10]\ : SLE
      port map(D => rptr_gray(10), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv is

    port( rptr_bin_sync  : inout std_logic_vector(11 downto 0) := (others => 'Z');
          rptr_gray_sync : in    std_logic_vector(10 downto 0)
        );

end FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv;

architecture DEF_ARCH of 
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    \bin_out_xhdl1_0_a2[1]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(3), B => rptr_gray_sync(1), C
         => rptr_bin_sync(4), D => rptr_gray_sync(2), Y => 
        rptr_bin_sync(1));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \bin_out_xhdl1_0_a2[5]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(7), B => rptr_gray_sync(6), C
         => rptr_gray_sync(5), D => rptr_bin_sync(8), Y => 
        rptr_bin_sync(5));
    
    \bin_out_xhdl1_0_a2[2]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(4), B => rptr_gray_sync(3), C
         => rptr_gray_sync(2), D => rptr_bin_sync(5), Y => 
        rptr_bin_sync(2));
    
    \bin_out_xhdl1_0_a2[0]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(2), B => rptr_bin_sync(3), C
         => rptr_gray_sync(0), D => rptr_gray_sync(1), Y => 
        rptr_bin_sync(0));
    
    \bin_out_xhdl1_i_o2[9]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(10), B => rptr_gray_sync(9), C
         => rptr_bin_sync(11), Y => rptr_bin_sync(9));
    
    \bin_out_xhdl1_i_o2[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(11), B => rptr_gray_sync(10), Y
         => rptr_bin_sync(10));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \bin_out_xhdl1_0_a2[6]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(8), B => rptr_gray_sync(7), C
         => rptr_gray_sync(6), D => rptr_bin_sync(9), Y => 
        rptr_bin_sync(6));
    
    \bin_out_xhdl1_0_a2[4]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(6), B => rptr_gray_sync(5), C
         => rptr_gray_sync(4), D => rptr_bin_sync(7), Y => 
        rptr_bin_sync(4));
    
    \bin_out_xhdl1_0_a2[8]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(10), B => rptr_gray_sync(9), C
         => rptr_gray_sync(8), D => rptr_bin_sync(11), Y => 
        rptr_bin_sync(8));
    
    \bin_out_xhdl1_0_a2[7]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(9), B => rptr_gray_sync(8), C
         => rptr_gray_sync(7), D => rptr_bin_sync(10), Y => 
        rptr_bin_sync(7));
    
    \bin_out_xhdl1_0_a2[3]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(5), B => rptr_gray_sync(4), C
         => rptr_gray_sync(3), D => rptr_bin_sync(6), Y => 
        rptr_bin_sync(3));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_2Kx8_FIFO_2Kx8_0_corefifo_async is

    port( fifo_MEMWADDR                   : out   std_logic_vector(10 downto 0);
          fifo_MEMRADDR                   : out   std_logic_vector(10 downto 0);
          N_432_i                         : out   std_logic;
          byte_clk_en                     : in    std_logic;
          TX_PreAmble                     : in    std_logic;
          un1_tx_packet_length_0_sqmuxa_o : in    std_logic;
          TX_DataEn_1_o                   : in    std_logic;
          TX_FIFO_wr_en                   : in    std_logic;
          fifo_MEMWE                      : out   std_logic;
          N_744_i                         : out   std_logic;
          TX_FIFO_Full                    : out   std_logic;
          TX_FIFO_Empty                   : out   std_logic;
          BIT_CLK                         : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz       : in    std_logic;
          itx_fifo_rst_i                  : in    std_logic;
          TX_FIFO_OVERFLOW_i              : out   std_logic;
          TX_FIFO_OVERFLOW                : out   std_logic;
          TX_FIFO_UNDERRUN_i              : out   std_logic;
          TX_FIFO_UNDERRUN                : out   std_logic
        );

end FIFO_2Kx8_FIFO_2Kx8_0_corefifo_async;

architecture DEF_ARCH of FIFO_2Kx8_FIFO_2Kx8_0_corefifo_async is 

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv_0
    port( wptr_bin_sync  : inout   std_logic_vector(11 downto 0);
          wptr_gray_sync : in    std_logic_vector(10 downto 0) := (others => 'U');
          bin_N_4_0_i    : out   std_logic
        );
  end component;

  component FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_1
    port( wptr_gray       : in    std_logic_vector(11 downto 0) := (others => 'U');
          wptr_gray_sync  : out   std_logic_vector(10 downto 0);
          wptr_bin_sync_0 : out   std_logic;
          BIT_CLK         : in    std_logic := 'U';
          itx_fifo_rst_i  : in    std_logic := 'U'
        );
  end component;

  component FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_0
    port( rptr_gray                 : in    std_logic_vector(11 downto 0) := (others => 'U');
          rptr_gray_sync            : out   std_logic_vector(10 downto 0);
          rptr_bin_sync_0           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          itx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv
    port( rptr_bin_sync  : inout   std_logic_vector(11 downto 0);
          rptr_gray_sync : in    std_logic_vector(10 downto 0) := (others => 'U')
        );
  end component;

    signal \wptr[0]_net_1\, \wptr_s[0]\, \fifo_MEMWADDR[0]\, 
        \memwaddr_r_s[0]\, \fifo_MEMRADDR[0]\, \memraddr_r_s[0]\, 
        \rptr[0]_net_1\, \rptr_s[0]\, \TX_FIFO_UNDERRUN\, 
        \TX_FIFO_OVERFLOW\, \wptr_gray[10]_net_1\, VCC_net_1, 
        \wptr_gray_1[10]_net_1\, GND_net_1, \wptr_gray[11]_net_1\, 
        \wptr[11]_net_1\, \rptr_gray[0]_net_1\, 
        \rptr_gray_1[0]_net_1\, \rptr_gray[1]_net_1\, 
        \rptr_gray_1[1]_net_1\, \rptr_gray[2]_net_1\, 
        \rptr_gray_1[2]_net_1\, \rptr_gray[3]_net_1\, 
        \rptr_gray_1[3]_net_1\, \rptr_gray[4]_net_1\, 
        \rptr_gray_1[4]_net_1\, \rptr_gray[5]_net_1\, 
        \rptr_gray_1[5]_net_1\, \rptr_gray[6]_net_1\, 
        \rptr_gray_1[6]_net_1\, \rptr_gray[7]_net_1\, 
        \rptr_gray_1[7]_net_1\, \rptr_gray[8]_net_1\, 
        \rptr_gray_1[8]_net_1\, \rptr_gray[9]_net_1\, 
        \rptr_gray_1[9]_net_1\, \rptr_gray[10]_net_1\, 
        \rptr_gray_1[10]_net_1\, \rptr_gray[11]_net_1\, 
        \rptr[11]_net_1\, \rptr_bin_sync2[7]_net_1\, 
        \rptr_bin_sync[7]\, \rptr_bin_sync2[8]_net_1\, 
        \rptr_bin_sync[8]\, \rptr_bin_sync2[9]_net_1\, 
        \rptr_bin_sync[9]\, \rptr_bin_sync2[10]_net_1\, 
        \rptr_bin_sync[10]\, \rptr_bin_sync2[11]_net_1\, 
        \rptr_bin_sync[11]\, \wptr_gray[0]_net_1\, 
        \wptr_gray_1[0]_net_1\, \wptr_gray[1]_net_1\, 
        \wptr_gray_1[1]_net_1\, \wptr_gray[2]_net_1\, 
        \wptr_gray_1[2]_net_1\, \wptr_gray[3]_net_1\, 
        \wptr_gray_1[3]_net_1\, \wptr_gray[4]_net_1\, 
        \wptr_gray_1[4]_net_1\, \wptr_gray[5]_net_1\, 
        \wptr_gray_1[5]_net_1\, \wptr_gray[6]_net_1\, 
        \wptr_gray_1[6]_net_1\, \wptr_gray[7]_net_1\, 
        \wptr_gray_1[7]_net_1\, \wptr_gray[8]_net_1\, 
        \wptr_gray_1[8]_net_1\, \wptr_gray[9]_net_1\, 
        \wptr_gray_1[9]_net_1\, \rptr_bin_sync2[0]_net_1\, 
        \rptr_bin_sync[0]\, \rptr_bin_sync2[1]_net_1\, 
        \rptr_bin_sync[1]\, \rptr_bin_sync2[2]_net_1\, 
        \rptr_bin_sync[2]\, \rptr_bin_sync2[3]_net_1\, 
        \rptr_bin_sync[3]\, \rptr_bin_sync2[4]_net_1\, 
        \rptr_bin_sync[4]\, \rptr_bin_sync2[5]_net_1\, 
        \rptr_bin_sync[5]\, \rptr_bin_sync2[6]_net_1\, 
        \rptr_bin_sync[6]\, \wptr_bin_sync2[7]_net_1\, 
        \wptr_bin_sync[7]\, \wptr_bin_sync2[8]_net_1\, 
        \wptr_bin_sync[8]\, \wptr_bin_sync2[9]_net_1\, 
        \wptr_bin_sync[9]\, \wptr_bin_sync2[10]_net_1\, 
        \wptr_bin_sync[10]\, \wptr_bin_sync2[11]_net_1\, 
        \wptr_bin_sync[11]\, N_416_i, rdiff_bus, 
        \wptr_bin_sync[0]\, \wptr_bin_sync2[1]_net_1\, 
        \wptr_bin_sync[1]\, \wptr_bin_sync2[2]_net_1\, 
        \wptr_bin_sync[2]\, \wptr_bin_sync2[3]_net_1\, 
        bin_N_4_0_i, \wptr_bin_sync2[4]_net_1\, 
        \wptr_bin_sync[4]\, \wptr_bin_sync2[5]_net_1\, 
        \wptr_bin_sync[5]\, \wptr_bin_sync2[6]_net_1\, 
        \wptr_bin_sync[6]\, \TX_FIFO_Empty\, empty_r_3, N_1349_i, 
        \TX_FIFO_Full\, \fulli\, \N_744_i\, \rptr[1]_net_1\, 
        \rptr_s[1]\, \rptr[2]_net_1\, \rptr_s[2]\, 
        \rptr[3]_net_1\, \rptr_s[3]\, \rptr[4]_net_1\, 
        \rptr_s[4]\, \rptr[5]_net_1\, \rptr_s[5]\, 
        \rptr[6]_net_1\, \rptr_s[6]\, \rptr[7]_net_1\, 
        \rptr_s[7]\, \rptr[8]_net_1\, \rptr_s[8]\, 
        \rptr[9]_net_1\, \rptr_s[9]\, \rptr[10]_net_1\, 
        \rptr_s[10]\, \rptr_s[11]_net_1\, \fifo_MEMRADDR[1]\, 
        \memraddr_r_s[1]\, \fifo_MEMRADDR[2]\, \memraddr_r_s[2]\, 
        \fifo_MEMRADDR[3]\, \memraddr_r_s[3]\, \fifo_MEMRADDR[4]\, 
        \memraddr_r_s[4]\, \fifo_MEMRADDR[5]\, \memraddr_r_s[5]\, 
        \fifo_MEMRADDR[6]\, \memraddr_r_s[6]\, \fifo_MEMRADDR[7]\, 
        \memraddr_r_s[7]\, \fifo_MEMRADDR[8]\, \memraddr_r_s[8]\, 
        \fifo_MEMRADDR[9]\, \memraddr_r_s[9]\, 
        \fifo_MEMRADDR[10]\, \memraddr_r_s[10]_net_1\, 
        \fifo_MEMWE\, \fifo_MEMWADDR[1]\, \memwaddr_r_s[1]\, 
        \fifo_MEMWADDR[2]\, \memwaddr_r_s[2]\, \fifo_MEMWADDR[3]\, 
        \memwaddr_r_s[3]\, \fifo_MEMWADDR[4]\, \memwaddr_r_s[4]\, 
        \fifo_MEMWADDR[5]\, \memwaddr_r_s[5]\, \fifo_MEMWADDR[6]\, 
        \memwaddr_r_s[6]\, \fifo_MEMWADDR[7]\, \memwaddr_r_s[7]\, 
        \fifo_MEMWADDR[8]\, \memwaddr_r_s[8]\, \fifo_MEMWADDR[9]\, 
        \memwaddr_r_s[9]\, \fifo_MEMWADDR[10]\, 
        \memwaddr_r_s[10]_net_1\, \wptr[1]_net_1\, \wptr_s[1]\, 
        \wptr[2]_net_1\, \wptr_s[2]\, \wptr[3]_net_1\, 
        \wptr_s[3]\, \wptr[4]_net_1\, \wptr_s[4]\, 
        \wptr[5]_net_1\, \wptr_s[5]\, \wptr[6]_net_1\, 
        \wptr_s[6]\, \wptr[7]_net_1\, \wptr_s[7]\, 
        \wptr[8]_net_1\, \wptr_s[8]\, \wptr[9]_net_1\, 
        \wptr_s[9]\, \wptr[10]_net_1\, \wptr_s[10]\, 
        \wptr_s[11]_net_1\, \wdiff_bus_cry_0\, wdiff_bus_cry_0_Y, 
        \wdiff_bus_cry_1\, \wdiff_bus[1]\, \wdiff_bus_cry_2\, 
        \wdiff_bus[2]\, \wdiff_bus_cry_3\, \wdiff_bus[3]\, 
        \wdiff_bus_cry_4\, \wdiff_bus[4]\, \wdiff_bus_cry_5\, 
        \wdiff_bus[5]\, \wdiff_bus_cry_6\, \wdiff_bus[6]\, 
        \wdiff_bus_cry_7\, \wdiff_bus[7]\, \wdiff_bus_cry_8\, 
        \wdiff_bus[8]\, \wdiff_bus_cry_9\, \wdiff_bus[9]\, 
        \wdiff_bus[11]\, \wdiff_bus_cry_10\, \wdiff_bus[10]\, 
        \rdiff_bus_cry_0\, rdiff_bus_cry_0_Y, \rdiff_bus_cry_1\, 
        \rdiff_bus[1]\, \rdiff_bus_cry_2\, \rdiff_bus[2]\, 
        \rdiff_bus_cry_3\, \rdiff_bus[3]\, \rdiff_bus_cry_4\, 
        \rdiff_bus[4]\, \rdiff_bus_cry_5\, \rdiff_bus[5]\, 
        \rdiff_bus_cry_6\, \rdiff_bus[6]\, \rdiff_bus_cry_7\, 
        \rdiff_bus[7]\, \rdiff_bus_cry_8\, \rdiff_bus[8]\, 
        \rdiff_bus_cry_9\, \rdiff_bus[9]\, \rdiff_bus[11]\, 
        \rdiff_bus_cry_10\, \rdiff_bus[10]\, wptr_s_386_FCO, 
        \wptr_cry[1]_net_1\, \wptr_cry[2]_net_1\, 
        \wptr_cry[3]_net_1\, \wptr_cry[4]_net_1\, 
        \wptr_cry[5]_net_1\, \wptr_cry[6]_net_1\, 
        \wptr_cry[7]_net_1\, \wptr_cry[8]_net_1\, 
        \wptr_cry[9]_net_1\, \wptr_cry[10]_net_1\, 
        memwaddr_r_s_387_FCO, \memwaddr_r_cry[1]_net_1\, 
        \memwaddr_r_cry[2]_net_1\, \memwaddr_r_cry[3]_net_1\, 
        \memwaddr_r_cry[4]_net_1\, \memwaddr_r_cry[5]_net_1\, 
        \memwaddr_r_cry[6]_net_1\, \memwaddr_r_cry[7]_net_1\, 
        \memwaddr_r_cry[8]_net_1\, \memwaddr_r_cry[9]_net_1\, 
        memraddr_r_s_388_FCO, \memraddr_r_cry[1]_net_1\, 
        \memraddr_r_cry[2]_net_1\, \memraddr_r_cry[3]_net_1\, 
        \memraddr_r_cry[4]_net_1\, \memraddr_r_cry[5]_net_1\, 
        \memraddr_r_cry[6]_net_1\, \memraddr_r_cry[7]_net_1\, 
        \memraddr_r_cry[8]_net_1\, \memraddr_r_cry[9]_net_1\, 
        rptr_s_389_FCO, \rptr_cry[1]_net_1\, \rptr_cry[2]_net_1\, 
        \rptr_cry[3]_net_1\, \rptr_cry[4]_net_1\, 
        \rptr_cry[5]_net_1\, \rptr_cry[6]_net_1\, 
        \rptr_cry[7]_net_1\, \rptr_cry[8]_net_1\, 
        \rptr_cry[9]_net_1\, \rptr_cry[10]_net_1\, 
        empty_r_3_0_a2_7, empty_r_3_0_a2_6, un4_fullilto10_i_a2_7, 
        un4_fullilto10_i_a2_6, empty_r_3_0_a2_8, \N_432_i\, 
        un4_fullilto10_i_a2_8, \wptr_gray_sync[0]\, 
        \wptr_gray_sync[1]\, \wptr_gray_sync[2]\, 
        \wptr_gray_sync[3]\, \wptr_gray_sync[4]\, 
        \wptr_gray_sync[5]\, \wptr_gray_sync[6]\, 
        \wptr_gray_sync[7]\, \wptr_gray_sync[8]\, 
        \wptr_gray_sync[9]\, \wptr_gray_sync[10]\, 
        \rptr_gray_sync[0]\, \rptr_gray_sync[1]\, 
        \rptr_gray_sync[2]\, \rptr_gray_sync[3]\, 
        \rptr_gray_sync[4]\, \rptr_gray_sync[5]\, 
        \rptr_gray_sync[6]\, \rptr_gray_sync[7]\, 
        \rptr_gray_sync[8]\, \rptr_gray_sync[9]\, 
        \rptr_gray_sync[10]\ : std_logic;
    signal nc1 : std_logic;

    for all : FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv_0
	Use entity work.
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv_0(DEF_ARCH);
    for all : FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_1
	Use entity work.
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_1(DEF_ARCH);
    for all : FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_0
	Use entity work.
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_0(DEF_ARCH);
    for all : FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv
	Use entity work.
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv(DEF_ARCH);
begin 

    fifo_MEMWADDR(10) <= \fifo_MEMWADDR[10]\;
    fifo_MEMWADDR(9) <= \fifo_MEMWADDR[9]\;
    fifo_MEMWADDR(8) <= \fifo_MEMWADDR[8]\;
    fifo_MEMWADDR(7) <= \fifo_MEMWADDR[7]\;
    fifo_MEMWADDR(6) <= \fifo_MEMWADDR[6]\;
    fifo_MEMWADDR(5) <= \fifo_MEMWADDR[5]\;
    fifo_MEMWADDR(4) <= \fifo_MEMWADDR[4]\;
    fifo_MEMWADDR(3) <= \fifo_MEMWADDR[3]\;
    fifo_MEMWADDR(2) <= \fifo_MEMWADDR[2]\;
    fifo_MEMWADDR(1) <= \fifo_MEMWADDR[1]\;
    fifo_MEMWADDR(0) <= \fifo_MEMWADDR[0]\;
    fifo_MEMRADDR(10) <= \fifo_MEMRADDR[10]\;
    fifo_MEMRADDR(9) <= \fifo_MEMRADDR[9]\;
    fifo_MEMRADDR(8) <= \fifo_MEMRADDR[8]\;
    fifo_MEMRADDR(7) <= \fifo_MEMRADDR[7]\;
    fifo_MEMRADDR(6) <= \fifo_MEMRADDR[6]\;
    fifo_MEMRADDR(5) <= \fifo_MEMRADDR[5]\;
    fifo_MEMRADDR(4) <= \fifo_MEMRADDR[4]\;
    fifo_MEMRADDR(3) <= \fifo_MEMRADDR[3]\;
    fifo_MEMRADDR(2) <= \fifo_MEMRADDR[2]\;
    fifo_MEMRADDR(1) <= \fifo_MEMRADDR[1]\;
    fifo_MEMRADDR(0) <= \fifo_MEMRADDR[0]\;
    N_432_i <= \N_432_i\;
    fifo_MEMWE <= \fifo_MEMWE\;
    N_744_i <= \N_744_i\;
    TX_FIFO_Full <= \TX_FIFO_Full\;
    TX_FIFO_Empty <= \TX_FIFO_Empty\;
    TX_FIFO_OVERFLOW <= \TX_FIFO_OVERFLOW\;
    TX_FIFO_UNDERRUN <= \TX_FIFO_UNDERRUN\;

    \rptr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[4]_net_1\, S
         => \rptr_s[5]\, Y => OPEN, FCO => \rptr_cry[5]_net_1\);
    
    underflow_r_RNIFFTA : CFG1
      generic map(INIT => "01")

      port map(A => \TX_FIFO_UNDERRUN\, Y => TX_FIFO_UNDERRUN_i);
    
    wdiff_bus_cry_8 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[8]_net_1\, B => 
        \rptr_bin_sync2[8]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_7\, S => \wdiff_bus[8]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_8\);
    
    wptr_s_386 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => wptr_s_386_FCO);
    
    \wptr_gray[4]\ : SLE
      port map(D => \wptr_gray_1[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[4]_net_1\);
    
    \rptr_gray_1[3]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[3]_net_1\, B => \rptr[4]_net_1\, Y => 
        \rptr_gray_1[3]_net_1\);
    
    \rptr_bin_sync2[6]\ : SLE
      port map(D => \rptr_bin_sync[6]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[6]_net_1\);
    
    \rptr[1]\ : SLE
      port map(D => \rptr_s[1]\, CLK => BIT_CLK, EN => \N_744_i\, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[1]_net_1\);
    
    \wptr_gray_1[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[9]_net_1\, B => \wptr[10]_net_1\, Y => 
        \wptr_gray_1[9]_net_1\);
    
    \rptr_gray_1[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[5]_net_1\, B => \rptr[6]_net_1\, Y => 
        \rptr_gray_1[5]_net_1\);
    
    \rptr_gray[9]\ : SLE
      port map(D => \rptr_gray_1[9]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[9]_net_1\);
    
    \rptr_gray[8]\ : SLE
      port map(D => \rptr_gray_1[8]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[8]_net_1\);
    
    \rptr_gray_1[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[2]_net_1\, B => \rptr[3]_net_1\, Y => 
        \rptr_gray_1[2]_net_1\);
    
    \rptr_bin_sync2[7]\ : SLE
      port map(D => \rptr_bin_sync[7]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[7]_net_1\);
    
    \memwaddr_r[1]\ : SLE
      port map(D => \memwaddr_r_s[1]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[1]\);
    
    fulli : CFG4
      generic map(INIT => x"EAAA")

      port map(A => \wdiff_bus[11]\, B => TX_FIFO_wr_en, C => 
        un4_fullilto10_i_a2_8, D => un4_fullilto10_i_a2_7, Y => 
        \fulli\);
    
    \memwaddr_r_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[5]_net_1\, S => \memwaddr_r_s[6]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[6]_net_1\);
    
    \memwaddr_r_s[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[9]_net_1\, S => \memwaddr_r_s[10]_net_1\, 
        Y => OPEN, FCO => OPEN);
    
    \wptr_gray_1[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[7]_net_1\, B => \wptr[8]_net_1\, Y => 
        \wptr_gray_1[7]_net_1\);
    
    \memraddr_r[0]\ : SLE
      port map(D => \memraddr_r_s[0]\, CLK => BIT_CLK, EN => 
        \N_744_i\, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[0]\);
    
    \wptr[0]\ : SLE
      port map(D => \wptr_s[0]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[0]_net_1\);
    
    \rptr_bin_sync2[8]\ : SLE
      port map(D => \rptr_bin_sync[8]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[8]_net_1\);
    
    \rptr_gray_1[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[1]_net_1\, B => \rptr[2]_net_1\, Y => 
        \rptr_gray_1[1]_net_1\);
    
    \rptr_gray[10]\ : SLE
      port map(D => \rptr_gray_1[10]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[10]_net_1\);
    
    \wptr_gray_1[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[0]_net_1\, B => \wptr[1]_net_1\, Y => 
        \wptr_gray_1[0]_net_1\);
    
    wdiff_bus_cry_9 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[9]_net_1\, B => 
        \rptr_bin_sync2[9]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_8\, S => \wdiff_bus[9]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_9\);
    
    \rptr[5]\ : SLE
      port map(D => \rptr_s[5]\, CLK => BIT_CLK, EN => \N_744_i\, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[5]_net_1\);
    
    \rptr_gray[3]\ : SLE
      port map(D => \rptr_gray_1[3]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[3]_net_1\);
    
    \rptr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[5]_net_1\, S
         => \rptr_s[6]\, Y => OPEN, FCO => \rptr_cry[6]_net_1\);
    
    \memwaddr_r_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[1]\, C => 
        GND_net_1, D => GND_net_1, FCI => memwaddr_r_s_387_FCO, S
         => \memwaddr_r_s[1]\, Y => OPEN, FCO => 
        \memwaddr_r_cry[1]_net_1\);
    
    \wptr_gray[3]\ : SLE
      port map(D => \wptr_gray_1[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[3]_net_1\);
    
    \rptr_gray_1[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[11]_net_1\, B => \rptr[10]_net_1\, Y
         => \rptr_gray_1[10]_net_1\);
    
    wdiff_bus_s_11 : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \rptr_bin_sync2[11]_net_1\, C
         => \wptr[11]_net_1\, D => GND_net_1, FCI => 
        \wdiff_bus_cry_10\, S => \wdiff_bus[11]\, Y => OPEN, FCO
         => OPEN);
    
    \rptr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[7]_net_1\, S
         => \rptr_s[8]\, Y => OPEN, FCO => \rptr_cry[8]_net_1\);
    
    \rptr[7]\ : SLE
      port map(D => \rptr_s[7]\, CLK => BIT_CLK, EN => \N_744_i\, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[7]_net_1\);
    
    rdiff_bus_cry_4 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[4]_net_1\, B => 
        \rptr[4]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_3\, S => \rdiff_bus[4]\, Y => OPEN, FCO
         => \rdiff_bus_cry_4\);
    
    \rptr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[9]_net_1\, S
         => \rptr_s[10]\, Y => OPEN, FCO => \rptr_cry[10]_net_1\);
    
    \rptr_bin_sync2[0]\ : SLE
      port map(D => \rptr_bin_sync[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[0]_net_1\);
    
    \L1.empty_r_3_0_a2_7\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \rdiff_bus[7]\, B => \rdiff_bus[8]\, C => 
        \rdiff_bus[9]\, D => \rdiff_bus[10]\, Y => 
        empty_r_3_0_a2_7);
    
    \wptr[11]\ : SLE
      port map(D => \wptr_s[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \wptr[11]_net_1\);
    
    rptr_s_389 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => rptr_s_389_FCO);
    
    rdiff_bus_cry_1 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[1]_net_1\, B => 
        \rptr[1]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_0\, S => \rdiff_bus[1]\, Y => OPEN, FCO
         => \rdiff_bus_cry_1\);
    
    \memraddr_r[1]\ : SLE
      port map(D => \memraddr_r_s[1]\, CLK => BIT_CLK, EN => 
        \N_744_i\, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[1]\);
    
    \rptr_bin_sync2[2]\ : SLE
      port map(D => \rptr_bin_sync[2]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[2]_net_1\);
    
    rdiff_bus_cry_6 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[6]_net_1\, B => 
        \rptr[6]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_5\, S => \rdiff_bus[6]\, Y => OPEN, FCO
         => \rdiff_bus_cry_6\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \memwaddr_r_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[3]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[2]_net_1\, S => \memwaddr_r_s[3]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[3]_net_1\);
    
    \rptr_gray[1]\ : SLE
      port map(D => \rptr_gray_1[1]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[1]_net_1\);
    
    \memwaddr_r[7]\ : SLE
      port map(D => \memwaddr_r_s[7]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[7]\);
    
    \memraddr_r_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[2]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[1]_net_1\, S => \memraddr_r_s[2]\, Y => 
        OPEN, FCO => \memraddr_r_cry[2]_net_1\);
    
    \wptr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[3]_net_1\, S
         => \wptr_s[4]\, Y => OPEN, FCO => \wptr_cry[4]_net_1\);
    
    \memraddr_r_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[8]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[7]_net_1\, S => \memraddr_r_s[8]\, Y => 
        OPEN, FCO => \memraddr_r_cry[8]_net_1\);
    
    \wptr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[9]_net_1\, S
         => \wptr_s[10]\, Y => OPEN, FCO => \wptr_cry[10]_net_1\);
    
    wdiff_bus_cry_5 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[5]_net_1\, B => 
        \rptr_bin_sync2[5]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_4\, S => \wdiff_bus[5]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_5\);
    
    \memwaddr_r[4]\ : SLE
      port map(D => \memwaddr_r_s[4]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[4]\);
    
    \wptr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[1]_net_1\, S
         => \wptr_s[2]\, Y => OPEN, FCO => \wptr_cry[2]_net_1\);
    
    wdiff_bus_cry_0 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[0]_net_1\, B => 
        \rptr_bin_sync2[0]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => VCC_net_1, S => OPEN, Y => wdiff_bus_cry_0_Y, FCO
         => \wdiff_bus_cry_0\);
    
    \wptr[1]\ : SLE
      port map(D => \wptr_s[1]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[1]_net_1\);
    
    \rptr_bin_sync2[4]\ : SLE
      port map(D => \rptr_bin_sync[4]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[4]_net_1\);
    
    \wptr_bin_sync2[6]\ : SLE
      port map(D => \wptr_bin_sync[6]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[6]_net_1\);
    
    \rptr[3]\ : SLE
      port map(D => \rptr_s[3]\, CLK => BIT_CLK, EN => \N_744_i\, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[3]_net_1\);
    
    \wptr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[2]_net_1\, S
         => \wptr_s[3]\, Y => OPEN, FCO => \wptr_cry[3]_net_1\);
    
    \L1.empty_r_3_0_a2_8\ : CFG4
      generic map(INIT => x"0004")

      port map(A => \rdiff_bus[11]\, B => empty_r_3_0_a2_6, C => 
        \rdiff_bus[2]\, D => \rdiff_bus[1]\, Y => 
        empty_r_3_0_a2_8);
    
    \rptr[6]\ : SLE
      port map(D => \rptr_s[6]\, CLK => BIT_CLK, EN => \N_744_i\, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[6]_net_1\);
    
    rdiff_bus_cry_8 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[8]_net_1\, B => 
        \rptr[8]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_7\, S => \rdiff_bus[8]\, Y => OPEN, FCO
         => \rdiff_bus_cry_8\);
    
    \wptr_gray[10]\ : SLE
      port map(D => \wptr_gray_1[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[10]_net_1\);
    
    rdiff_bus_cry_7 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[7]_net_1\, B => 
        \rptr[7]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_6\, S => \rdiff_bus[7]\, Y => OPEN, FCO
         => \rdiff_bus_cry_7\);
    
    \wptr_bin_sync2[7]\ : SLE
      port map(D => \wptr_bin_sync[7]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[7]_net_1\);
    
    overflow_r_RNIDBD3 : CFG1
      generic map(INIT => "01")

      port map(A => \TX_FIFO_OVERFLOW\, Y => TX_FIFO_OVERFLOW_i);
    
    \rptr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[8]_net_1\, S
         => \rptr_s[9]\, Y => OPEN, FCO => \rptr_cry[9]_net_1\);
    
    \T11.un4_fullilto10_i_a2_8\ : CFG4
      generic map(INIT => x"4000")

      port map(A => wdiff_bus_cry_0_Y, B => \wdiff_bus[1]\, C => 
        \wdiff_bus[10]\, D => un4_fullilto10_i_a2_6, Y => 
        un4_fullilto10_i_a2_8);
    
    \rptr_gray[5]\ : SLE
      port map(D => \rptr_gray_1[5]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[5]_net_1\);
    
    \wptr_gray_1[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[2]_net_1\, B => \wptr[3]_net_1\, Y => 
        \wptr_gray_1[2]_net_1\);
    
    \wptr[5]\ : SLE
      port map(D => \wptr_s[5]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[5]_net_1\);
    
    rdiff_bus_cry_5 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[5]_net_1\, B => 
        \rptr[5]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_4\, S => \rdiff_bus[5]\, Y => OPEN, FCO
         => \rdiff_bus_cry_5\);
    
    \wptr_bin_sync2[8]\ : SLE
      port map(D => \wptr_bin_sync[8]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[8]_net_1\);
    
    \wptr[7]\ : SLE
      port map(D => \wptr_s[7]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[7]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \wptr_gray[1]\ : SLE
      port map(D => \wptr_gray_1[1]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[1]_net_1\);
    
    \rptr_gray_1[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[9]_net_1\, B => \rptr[10]_net_1\, Y => 
        \rptr_gray_1[9]_net_1\);
    
    \rptr_bin_sync2[5]\ : SLE
      port map(D => \rptr_bin_sync[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[5]_net_1\);
    
    \rptr_bin_sync2[1]\ : SLE
      port map(D => \rptr_bin_sync[1]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[1]_net_1\);
    
    \memwaddr_r[10]\ : SLE
      port map(D => \memwaddr_r_s[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[10]\);
    
    wdiff_bus_cry_7 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[7]_net_1\, B => 
        \rptr_bin_sync2[7]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_6\, S => \wdiff_bus[7]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_7\);
    
    \wptr_bin_sync2[0]\ : SLE
      port map(D => \wptr_bin_sync[0]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        rdiff_bus);
    
    rdiff_bus_s_11 : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \rptr[11]_net_1\, C => 
        \wptr_bin_sync2[11]_net_1\, D => GND_net_1, FCI => 
        \rdiff_bus_cry_10\, S => \rdiff_bus[11]\, Y => OPEN, FCO
         => OPEN);
    
    \memwaddr_r_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[8]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[7]_net_1\, S => \memwaddr_r_s[8]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[8]_net_1\);
    
    \wptr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => wptr_s_386_FCO, S => 
        \wptr_s[1]\, Y => OPEN, FCO => \wptr_cry[1]_net_1\);
    
    \memraddr_r[8]\ : SLE
      port map(D => \memraddr_r_s[8]\, CLK => BIT_CLK, EN => 
        \N_744_i\, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[8]\);
    
    \rptr[9]\ : SLE
      port map(D => \rptr_s[9]\, CLK => BIT_CLK, EN => \N_744_i\, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[9]_net_1\);
    
    \wptr_gray_1[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[6]_net_1\, B => \wptr[7]_net_1\, Y => 
        \wptr_gray_1[6]_net_1\);
    
    \wptr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[6]_net_1\, S
         => \wptr_s[7]\, Y => OPEN, FCO => \wptr_cry[7]_net_1\);
    
    \wptr_bin_sync2[2]\ : SLE
      port map(D => \wptr_bin_sync[2]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[2]_net_1\);
    
    \T11.un4_fullilto10_i_a2_6\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \wdiff_bus[2]\, B => \wdiff_bus[3]\, C => 
        \wdiff_bus[5]\, D => \wdiff_bus[4]\, Y => 
        un4_fullilto10_i_a2_6);
    
    \rptr_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \rptr[0]_net_1\, Y => \rptr_s[0]\);
    
    \rptr[4]\ : SLE
      port map(D => \rptr_s[4]\, CLK => BIT_CLK, EN => \N_744_i\, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[4]_net_1\);
    
    \memwaddr_r_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[4]_net_1\, S => \memwaddr_r_s[5]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[5]_net_1\);
    
    \memraddr_r_s[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[9]_net_1\, S => \memraddr_r_s[10]_net_1\, 
        Y => OPEN, FCO => OPEN);
    
    \wptr_gray[6]\ : SLE
      port map(D => \wptr_gray_1[6]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[6]_net_1\);
    
    \wptr_gray_1[3]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[3]_net_1\, B => \wptr[4]_net_1\, Y => 
        \wptr_gray_1[3]_net_1\);
    
    \wptr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[4]_net_1\, S
         => \wptr_s[5]\, Y => OPEN, FCO => \wptr_cry[5]_net_1\);
    
    \memraddr_r_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[4]_net_1\, S => \memraddr_r_s[5]\, Y => 
        OPEN, FCO => \memraddr_r_cry[5]_net_1\);
    
    \memraddr_r_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[1]\, C => 
        GND_net_1, D => GND_net_1, FCI => memraddr_r_s_388_FCO, S
         => \memraddr_r_s[1]\, Y => OPEN, FCO => 
        \memraddr_r_cry[1]_net_1\);
    
    \rptr_gray[4]\ : SLE
      port map(D => \rptr_gray_1[4]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[4]_net_1\);
    
    \wptr_bin_sync2[4]\ : SLE
      port map(D => \wptr_bin_sync[4]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[4]_net_1\);
    
    \L1.empty_r_3_0_a2_6\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \rdiff_bus[3]\, B => \rdiff_bus[4]\, C => 
        \rdiff_bus[5]\, D => \rdiff_bus[6]\, Y => 
        empty_r_3_0_a2_6);
    
    \wptr[3]\ : SLE
      port map(D => \wptr_s[3]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[3]_net_1\);
    
    \memwaddr_r[6]\ : SLE
      port map(D => \memwaddr_r_s[6]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[6]\);
    
    memwe_0_a2 : CFG2
      generic map(INIT => x"4")

      port map(A => \TX_FIFO_Full\, B => TX_FIFO_wr_en, Y => 
        \fifo_MEMWE\);
    
    \wptr_s[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[10]_net_1\, S
         => \wptr_s[11]_net_1\, Y => OPEN, FCO => OPEN);
    
    \wptr[6]\ : SLE
      port map(D => \wptr_s[6]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[6]_net_1\);
    
    \memwaddr_r[9]\ : SLE
      port map(D => \memwaddr_r_s[9]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[9]\);
    
    \memraddr_r_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[3]_net_1\, S => \memraddr_r_s[4]\, Y => 
        OPEN, FCO => \memraddr_r_cry[4]_net_1\);
    
    \memraddr_r[10]\ : SLE
      port map(D => \memraddr_r_s[10]_net_1\, CLK => BIT_CLK, EN
         => \N_744_i\, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \fifo_MEMRADDR[10]\);
    
    \memwaddr_r[3]\ : SLE
      port map(D => \memwaddr_r_s[3]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[3]\);
    
    full_r : SLE
      port map(D => \fulli\, CLK => m2s010_som_sb_0_CCC_71MHz, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \TX_FIFO_Full\);
    
    \rptr_bin_sync2[3]\ : SLE
      port map(D => \rptr_bin_sync[3]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[3]_net_1\);
    
    \wptr_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \wptr[0]_net_1\, Y => \wptr_s[0]\);
    
    \rptr[2]\ : SLE
      port map(D => \rptr_s[2]\, CLK => BIT_CLK, EN => \N_744_i\, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[2]_net_1\);
    
    \memraddr_r[3]\ : SLE
      port map(D => \memraddr_r_s[3]\, CLK => BIT_CLK, EN => 
        \N_744_i\, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[3]\);
    
    \rptr_bin_sync2[9]\ : SLE
      port map(D => \rptr_bin_sync[9]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[9]_net_1\);
    
    \rptr[11]\ : SLE
      port map(D => \rptr_s[11]_net_1\, CLK => BIT_CLK, EN => 
        \N_744_i\, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rptr[11]_net_1\);
    
    \L1.un2_re_p_i_0_o2_RNICFVI\ : CFG2
      generic map(INIT => x"2")

      port map(A => \N_432_i\, B => \TX_FIFO_Empty\, Y => 
        \N_744_i\);
    
    \wptr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[5]_net_1\, S
         => \wptr_s[6]\, Y => OPEN, FCO => \wptr_cry[6]_net_1\);
    
    \rptr_bin_sync2[11]\ : SLE
      port map(D => \rptr_bin_sync[11]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[11]_net_1\);
    
    \wptr_bin_sync2[5]\ : SLE
      port map(D => \wptr_bin_sync[5]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[5]_net_1\);
    
    \wptr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[7]_net_1\, S
         => \wptr_s[8]\, Y => OPEN, FCO => \wptr_cry[8]_net_1\);
    
    \wptr_bin_sync2[1]\ : SLE
      port map(D => \wptr_bin_sync[1]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[1]_net_1\);
    
    Wr_corefifo_grayToBinConv : 
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv_0
      port map(wptr_bin_sync(11) => \wptr_bin_sync[11]\, 
        wptr_bin_sync(10) => \wptr_bin_sync[10]\, 
        wptr_bin_sync(9) => \wptr_bin_sync[9]\, wptr_bin_sync(8)
         => \wptr_bin_sync[8]\, wptr_bin_sync(7) => 
        \wptr_bin_sync[7]\, wptr_bin_sync(6) => 
        \wptr_bin_sync[6]\, wptr_bin_sync(5) => 
        \wptr_bin_sync[5]\, wptr_bin_sync(4) => 
        \wptr_bin_sync[4]\, wptr_bin_sync(3) => nc1, 
        wptr_bin_sync(2) => \wptr_bin_sync[2]\, wptr_bin_sync(1)
         => \wptr_bin_sync[1]\, wptr_bin_sync(0) => 
        \wptr_bin_sync[0]\, wptr_gray_sync(10) => 
        \wptr_gray_sync[10]\, wptr_gray_sync(9) => 
        \wptr_gray_sync[9]\, wptr_gray_sync(8) => 
        \wptr_gray_sync[8]\, wptr_gray_sync(7) => 
        \wptr_gray_sync[7]\, wptr_gray_sync(6) => 
        \wptr_gray_sync[6]\, wptr_gray_sync(5) => 
        \wptr_gray_sync[5]\, wptr_gray_sync(4) => 
        \wptr_gray_sync[4]\, wptr_gray_sync(3) => 
        \wptr_gray_sync[3]\, wptr_gray_sync(2) => 
        \wptr_gray_sync[2]\, wptr_gray_sync(1) => 
        \wptr_gray_sync[1]\, wptr_gray_sync(0) => 
        \wptr_gray_sync[0]\, bin_N_4_0_i => bin_N_4_0_i);
    
    \wptr_gray_1[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[4]_net_1\, B => \wptr[5]_net_1\, Y => 
        \wptr_gray_1[4]_net_1\);
    
    overflow_r : SLE
      port map(D => N_1349_i, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \TX_FIFO_OVERFLOW\);
    
    \memraddr_r_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \fifo_MEMRADDR[0]\, Y => \memraddr_r_s[0]\);
    
    \rptr_gray[11]\ : SLE
      port map(D => \rptr[11]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[11]_net_1\);
    
    \wptr_bin_sync2[10]\ : SLE
      port map(D => \wptr_bin_sync[10]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[10]_net_1\);
    
    \rptr[10]\ : SLE
      port map(D => \rptr_s[10]\, CLK => BIT_CLK, EN => \N_744_i\, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[10]_net_1\);
    
    \wptr[9]\ : SLE
      port map(D => \wptr_s[9]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[9]_net_1\);
    
    Wr_corefifo_doubleSync : 
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_1
      port map(wptr_gray(11) => \wptr_gray[11]_net_1\, 
        wptr_gray(10) => \wptr_gray[10]_net_1\, wptr_gray(9) => 
        \wptr_gray[9]_net_1\, wptr_gray(8) => 
        \wptr_gray[8]_net_1\, wptr_gray(7) => 
        \wptr_gray[7]_net_1\, wptr_gray(6) => 
        \wptr_gray[6]_net_1\, wptr_gray(5) => 
        \wptr_gray[5]_net_1\, wptr_gray(4) => 
        \wptr_gray[4]_net_1\, wptr_gray(3) => 
        \wptr_gray[3]_net_1\, wptr_gray(2) => 
        \wptr_gray[2]_net_1\, wptr_gray(1) => 
        \wptr_gray[1]_net_1\, wptr_gray(0) => 
        \wptr_gray[0]_net_1\, wptr_gray_sync(10) => 
        \wptr_gray_sync[10]\, wptr_gray_sync(9) => 
        \wptr_gray_sync[9]\, wptr_gray_sync(8) => 
        \wptr_gray_sync[8]\, wptr_gray_sync(7) => 
        \wptr_gray_sync[7]\, wptr_gray_sync(6) => 
        \wptr_gray_sync[6]\, wptr_gray_sync(5) => 
        \wptr_gray_sync[5]\, wptr_gray_sync(4) => 
        \wptr_gray_sync[4]\, wptr_gray_sync(3) => 
        \wptr_gray_sync[3]\, wptr_gray_sync(2) => 
        \wptr_gray_sync[2]\, wptr_gray_sync(1) => 
        \wptr_gray_sync[1]\, wptr_gray_sync(0) => 
        \wptr_gray_sync[0]\, wptr_bin_sync_0 => 
        \wptr_bin_sync[11]\, BIT_CLK => BIT_CLK, itx_fifo_rst_i
         => itx_fifo_rst_i);
    
    \rptr_gray[0]\ : SLE
      port map(D => \rptr_gray_1[0]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[0]_net_1\);
    
    empty_r : SLE
      port map(D => empty_r_3, CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => GND_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \TX_FIFO_Empty\);
    
    \memwaddr_r_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \fifo_MEMWADDR[0]\, Y => \memwaddr_r_s[0]\);
    
    \T11.un4_fullilto10_i_a2_7\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \wdiff_bus[6]\, B => \wdiff_bus[7]\, C => 
        \wdiff_bus[8]\, D => \wdiff_bus[9]\, Y => 
        un4_fullilto10_i_a2_7);
    
    \rptr_gray_1[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[7]_net_1\, B => \rptr[8]_net_1\, Y => 
        \rptr_gray_1[7]_net_1\);
    
    \wptr[4]\ : SLE
      port map(D => \wptr_s[4]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[4]_net_1\);
    
    \memwaddr_r[8]\ : SLE
      port map(D => \memwaddr_r_s[8]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[8]\);
    
    \memwaddr_r[2]\ : SLE
      port map(D => \memwaddr_r_s[2]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[2]\);
    
    \wptr_bin_sync2[11]\ : SLE
      port map(D => \wptr_bin_sync[11]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[11]_net_1\);
    
    \wptr_gray_1[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[1]_net_1\, B => \wptr[2]_net_1\, Y => 
        \wptr_gray_1[1]_net_1\);
    
    underflow_r : SLE
      port map(D => N_416_i, CLK => BIT_CLK, EN => VCC_net_1, ALn
         => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_FIFO_UNDERRUN\);
    
    \memwaddr_r_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[6]_net_1\, S => \memwaddr_r_s[7]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[7]_net_1\);
    
    \wptr_gray[5]\ : SLE
      port map(D => \wptr_gray_1[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[5]_net_1\);
    
    overflow_r_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => \TX_FIFO_Full\, B => TX_FIFO_wr_en, Y => 
        N_1349_i);
    
    \memraddr_r[7]\ : SLE
      port map(D => \memraddr_r_s[7]\, CLK => BIT_CLK, EN => 
        \N_744_i\, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[7]\);
    
    \rptr_bin_sync2[10]\ : SLE
      port map(D => \rptr_bin_sync[10]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[10]_net_1\);
    
    wdiff_bus_cry_10 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[10]_net_1\, B => 
        \rptr_bin_sync2[10]_net_1\, C => GND_net_1, D => 
        GND_net_1, FCI => \wdiff_bus_cry_9\, S => \wdiff_bus[10]\, 
        Y => OPEN, FCO => \wdiff_bus_cry_10\);
    
    \memwaddr_r_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[9]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[8]_net_1\, S => \memwaddr_r_s[9]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[9]_net_1\);
    
    \wptr_gray[8]\ : SLE
      port map(D => \wptr_gray_1[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[8]_net_1\);
    
    \wptr_gray[7]\ : SLE
      port map(D => \wptr_gray_1[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[7]_net_1\);
    
    \wptr_gray_1[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[5]_net_1\, B => \wptr[6]_net_1\, Y => 
        \wptr_gray_1[5]_net_1\);
    
    \memwaddr_r[5]\ : SLE
      port map(D => \memwaddr_r_s[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[5]\);
    
    \L1.empty_r_3_0_a2\ : CFG4
      generic map(INIT => x"E000")

      port map(A => rdiff_bus_cry_0_Y, B => \N_432_i\, C => 
        empty_r_3_0_a2_7, D => empty_r_3_0_a2_8, Y => empty_r_3);
    
    \rptr[8]\ : SLE
      port map(D => \rptr_s[8]\, CLK => BIT_CLK, EN => \N_744_i\, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[8]_net_1\);
    
    Rd_corefifo_doubleSync : 
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_0
      port map(rptr_gray(11) => \rptr_gray[11]_net_1\, 
        rptr_gray(10) => \rptr_gray[10]_net_1\, rptr_gray(9) => 
        \rptr_gray[9]_net_1\, rptr_gray(8) => 
        \rptr_gray[8]_net_1\, rptr_gray(7) => 
        \rptr_gray[7]_net_1\, rptr_gray(6) => 
        \rptr_gray[6]_net_1\, rptr_gray(5) => 
        \rptr_gray[5]_net_1\, rptr_gray(4) => 
        \rptr_gray[4]_net_1\, rptr_gray(3) => 
        \rptr_gray[3]_net_1\, rptr_gray(2) => 
        \rptr_gray[2]_net_1\, rptr_gray(1) => 
        \rptr_gray[1]_net_1\, rptr_gray(0) => 
        \rptr_gray[0]_net_1\, rptr_gray_sync(10) => 
        \rptr_gray_sync[10]\, rptr_gray_sync(9) => 
        \rptr_gray_sync[9]\, rptr_gray_sync(8) => 
        \rptr_gray_sync[8]\, rptr_gray_sync(7) => 
        \rptr_gray_sync[7]\, rptr_gray_sync(6) => 
        \rptr_gray_sync[6]\, rptr_gray_sync(5) => 
        \rptr_gray_sync[5]\, rptr_gray_sync(4) => 
        \rptr_gray_sync[4]\, rptr_gray_sync(3) => 
        \rptr_gray_sync[3]\, rptr_gray_sync(2) => 
        \rptr_gray_sync[2]\, rptr_gray_sync(1) => 
        \rptr_gray_sync[1]\, rptr_gray_sync(0) => 
        \rptr_gray_sync[0]\, rptr_bin_sync_0 => 
        \rptr_bin_sync[11]\, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, itx_fifo_rst_i => 
        itx_fifo_rst_i);
    
    underflow_r_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => \N_432_i\, B => \TX_FIFO_Empty\, Y => N_416_i);
    
    \rptr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[3]_net_1\, S
         => \rptr_s[4]\, Y => OPEN, FCO => \rptr_cry[4]_net_1\);
    
    wdiff_bus_cry_2 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[2]_net_1\, B => 
        \rptr_bin_sync2[2]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_1\, S => \wdiff_bus[2]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_2\);
    
    \rptr_gray[2]\ : SLE
      port map(D => \rptr_gray_1[2]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[2]_net_1\);
    
    \wptr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[8]_net_1\, S
         => \wptr_s[9]\, Y => OPEN, FCO => \wptr_cry[9]_net_1\);
    
    \wptr_bin_sync2[3]\ : SLE
      port map(D => bin_N_4_0_i, CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[3]_net_1\);
    
    \wptr[2]\ : SLE
      port map(D => \wptr_s[2]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[2]_net_1\);
    
    \rptr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[1]_net_1\, S
         => \rptr_s[2]\, Y => OPEN, FCO => \rptr_cry[2]_net_1\);
    
    rdiff_bus_cry_9 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[9]_net_1\, B => 
        \rptr[9]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_8\, S => \rdiff_bus[9]\, Y => OPEN, FCO
         => \rdiff_bus_cry_9\);
    
    \memwaddr_r[0]\ : SLE
      port map(D => \memwaddr_r_s[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[0]\);
    
    \wptr_gray[2]\ : SLE
      port map(D => \wptr_gray_1[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[2]_net_1\);
    
    wdiff_bus_cry_4 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[4]_net_1\, B => 
        \rptr_bin_sync2[4]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_3\, S => \wdiff_bus[4]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_4\);
    
    \memwaddr_r_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[2]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[1]_net_1\, S => \memwaddr_r_s[2]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[2]_net_1\);
    
    \wptr_gray[11]\ : SLE
      port map(D => \wptr[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[11]_net_1\);
    
    \wptr_bin_sync2[9]\ : SLE
      port map(D => \wptr_bin_sync[9]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[9]_net_1\);
    
    \rptr_gray_1[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[6]_net_1\, B => \rptr[7]_net_1\, Y => 
        \rptr_gray_1[6]_net_1\);
    
    \wptr_gray_1[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[11]_net_1\, B => \wptr[10]_net_1\, Y
         => \wptr_gray_1[10]_net_1\);
    
    wdiff_bus_cry_6 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[6]_net_1\, B => 
        \rptr_bin_sync2[6]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_5\, S => \wdiff_bus[6]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_6\);
    
    \rptr_s[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[10]_net_1\, S
         => \rptr_s[11]_net_1\, Y => OPEN, FCO => OPEN);
    
    \rptr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[2]_net_1\, S
         => \rptr_s[3]\, Y => OPEN, FCO => \rptr_cry[3]_net_1\);
    
    \memraddr_r[4]\ : SLE
      port map(D => \memraddr_r_s[4]\, CLK => BIT_CLK, EN => 
        \N_744_i\, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[4]\);
    
    \memraddr_r_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[6]_net_1\, S => \memraddr_r_s[7]\, Y => 
        OPEN, FCO => \memraddr_r_cry[7]_net_1\);
    
    memraddr_r_s_388 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[0]\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => memraddr_r_s_388_FCO);
    
    \memraddr_r_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[9]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[8]_net_1\, S => \memraddr_r_s[9]\, Y => 
        OPEN, FCO => \memraddr_r_cry[9]_net_1\);
    
    \memraddr_r[5]\ : SLE
      port map(D => \memraddr_r_s[5]\, CLK => BIT_CLK, EN => 
        \N_744_i\, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[5]\);
    
    \rptr_gray[6]\ : SLE
      port map(D => \rptr_gray_1[6]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[6]_net_1\);
    
    \memraddr_r[9]\ : SLE
      port map(D => \memraddr_r_s[9]\, CLK => BIT_CLK, EN => 
        \N_744_i\, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[9]\);
    
    \rptr[0]\ : SLE
      port map(D => \rptr_s[0]\, CLK => BIT_CLK, EN => \N_744_i\, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[0]_net_1\);
    
    \wptr[10]\ : SLE
      port map(D => \wptr_s[10]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \wptr[10]_net_1\);
    
    \memwaddr_r_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[3]_net_1\, S => \memwaddr_r_s[4]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[4]_net_1\);
    
    \memraddr_r_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[3]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[2]_net_1\, S => \memraddr_r_s[3]\, Y => 
        OPEN, FCO => \memraddr_r_cry[3]_net_1\);
    
    wdiff_bus_cry_1 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[1]_net_1\, B => 
        \rptr_bin_sync2[1]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_0\, S => \wdiff_bus[1]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_1\);
    
    rdiff_bus_cry_2 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[2]_net_1\, B => 
        \rptr[2]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_1\, S => \rdiff_bus[2]\, Y => OPEN, FCO
         => \rdiff_bus_cry_2\);
    
    \wptr_gray[9]\ : SLE
      port map(D => \wptr_gray_1[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[9]_net_1\);
    
    \rptr_gray_1[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[4]_net_1\, B => \rptr[5]_net_1\, Y => 
        \rptr_gray_1[4]_net_1\);
    
    \wptr_gray_1[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[8]_net_1\, B => \wptr[9]_net_1\, Y => 
        \wptr_gray_1[8]_net_1\);
    
    Rd_corefifo_grayToBinConv : 
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv
      port map(rptr_bin_sync(11) => \rptr_bin_sync[11]\, 
        rptr_bin_sync(10) => \rptr_bin_sync[10]\, 
        rptr_bin_sync(9) => \rptr_bin_sync[9]\, rptr_bin_sync(8)
         => \rptr_bin_sync[8]\, rptr_bin_sync(7) => 
        \rptr_bin_sync[7]\, rptr_bin_sync(6) => 
        \rptr_bin_sync[6]\, rptr_bin_sync(5) => 
        \rptr_bin_sync[5]\, rptr_bin_sync(4) => 
        \rptr_bin_sync[4]\, rptr_bin_sync(3) => 
        \rptr_bin_sync[3]\, rptr_bin_sync(2) => 
        \rptr_bin_sync[2]\, rptr_bin_sync(1) => 
        \rptr_bin_sync[1]\, rptr_bin_sync(0) => 
        \rptr_bin_sync[0]\, rptr_gray_sync(10) => 
        \rptr_gray_sync[10]\, rptr_gray_sync(9) => 
        \rptr_gray_sync[9]\, rptr_gray_sync(8) => 
        \rptr_gray_sync[8]\, rptr_gray_sync(7) => 
        \rptr_gray_sync[7]\, rptr_gray_sync(6) => 
        \rptr_gray_sync[6]\, rptr_gray_sync(5) => 
        \rptr_gray_sync[5]\, rptr_gray_sync(4) => 
        \rptr_gray_sync[4]\, rptr_gray_sync(3) => 
        \rptr_gray_sync[3]\, rptr_gray_sync(2) => 
        \rptr_gray_sync[2]\, rptr_gray_sync(1) => 
        \rptr_gray_sync[1]\, rptr_gray_sync(0) => 
        \rptr_gray_sync[0]\);
    
    \L1.un2_re_p_i_0_o2\ : CFG4
      generic map(INIT => x"EC00")

      port map(A => TX_DataEn_1_o, B => 
        un1_tx_packet_length_0_sqmuxa_o, C => TX_PreAmble, D => 
        byte_clk_en, Y => \N_432_i\);
    
    \rptr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => rptr_s_389_FCO, S => 
        \rptr_s[1]\, Y => OPEN, FCO => \rptr_cry[1]_net_1\);
    
    rdiff_bus_cry_3 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[3]_net_1\, B => 
        \rptr[3]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_2\, S => \rdiff_bus[3]\, Y => OPEN, FCO
         => \rdiff_bus_cry_3\);
    
    rdiff_bus_cry_10 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[10]_net_1\, B => 
        \rptr[10]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_9\, S => \rdiff_bus[10]\, Y => OPEN, FCO
         => \rdiff_bus_cry_10\);
    
    \memraddr_r_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[5]_net_1\, S => \memraddr_r_s[6]\, Y => 
        OPEN, FCO => \memraddr_r_cry[6]_net_1\);
    
    \memraddr_r[6]\ : SLE
      port map(D => \memraddr_r_s[6]\, CLK => BIT_CLK, EN => 
        \N_744_i\, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[6]\);
    
    \rptr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[6]_net_1\, S
         => \rptr_s[7]\, Y => OPEN, FCO => \rptr_cry[7]_net_1\);
    
    rdiff_bus_cry_0 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => rdiff_bus, B => \rptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => rdiff_bus_cry_0_Y, FCO => \rdiff_bus_cry_0\);
    
    \memraddr_r[2]\ : SLE
      port map(D => \memraddr_r_s[2]\, CLK => BIT_CLK, EN => 
        \N_744_i\, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[2]\);
    
    \wptr[8]\ : SLE
      port map(D => \wptr_s[8]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[8]_net_1\);
    
    wdiff_bus_cry_3 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[3]_net_1\, B => 
        \rptr_bin_sync2[3]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_2\, S => \wdiff_bus[3]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_3\);
    
    memwaddr_r_s_387 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[0]\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => memwaddr_r_s_387_FCO);
    
    \rptr_gray[7]\ : SLE
      port map(D => \rptr_gray_1[7]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[7]_net_1\);
    
    \wptr_gray[0]\ : SLE
      port map(D => \wptr_gray_1[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[0]_net_1\);
    
    \rptr_gray_1[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[0]_net_1\, B => \rptr[1]_net_1\, Y => 
        \rptr_gray_1[0]_net_1\);
    
    \rptr_gray_1[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[8]_net_1\, B => \rptr[9]_net_1\, Y => 
        \rptr_gray_1[8]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_2Kx8_FIFO_2Kx8_0_COREFIFO is

    port( CoreAPB3_0_APBmslave0_PWDATA    : in    std_logic_vector(7 downto 0);
          TX_FIFO_UNDERRUN                : out   std_logic;
          TX_FIFO_UNDERRUN_i              : out   std_logic;
          TX_FIFO_OVERFLOW                : out   std_logic;
          TX_FIFO_OVERFLOW_i              : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz       : in    std_logic;
          TX_FIFO_Full                    : out   std_logic;
          TX_FIFO_wr_en                   : in    std_logic;
          un1_tx_packet_length_0_sqmuxa_o : in    std_logic;
          TX_DataEn_1_o                   : in    std_logic;
          TX_PreAmble                     : in    std_logic;
          N_704                           : out   std_logic;
          N_705                           : out   std_logic;
          N_706                           : out   std_logic;
          N_707                           : out   std_logic;
          N_708                           : out   std_logic;
          N_709                           : out   std_logic;
          N_710                           : out   std_logic;
          N_711                           : out   std_logic;
          byte_clk_en                     : in    std_logic;
          TX_FIFO_Empty                   : out   std_logic;
          BIT_CLK                         : in    std_logic;
          itx_fifo_rst_i                  : in    std_logic
        );

end FIFO_2Kx8_FIFO_2Kx8_0_COREFIFO;

architecture DEF_ARCH of FIFO_2Kx8_FIFO_2Kx8_0_COREFIFO is 

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component FIFO_2Kx8_FIFO_2Kx8_0_ram_wrapper
    port( RDATA_int                    : out   std_logic_vector(7 downto 0);
          fifo_MEMRADDR                : in    std_logic_vector(10 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0) := (others => 'U');
          fifo_MEMWADDR                : in    std_logic_vector(10 downto 0) := (others => 'U');
          BIT_CLK                      : in    std_logic := 'U';
          N_744_i                      : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic := 'U';
          fifo_MEMWE                   : in    std_logic := 'U'
        );
  end component;

  component FIFO_2Kx8_FIFO_2Kx8_0_corefifo_async
    port( fifo_MEMWADDR                   : out   std_logic_vector(10 downto 0);
          fifo_MEMRADDR                   : out   std_logic_vector(10 downto 0);
          N_432_i                         : out   std_logic;
          byte_clk_en                     : in    std_logic := 'U';
          TX_PreAmble                     : in    std_logic := 'U';
          un1_tx_packet_length_0_sqmuxa_o : in    std_logic := 'U';
          TX_DataEn_1_o                   : in    std_logic := 'U';
          TX_FIFO_wr_en                   : in    std_logic := 'U';
          fifo_MEMWE                      : out   std_logic;
          N_744_i                         : out   std_logic;
          TX_FIFO_Full                    : out   std_logic;
          TX_FIFO_Empty                   : out   std_logic;
          BIT_CLK                         : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz       : in    std_logic := 'U';
          itx_fifo_rst_i                  : in    std_logic := 'U';
          TX_FIFO_OVERFLOW_i              : out   std_logic;
          TX_FIFO_OVERFLOW                : out   std_logic;
          TX_FIFO_UNDERRUN_i              : out   std_logic;
          TX_FIFO_UNDERRUN                : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \RDATA_r[5]_net_1\, VCC_net_1, \RDATA_int[5]\, 
        N_415_i, GND_net_1, \RDATA_r[6]_net_1\, \RDATA_int[6]\, 
        \RDATA_r[7]_net_1\, \RDATA_int[7]\, \re_set\, 
        \re_set_ldmx\, N_769_i, \RDATA_r[0]_net_1\, 
        \RDATA_int[0]\, \RDATA_r[1]_net_1\, \RDATA_int[1]\, 
        \RDATA_r[2]_net_1\, \RDATA_int[2]\, \RDATA_r[3]_net_1\, 
        \RDATA_int[3]\, \RDATA_r[4]_net_1\, \RDATA_int[4]\, 
        \REN_d1\, N_744_i, \RE_d1\, N_432_i, \re_pulse_d1\, 
        \re_pulse\, \TX_FIFO_Empty\, \un9_fifo_memre_i_0_a2_0_1\, 
        N_770, \fifo_MEMWADDR[0]\, \fifo_MEMWADDR[1]\, 
        \fifo_MEMWADDR[2]\, \fifo_MEMWADDR[3]\, 
        \fifo_MEMWADDR[4]\, \fifo_MEMWADDR[5]\, 
        \fifo_MEMWADDR[6]\, \fifo_MEMWADDR[7]\, 
        \fifo_MEMWADDR[8]\, \fifo_MEMWADDR[9]\, 
        \fifo_MEMWADDR[10]\, \fifo_MEMRADDR[0]\, 
        \fifo_MEMRADDR[1]\, \fifo_MEMRADDR[2]\, 
        \fifo_MEMRADDR[3]\, \fifo_MEMRADDR[4]\, 
        \fifo_MEMRADDR[5]\, \fifo_MEMRADDR[6]\, 
        \fifo_MEMRADDR[7]\, \fifo_MEMRADDR[8]\, 
        \fifo_MEMRADDR[9]\, \fifo_MEMRADDR[10]\, fifo_MEMWE
         : std_logic;

    for all : FIFO_2Kx8_FIFO_2Kx8_0_ram_wrapper
	Use entity work.FIFO_2Kx8_FIFO_2Kx8_0_ram_wrapper(DEF_ARCH);
    for all : FIFO_2Kx8_FIFO_2Kx8_0_corefifo_async
	Use entity work.FIFO_2Kx8_FIFO_2Kx8_0_corefifo_async(DEF_ARCH);
begin 

    TX_FIFO_Empty <= \TX_FIFO_Empty\;

    un9_fifo_memre_i_0_a2_0_1 : CFG3
      generic map(INIT => x"20")

      port map(A => \REN_d1\, B => \TX_FIFO_Empty\, C => 
        byte_clk_en, Y => \un9_fifo_memre_i_0_a2_0_1\);
    
    re_pulse : CFG4
      generic map(INIT => x"EAEE")

      port map(A => \re_set\, B => \REN_d1\, C => \TX_FIFO_Empty\, 
        D => N_432_i, Y => \re_pulse\);
    
    \RDATA_r[3]\ : SLE
      port map(D => \RDATA_int[3]\, CLK => BIT_CLK, EN => N_415_i, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[3]_net_1\);
    
    re_pulse_d1 : SLE
      port map(D => \re_pulse\, CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \re_pulse_d1\);
    
    \RDATA_r[5]\ : SLE
      port map(D => \RDATA_int[5]\, CLK => BIT_CLK, EN => N_415_i, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[5]_net_1\);
    
    \Q_i_m2_i_m2_i_m2[1]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[1]_net_1\, C => 
        \RDATA_int[1]\, D => \RE_d1\, Y => N_711);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \RW1.UI_ram_wrapper_1\ : FIFO_2Kx8_FIFO_2Kx8_0_ram_wrapper
      port map(RDATA_int(7) => \RDATA_int[7]\, RDATA_int(6) => 
        \RDATA_int[6]\, RDATA_int(5) => \RDATA_int[5]\, 
        RDATA_int(4) => \RDATA_int[4]\, RDATA_int(3) => 
        \RDATA_int[3]\, RDATA_int(2) => \RDATA_int[2]\, 
        RDATA_int(1) => \RDATA_int[1]\, RDATA_int(0) => 
        \RDATA_int[0]\, fifo_MEMRADDR(10) => \fifo_MEMRADDR[10]\, 
        fifo_MEMRADDR(9) => \fifo_MEMRADDR[9]\, fifo_MEMRADDR(8)
         => \fifo_MEMRADDR[8]\, fifo_MEMRADDR(7) => 
        \fifo_MEMRADDR[7]\, fifo_MEMRADDR(6) => 
        \fifo_MEMRADDR[6]\, fifo_MEMRADDR(5) => 
        \fifo_MEMRADDR[5]\, fifo_MEMRADDR(4) => 
        \fifo_MEMRADDR[4]\, fifo_MEMRADDR(3) => 
        \fifo_MEMRADDR[3]\, fifo_MEMRADDR(2) => 
        \fifo_MEMRADDR[2]\, fifo_MEMRADDR(1) => 
        \fifo_MEMRADDR[1]\, fifo_MEMRADDR(0) => 
        \fifo_MEMRADDR[0]\, CoreAPB3_0_APBmslave0_PWDATA(7) => 
        CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), fifo_MEMWADDR(10) => 
        \fifo_MEMWADDR[10]\, fifo_MEMWADDR(9) => 
        \fifo_MEMWADDR[9]\, fifo_MEMWADDR(8) => 
        \fifo_MEMWADDR[8]\, fifo_MEMWADDR(7) => 
        \fifo_MEMWADDR[7]\, fifo_MEMWADDR(6) => 
        \fifo_MEMWADDR[6]\, fifo_MEMWADDR(5) => 
        \fifo_MEMWADDR[5]\, fifo_MEMWADDR(4) => 
        \fifo_MEMWADDR[4]\, fifo_MEMWADDR(3) => 
        \fifo_MEMWADDR[3]\, fifo_MEMWADDR(2) => 
        \fifo_MEMWADDR[2]\, fifo_MEMWADDR(1) => 
        \fifo_MEMWADDR[1]\, fifo_MEMWADDR(0) => 
        \fifo_MEMWADDR[0]\, BIT_CLK => BIT_CLK, N_744_i => 
        N_744_i, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, fifo_MEMWE => fifo_MEMWE);
    
    \Q_i_m2_i_m2_i_m2[5]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[5]_net_1\, C => 
        \RDATA_int[5]\, D => \RE_d1\, Y => N_708);
    
    \RDATA_r[0]\ : SLE
      port map(D => \RDATA_int[0]\, CLK => BIT_CLK, EN => N_415_i, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[0]_net_1\);
    
    \RDATA_r[2]\ : SLE
      port map(D => \RDATA_int[2]\, CLK => BIT_CLK, EN => N_415_i, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[2]_net_1\);
    
    \Q_i_m2_i_m2_i_m2[4]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[4]_net_1\, C => 
        \RDATA_int[4]\, D => \RE_d1\, Y => N_704);
    
    re_set_ldmx : CFG3
      generic map(INIT => x"E2")

      port map(A => \REN_d1\, B => N_770, C => \re_set\, Y => 
        \re_set_ldmx\);
    
    \RDATA_r[6]\ : SLE
      port map(D => \RDATA_int[6]\, CLK => BIT_CLK, EN => N_415_i, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[6]_net_1\);
    
    \Q_i_m2_i_m2_i_m2[7]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[7]_net_1\, C => 
        \RDATA_int[7]\, D => \RE_d1\, Y => N_706);
    
    \Q_i_m2_i_m2_i_m2[3]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[3]_net_1\, C => 
        \RDATA_int[3]\, D => \RE_d1\, Y => N_709);
    
    \Q_i_m2_i_m2_i_m2[2]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[2]_net_1\, C => 
        \RDATA_int[2]\, D => \RE_d1\, Y => N_710);
    
    \Q_i_m2_i_m2_i_m2[6]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[6]_net_1\, C => 
        \RDATA_int[6]\, D => \RE_d1\, Y => N_707);
    
    \L31.U_corefifo_async\ : FIFO_2Kx8_FIFO_2Kx8_0_corefifo_async
      port map(fifo_MEMWADDR(10) => \fifo_MEMWADDR[10]\, 
        fifo_MEMWADDR(9) => \fifo_MEMWADDR[9]\, fifo_MEMWADDR(8)
         => \fifo_MEMWADDR[8]\, fifo_MEMWADDR(7) => 
        \fifo_MEMWADDR[7]\, fifo_MEMWADDR(6) => 
        \fifo_MEMWADDR[6]\, fifo_MEMWADDR(5) => 
        \fifo_MEMWADDR[5]\, fifo_MEMWADDR(4) => 
        \fifo_MEMWADDR[4]\, fifo_MEMWADDR(3) => 
        \fifo_MEMWADDR[3]\, fifo_MEMWADDR(2) => 
        \fifo_MEMWADDR[2]\, fifo_MEMWADDR(1) => 
        \fifo_MEMWADDR[1]\, fifo_MEMWADDR(0) => 
        \fifo_MEMWADDR[0]\, fifo_MEMRADDR(10) => 
        \fifo_MEMRADDR[10]\, fifo_MEMRADDR(9) => 
        \fifo_MEMRADDR[9]\, fifo_MEMRADDR(8) => 
        \fifo_MEMRADDR[8]\, fifo_MEMRADDR(7) => 
        \fifo_MEMRADDR[7]\, fifo_MEMRADDR(6) => 
        \fifo_MEMRADDR[6]\, fifo_MEMRADDR(5) => 
        \fifo_MEMRADDR[5]\, fifo_MEMRADDR(4) => 
        \fifo_MEMRADDR[4]\, fifo_MEMRADDR(3) => 
        \fifo_MEMRADDR[3]\, fifo_MEMRADDR(2) => 
        \fifo_MEMRADDR[2]\, fifo_MEMRADDR(1) => 
        \fifo_MEMRADDR[1]\, fifo_MEMRADDR(0) => 
        \fifo_MEMRADDR[0]\, N_432_i => N_432_i, byte_clk_en => 
        byte_clk_en, TX_PreAmble => TX_PreAmble, 
        un1_tx_packet_length_0_sqmuxa_o => 
        un1_tx_packet_length_0_sqmuxa_o, TX_DataEn_1_o => 
        TX_DataEn_1_o, TX_FIFO_wr_en => TX_FIFO_wr_en, fifo_MEMWE
         => fifo_MEMWE, N_744_i => N_744_i, TX_FIFO_Full => 
        TX_FIFO_Full, TX_FIFO_Empty => \TX_FIFO_Empty\, BIT_CLK
         => BIT_CLK, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, itx_fifo_rst_i => 
        itx_fifo_rst_i, TX_FIFO_OVERFLOW_i => TX_FIFO_OVERFLOW_i, 
        TX_FIFO_OVERFLOW => TX_FIFO_OVERFLOW, TX_FIFO_UNDERRUN_i
         => TX_FIFO_UNDERRUN_i, TX_FIFO_UNDERRUN => 
        TX_FIFO_UNDERRUN);
    
    re_set : SLE
      port map(D => \re_set_ldmx\, CLK => BIT_CLK, EN => N_769_i, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \re_set\);
    
    REN_d1_RNI3O3L : CFG3
      generic map(INIT => x"C4")

      port map(A => N_432_i, B => \REN_d1\, C => \TX_FIFO_Empty\, 
        Y => N_415_i);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    RE_d1 : SLE
      port map(D => N_432_i, CLK => BIT_CLK, EN => VCC_net_1, ALn
         => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \RE_d1\);
    
    \RDATA_r[7]\ : SLE
      port map(D => \RDATA_int[7]\, CLK => BIT_CLK, EN => N_415_i, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[7]_net_1\);
    
    \RDATA_r[4]\ : SLE
      port map(D => \RDATA_int[4]\, CLK => BIT_CLK, EN => N_415_i, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[4]_net_1\);
    
    un9_fifo_memre_i_0_a2_0 : CFG4
      generic map(INIT => x"CC80")

      port map(A => TX_PreAmble, B => \un9_fifo_memre_i_0_a2_0_1\, 
        C => TX_DataEn_1_o, D => un1_tx_packet_length_0_sqmuxa_o, 
        Y => N_770);
    
    \Q_i_m2_i_m2_i_m2[0]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[0]_net_1\, C => 
        \RDATA_int[0]\, D => \RE_d1\, Y => N_705);
    
    REN_d1 : SLE
      port map(D => N_744_i, CLK => BIT_CLK, EN => VCC_net_1, ALn
         => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \REN_d1\);
    
    re_set_RNO : CFG3
      generic map(INIT => x"CE")

      port map(A => N_432_i, B => \REN_d1\, C => \TX_FIFO_Empty\, 
        Y => N_769_i);
    
    \RDATA_r[1]\ : SLE
      port map(D => \RDATA_int[1]\, CLK => BIT_CLK, EN => N_415_i, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[1]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_2Kx8 is

    port( CoreAPB3_0_APBmslave0_PWDATA    : in    std_logic_vector(7 downto 0);
          itx_fifo_rst_i                  : in    std_logic;
          BIT_CLK                         : in    std_logic;
          TX_FIFO_Empty                   : out   std_logic;
          byte_clk_en                     : in    std_logic;
          N_711                           : out   std_logic;
          N_710                           : out   std_logic;
          N_709                           : out   std_logic;
          N_708                           : out   std_logic;
          N_707                           : out   std_logic;
          N_706                           : out   std_logic;
          N_705                           : out   std_logic;
          N_704                           : out   std_logic;
          TX_PreAmble                     : in    std_logic;
          TX_DataEn_1_o                   : in    std_logic;
          un1_tx_packet_length_0_sqmuxa_o : in    std_logic;
          TX_FIFO_wr_en                   : in    std_logic;
          TX_FIFO_Full                    : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz       : in    std_logic;
          TX_FIFO_OVERFLOW_i              : out   std_logic;
          TX_FIFO_OVERFLOW                : out   std_logic;
          TX_FIFO_UNDERRUN_i              : out   std_logic;
          TX_FIFO_UNDERRUN                : out   std_logic
        );

end FIFO_2Kx8;

architecture DEF_ARCH of FIFO_2Kx8 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component FIFO_2Kx8_FIFO_2Kx8_0_COREFIFO
    port( CoreAPB3_0_APBmslave0_PWDATA    : in    std_logic_vector(7 downto 0) := (others => 'U');
          TX_FIFO_UNDERRUN                : out   std_logic;
          TX_FIFO_UNDERRUN_i              : out   std_logic;
          TX_FIFO_OVERFLOW                : out   std_logic;
          TX_FIFO_OVERFLOW_i              : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz       : in    std_logic := 'U';
          TX_FIFO_Full                    : out   std_logic;
          TX_FIFO_wr_en                   : in    std_logic := 'U';
          un1_tx_packet_length_0_sqmuxa_o : in    std_logic := 'U';
          TX_DataEn_1_o                   : in    std_logic := 'U';
          TX_PreAmble                     : in    std_logic := 'U';
          N_704                           : out   std_logic;
          N_705                           : out   std_logic;
          N_706                           : out   std_logic;
          N_707                           : out   std_logic;
          N_708                           : out   std_logic;
          N_709                           : out   std_logic;
          N_710                           : out   std_logic;
          N_711                           : out   std_logic;
          byte_clk_en                     : in    std_logic := 'U';
          TX_FIFO_Empty                   : out   std_logic;
          BIT_CLK                         : in    std_logic := 'U';
          itx_fifo_rst_i                  : in    std_logic := 'U'
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : FIFO_2Kx8_FIFO_2Kx8_0_COREFIFO
	Use entity work.FIFO_2Kx8_FIFO_2Kx8_0_COREFIFO(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    FIFO_2Kx8_0 : FIFO_2Kx8_FIFO_2Kx8_0_COREFIFO
      port map(CoreAPB3_0_APBmslave0_PWDATA(7) => 
        CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), TX_FIFO_UNDERRUN => 
        TX_FIFO_UNDERRUN, TX_FIFO_UNDERRUN_i => 
        TX_FIFO_UNDERRUN_i, TX_FIFO_OVERFLOW => TX_FIFO_OVERFLOW, 
        TX_FIFO_OVERFLOW_i => TX_FIFO_OVERFLOW_i, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz, 
        TX_FIFO_Full => TX_FIFO_Full, TX_FIFO_wr_en => 
        TX_FIFO_wr_en, un1_tx_packet_length_0_sqmuxa_o => 
        un1_tx_packet_length_0_sqmuxa_o, TX_DataEn_1_o => 
        TX_DataEn_1_o, TX_PreAmble => TX_PreAmble, N_704 => N_704, 
        N_705 => N_705, N_706 => N_706, N_707 => N_707, N_708 => 
        N_708, N_709 => N_709, N_710 => N_710, N_711 => N_711, 
        byte_clk_en => byte_clk_en, TX_FIFO_Empty => 
        TX_FIFO_Empty, BIT_CLK => BIT_CLK, itx_fifo_rst_i => 
        itx_fifo_rst_i);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_0 is

    port( fifo_MEMWADDR             : in    std_logic_vector(10 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          fifo_MEMRADDR             : in    std_logic_vector(10 downto 0);
          RDATA_int                 : out   std_logic_vector(8 downto 0);
          fifo_MEMWE                : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          N_140_i                   : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_0;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component RAM1K18
    generic (MEMORYFILE:string := "");

    port( A_DOUT        : out   std_logic_vector(17 downto 0);
          B_DOUT        : out   std_logic_vector(17 downto 0);
          BUSY          : out   std_logic;
          A_CLK         : in    std_logic := 'U';
          A_DOUT_CLK    : in    std_logic := 'U';
          A_ARST_N      : in    std_logic := 'U';
          A_DOUT_EN     : in    std_logic := 'U';
          A_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_DOUT_ARST_N : in    std_logic := 'U';
          A_DOUT_SRST_N : in    std_logic := 'U';
          A_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          A_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          A_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          B_CLK         : in    std_logic := 'U';
          B_DOUT_CLK    : in    std_logic := 'U';
          B_ARST_N      : in    std_logic := 'U';
          B_DOUT_EN     : in    std_logic := 'U';
          B_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_DOUT_ARST_N : in    std_logic := 'U';
          B_DOUT_SRST_N : in    std_logic := 'U';
          B_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          B_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          B_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          A_EN          : in    std_logic := 'U';
          A_DOUT_LAT    : in    std_logic := 'U';
          A_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_WMODE       : in    std_logic := 'U';
          B_EN          : in    std_logic := 'U';
          B_DOUT_LAT    : in    std_logic := 'U';
          B_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_WMODE       : in    std_logic := 'U';
          SII_LOCK      : in    std_logic := 'U'
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;
    signal nc24, nc1, nc8, nc13, nc16, nc19, nc25, nc20, nc27, 
        nc9, nc22, nc14, nc5, nc21, nc15, nc3, nc10, nc7, nc17, 
        nc4, nc12, nc2, nc23, nc18, nc26, nc6, nc11 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C0 : RAM1K18
      port map(A_DOUT(17) => nc24, A_DOUT(16) => nc1, A_DOUT(15)
         => nc8, A_DOUT(14) => nc13, A_DOUT(13) => nc16, 
        A_DOUT(12) => nc19, A_DOUT(11) => nc25, A_DOUT(10) => 
        nc20, A_DOUT(9) => nc27, A_DOUT(8) => RDATA_int(8), 
        A_DOUT(7) => RDATA_int(7), A_DOUT(6) => RDATA_int(6), 
        A_DOUT(5) => RDATA_int(5), A_DOUT(4) => RDATA_int(4), 
        A_DOUT(3) => RDATA_int(3), A_DOUT(2) => RDATA_int(2), 
        A_DOUT(1) => RDATA_int(1), A_DOUT(0) => RDATA_int(0), 
        B_DOUT(17) => nc9, B_DOUT(16) => nc22, B_DOUT(15) => nc14, 
        B_DOUT(14) => nc5, B_DOUT(13) => nc21, B_DOUT(12) => nc15, 
        B_DOUT(11) => nc3, B_DOUT(10) => nc10, B_DOUT(9) => nc7, 
        B_DOUT(8) => nc17, B_DOUT(7) => nc4, B_DOUT(6) => nc12, 
        B_DOUT(5) => nc2, B_DOUT(4) => nc23, B_DOUT(3) => nc18, 
        B_DOUT(2) => nc26, B_DOUT(1) => nc6, B_DOUT(0) => nc11, 
        BUSY => OPEN, A_CLK => m2s010_som_sb_0_CCC_71MHz, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => VCC_net_1, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_140_i, A_BLK(1) => VCC_net_1, 
        A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => VCC_net_1, 
        A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => GND_net_1, 
        A_DIN(16) => GND_net_1, A_DIN(15) => GND_net_1, A_DIN(14)
         => GND_net_1, A_DIN(13) => GND_net_1, A_DIN(12) => 
        GND_net_1, A_DIN(11) => GND_net_1, A_DIN(10) => GND_net_1, 
        A_DIN(9) => GND_net_1, A_DIN(8) => GND_net_1, A_DIN(7)
         => GND_net_1, A_DIN(6) => GND_net_1, A_DIN(5) => 
        GND_net_1, A_DIN(4) => GND_net_1, A_DIN(3) => GND_net_1, 
        A_DIN(2) => GND_net_1, A_DIN(1) => GND_net_1, A_DIN(0)
         => GND_net_1, A_ADDR(13) => fifo_MEMRADDR(10), 
        A_ADDR(12) => fifo_MEMRADDR(9), A_ADDR(11) => 
        fifo_MEMRADDR(8), A_ADDR(10) => fifo_MEMRADDR(7), 
        A_ADDR(9) => fifo_MEMRADDR(6), A_ADDR(8) => 
        fifo_MEMRADDR(5), A_ADDR(7) => fifo_MEMRADDR(4), 
        A_ADDR(6) => fifo_MEMRADDR(3), A_ADDR(5) => 
        fifo_MEMRADDR(2), A_ADDR(4) => fifo_MEMRADDR(1), 
        A_ADDR(3) => fifo_MEMRADDR(0), A_ADDR(2) => GND_net_1, 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => RX_FIFO_DIN_pipe(8), B_DIN(7) => RX_FIFO_DIN_pipe(7), 
        B_DIN(6) => RX_FIFO_DIN_pipe(6), B_DIN(5) => 
        RX_FIFO_DIN_pipe(5), B_DIN(4) => RX_FIFO_DIN_pipe(4), 
        B_DIN(3) => RX_FIFO_DIN_pipe(3), B_DIN(2) => 
        RX_FIFO_DIN_pipe(2), B_DIN(1) => RX_FIFO_DIN_pipe(1), 
        B_DIN(0) => RX_FIFO_DIN_pipe(0), B_ADDR(13) => 
        fifo_MEMWADDR(10), B_ADDR(12) => fifo_MEMWADDR(9), 
        B_ADDR(11) => fifo_MEMWADDR(8), B_ADDR(10) => 
        fifo_MEMWADDR(7), B_ADDR(9) => fifo_MEMWADDR(6), 
        B_ADDR(8) => fifo_MEMWADDR(5), B_ADDR(7) => 
        fifo_MEMWADDR(4), B_ADDR(6) => fifo_MEMWADDR(3), 
        B_ADDR(5) => fifo_MEMWADDR(2), B_ADDR(4) => 
        fifo_MEMWADDR(1), B_ADDR(3) => fifo_MEMWADDR(0), 
        B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, B_ADDR(0)
         => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0) => 
        VCC_net_1, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_0 is

    port( RDATA_int                 : out   std_logic_vector(8 downto 0);
          fifo_MEMRADDR             : in    std_logic_vector(10 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          fifo_MEMWADDR             : in    std_logic_vector(10 downto 0);
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          N_140_i                   : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          fifo_MEMWE                : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_0;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_0
    port( fifo_MEMWADDR             : in    std_logic_vector(10 downto 0) := (others => 'U');
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          fifo_MEMRADDR             : in    std_logic_vector(10 downto 0) := (others => 'U');
          RDATA_int                 : out   std_logic_vector(8 downto 0);
          fifo_MEMWE                : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          N_140_i                   : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_0
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_0(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    L1_asyncnonpipe : FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_0
      port map(fifo_MEMWADDR(10) => fifo_MEMWADDR(10), 
        fifo_MEMWADDR(9) => fifo_MEMWADDR(9), fifo_MEMWADDR(8)
         => fifo_MEMWADDR(8), fifo_MEMWADDR(7) => 
        fifo_MEMWADDR(7), fifo_MEMWADDR(6) => fifo_MEMWADDR(6), 
        fifo_MEMWADDR(5) => fifo_MEMWADDR(5), fifo_MEMWADDR(4)
         => fifo_MEMWADDR(4), fifo_MEMWADDR(3) => 
        fifo_MEMWADDR(3), fifo_MEMWADDR(2) => fifo_MEMWADDR(2), 
        fifo_MEMWADDR(1) => fifo_MEMWADDR(1), fifo_MEMWADDR(0)
         => fifo_MEMWADDR(0), RX_FIFO_DIN_pipe(8) => 
        RX_FIFO_DIN_pipe(8), RX_FIFO_DIN_pipe(7) => 
        RX_FIFO_DIN_pipe(7), RX_FIFO_DIN_pipe(6) => 
        RX_FIFO_DIN_pipe(6), RX_FIFO_DIN_pipe(5) => 
        RX_FIFO_DIN_pipe(5), RX_FIFO_DIN_pipe(4) => 
        RX_FIFO_DIN_pipe(4), RX_FIFO_DIN_pipe(3) => 
        RX_FIFO_DIN_pipe(3), RX_FIFO_DIN_pipe(2) => 
        RX_FIFO_DIN_pipe(2), RX_FIFO_DIN_pipe(1) => 
        RX_FIFO_DIN_pipe(1), RX_FIFO_DIN_pipe(0) => 
        RX_FIFO_DIN_pipe(0), fifo_MEMRADDR(10) => 
        fifo_MEMRADDR(10), fifo_MEMRADDR(9) => fifo_MEMRADDR(9), 
        fifo_MEMRADDR(8) => fifo_MEMRADDR(8), fifo_MEMRADDR(7)
         => fifo_MEMRADDR(7), fifo_MEMRADDR(6) => 
        fifo_MEMRADDR(6), fifo_MEMRADDR(5) => fifo_MEMRADDR(5), 
        fifo_MEMRADDR(4) => fifo_MEMRADDR(4), fifo_MEMRADDR(3)
         => fifo_MEMRADDR(3), fifo_MEMRADDR(2) => 
        fifo_MEMRADDR(2), fifo_MEMRADDR(1) => fifo_MEMRADDR(1), 
        fifo_MEMRADDR(0) => fifo_MEMRADDR(0), RDATA_int(8) => 
        RDATA_int(8), RDATA_int(7) => RDATA_int(7), RDATA_int(6)
         => RDATA_int(6), RDATA_int(5) => RDATA_int(5), 
        RDATA_int(4) => RDATA_int(4), RDATA_int(3) => 
        RDATA_int(3), RDATA_int(2) => RDATA_int(2), RDATA_int(1)
         => RDATA_int(1), RDATA_int(0) => RDATA_int(0), 
        fifo_MEMWE => fifo_MEMWE, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, N_140_i => N_140_i, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_2 is

    port( wptr_bin_sync  : inout std_logic_vector(11 downto 0) := (others => 'Z');
          wptr_gray_sync : in    std_logic_vector(10 downto 0)
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_2;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_2 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    \bin_out_xhdl1_0_a2[1]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(3), B => wptr_gray_sync(1), C
         => wptr_bin_sync(4), D => wptr_gray_sync(2), Y => 
        wptr_bin_sync(1));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \bin_out_xhdl1_0_a2[5]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(7), B => wptr_gray_sync(6), C
         => wptr_gray_sync(5), D => wptr_bin_sync(8), Y => 
        wptr_bin_sync(5));
    
    \bin_out_xhdl1_0_a2[2]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(4), B => wptr_gray_sync(3), C
         => wptr_gray_sync(2), D => wptr_bin_sync(5), Y => 
        wptr_bin_sync(2));
    
    \bin_out_xhdl1_0_a2[0]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(2), B => wptr_bin_sync(3), C
         => wptr_gray_sync(0), D => wptr_gray_sync(1), Y => 
        wptr_bin_sync(0));
    
    \bin_out_xhdl1_i_o2[9]\ : CFG3
      generic map(INIT => x"96")

      port map(A => wptr_gray_sync(10), B => wptr_gray_sync(9), C
         => wptr_bin_sync(11), Y => wptr_bin_sync(9));
    
    \bin_out_xhdl1_i_o2[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => wptr_bin_sync(11), B => wptr_gray_sync(10), Y
         => wptr_bin_sync(10));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \bin_out_xhdl1_0_a2[6]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(8), B => wptr_gray_sync(7), C
         => wptr_gray_sync(6), D => wptr_bin_sync(9), Y => 
        wptr_bin_sync(6));
    
    \bin_out_xhdl1_0_a2[4]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(6), B => wptr_gray_sync(5), C
         => wptr_gray_sync(4), D => wptr_bin_sync(7), Y => 
        wptr_bin_sync(4));
    
    \bin_out_xhdl1_0_a2[8]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(10), B => wptr_gray_sync(9), C
         => wptr_gray_sync(8), D => wptr_bin_sync(11), Y => 
        wptr_bin_sync(8));
    
    \bin_out_xhdl1_0_a2[7]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(9), B => wptr_gray_sync(8), C
         => wptr_gray_sync(7), D => wptr_bin_sync(10), Y => 
        wptr_bin_sync(7));
    
    \bin_out_xhdl1_0_a2[3]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(5), B => wptr_gray_sync(4), C
         => wptr_gray_sync(3), D => wptr_bin_sync(6), Y => 
        wptr_bin_sync(3));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_1 is

    port( wptr_gray                 : in    std_logic_vector(11 downto 0);
          wptr_gray_sync            : out   std_logic_vector(10 downto 0);
          wptr_bin_sync_0           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          irx_fifo_rst_i            : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_1;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_1 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \sync_int[10]_net_1\, VCC_net_1, GND_net_1, 
        \sync_int[11]_net_1\, \sync_int[0]_net_1\, 
        \sync_int[1]_net_1\, \sync_int[2]_net_1\, 
        \sync_int[3]_net_1\, \sync_int[4]_net_1\, 
        \sync_int[5]_net_1\, \sync_int[6]_net_1\, 
        \sync_int[7]_net_1\, \sync_int[8]_net_1\, 
        \sync_int[9]_net_1\ : std_logic;

begin 


    \sync_int[9]\ : SLE
      port map(D => wptr_gray(9), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[9]_net_1\);
    
    \sync_int[4]\ : SLE
      port map(D => wptr_gray(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[4]_net_1\);
    
    \sync_out_xhdl1[10]\ : SLE
      port map(D => \sync_int[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(10));
    
    \sync_int[1]\ : SLE
      port map(D => wptr_gray(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[1]_net_1\);
    
    \sync_int[11]\ : SLE
      port map(D => wptr_gray(11), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[11]_net_1\);
    
    \sync_out_xhdl1[6]\ : SLE
      port map(D => \sync_int[6]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(6));
    
    \sync_out_xhdl1[3]\ : SLE
      port map(D => \sync_int[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(3));
    
    \sync_int[6]\ : SLE
      port map(D => wptr_gray(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[6]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \sync_out_xhdl1[11]\ : SLE
      port map(D => \sync_int[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_bin_sync_0);
    
    \sync_int[3]\ : SLE
      port map(D => wptr_gray(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[3]_net_1\);
    
    \sync_out_xhdl1[4]\ : SLE
      port map(D => \sync_int[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(4));
    
    \sync_int[0]\ : SLE
      port map(D => wptr_gray(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[0]_net_1\);
    
    \sync_out_xhdl1[1]\ : SLE
      port map(D => \sync_int[1]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(1));
    
    \sync_int[5]\ : SLE
      port map(D => wptr_gray(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[5]_net_1\);
    
    \sync_int[2]\ : SLE
      port map(D => wptr_gray(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[2]_net_1\);
    
    \sync_out_xhdl1[9]\ : SLE
      port map(D => \sync_int[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(9));
    
    \sync_out_xhdl1[2]\ : SLE
      port map(D => \sync_int[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(2));
    
    \sync_int[8]\ : SLE
      port map(D => wptr_gray(8), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[8]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sync_out_xhdl1[7]\ : SLE
      port map(D => \sync_int[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(7));
    
    \sync_out_xhdl1[5]\ : SLE
      port map(D => \sync_int[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(5));
    
    \sync_out_xhdl1[0]\ : SLE
      port map(D => \sync_int[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(0));
    
    \sync_out_xhdl1[8]\ : SLE
      port map(D => \sync_int[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(8));
    
    \sync_int[7]\ : SLE
      port map(D => wptr_gray(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[7]_net_1\);
    
    \sync_int[10]\ : SLE
      port map(D => wptr_gray(10), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_0 is

    port( rptr_gray           : in    std_logic_vector(11 downto 0);
          rptr_gray_sync      : out   std_logic_vector(10 downto 0);
          rptr_bin_sync_0     : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          irx_fifo_rst_i      : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_0;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_0 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \sync_int[4]_net_1\, GND_net_1, 
        \sync_int[5]_net_1\, \sync_int[6]_net_1\, 
        \sync_int[7]_net_1\, \sync_int[8]_net_1\, 
        \sync_int[9]_net_1\, \sync_int[10]_net_1\, 
        \sync_int[11]_net_1\, \sync_int[1]_net_1\, 
        \sync_int[2]_net_1\, \sync_int[3]_net_1\, 
        \sync_int[0]_net_1\ : std_logic;

begin 


    \sync_int[9]\ : SLE
      port map(D => rptr_gray(9), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[9]_net_1\);
    
    \sync_int[4]\ : SLE
      port map(D => rptr_gray(4), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[4]_net_1\);
    
    \sync_out_xhdl1[10]\ : SLE
      port map(D => \sync_int[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(10));
    
    \sync_int[1]\ : SLE
      port map(D => rptr_gray(1), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[1]_net_1\);
    
    \sync_int[11]\ : SLE
      port map(D => rptr_gray(11), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[11]_net_1\);
    
    \sync_out_xhdl1[6]\ : SLE
      port map(D => \sync_int[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(6));
    
    \sync_out_xhdl1[3]\ : SLE
      port map(D => \sync_int[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(3));
    
    \sync_int[6]\ : SLE
      port map(D => rptr_gray(6), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[6]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \sync_out_xhdl1[11]\ : SLE
      port map(D => \sync_int[11]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_bin_sync_0);
    
    \sync_int[3]\ : SLE
      port map(D => rptr_gray(3), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[3]_net_1\);
    
    \sync_out_xhdl1[4]\ : SLE
      port map(D => \sync_int[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(4));
    
    \sync_int[0]\ : SLE
      port map(D => rptr_gray(0), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[0]_net_1\);
    
    \sync_out_xhdl1[1]\ : SLE
      port map(D => \sync_int[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(1));
    
    \sync_int[5]\ : SLE
      port map(D => rptr_gray(5), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[5]_net_1\);
    
    \sync_int[2]\ : SLE
      port map(D => rptr_gray(2), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[2]_net_1\);
    
    \sync_out_xhdl1[9]\ : SLE
      port map(D => \sync_int[9]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(9));
    
    \sync_out_xhdl1[2]\ : SLE
      port map(D => \sync_int[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(2));
    
    \sync_int[8]\ : SLE
      port map(D => rptr_gray(8), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[8]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sync_out_xhdl1[7]\ : SLE
      port map(D => \sync_int[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(7));
    
    \sync_out_xhdl1[5]\ : SLE
      port map(D => \sync_int[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(5));
    
    \sync_out_xhdl1[0]\ : SLE
      port map(D => \sync_int[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(0));
    
    \sync_out_xhdl1[8]\ : SLE
      port map(D => \sync_int[8]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(8));
    
    \sync_int[7]\ : SLE
      port map(D => rptr_gray(7), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[7]_net_1\);
    
    \sync_int[10]\ : SLE
      port map(D => rptr_gray(10), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_1 is

    port( rptr_bin_sync  : inout std_logic_vector(11 downto 0) := (others => 'Z');
          rptr_gray_sync : in    std_logic_vector(10 downto 0)
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_1;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_1 is 

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    \bin_out_xhdl1_0_a2[1]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(1), B => rptr_gray_sync(2), C
         => rptr_bin_sync(3), Y => rptr_bin_sync(1));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \bin_out_xhdl1_0_a2[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(6), B => rptr_gray_sync(5), Y
         => rptr_bin_sync(5));
    
    \bin_out_xhdl1_0_a2[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(3), B => rptr_gray_sync(2), Y
         => rptr_bin_sync(2));
    
    \bin_out_xhdl1_0_a2[0]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(1), B => rptr_gray_sync(0), C
         => rptr_bin_sync(3), D => rptr_gray_sync(2), Y => 
        rptr_bin_sync(0));
    
    \bin_out_xhdl1_i_o2[9]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(9), B => rptr_gray_sync(10), C
         => rptr_bin_sync(11), Y => rptr_bin_sync(9));
    
    \bin_out_xhdl1_i_o2[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(11), B => rptr_gray_sync(10), Y
         => rptr_bin_sync(10));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \bin_out_xhdl1_0_a2[6]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(6), B => rptr_gray_sync(7), C
         => rptr_gray_sync(8), D => rptr_bin_sync(9), Y => 
        rptr_bin_sync(6));
    
    \bin_out_xhdl1_0_a2[4]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(5), B => rptr_bin_sync(6), C
         => rptr_gray_sync(4), Y => rptr_bin_sync(4));
    
    \bin_out_xhdl1_0_a2[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(9), B => rptr_gray_sync(8), Y
         => rptr_bin_sync(8));
    
    \bin_out_xhdl1_0_a2[7]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(8), B => rptr_bin_sync(9), C
         => rptr_gray_sync(7), Y => rptr_bin_sync(7));
    
    \bin_out_xhdl1_0_a2[3]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(5), B => rptr_bin_sync(6), C
         => rptr_gray_sync(3), D => rptr_gray_sync(4), Y => 
        rptr_bin_sync(3));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_0 is

    port( ReadFIFO_Write_Ptr        : in    std_logic_vector(1 downto 0);
          fifo_MEMWADDR             : out   std_logic_vector(10 downto 0);
          fifo_MEMRADDR             : out   std_logic_vector(10 downto 0);
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          N_152_i_i                 : out   std_logic;
          N_89_i                    : out   std_logic;
          REN_d1                    : in    std_logic;
          N_1003                    : in    std_logic;
          N_1466                    : in    std_logic;
          N_140_i                   : out   std_logic;
          fifo_MEMWE                : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          irx_fifo_rst_i            : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_0;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_0 is 

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_2
    port( wptr_bin_sync  : inout   std_logic_vector(11 downto 0);
          wptr_gray_sync : in    std_logic_vector(10 downto 0) := (others => 'U')
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_1
    port( wptr_gray                 : in    std_logic_vector(11 downto 0) := (others => 'U');
          wptr_gray_sync            : out   std_logic_vector(10 downto 0);
          wptr_bin_sync_0           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          irx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_0
    port( rptr_gray           : in    std_logic_vector(11 downto 0) := (others => 'U');
          rptr_gray_sync      : out   std_logic_vector(10 downto 0);
          rptr_bin_sync_0     : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          irx_fifo_rst_i      : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_1
    port( rptr_bin_sync  : inout   std_logic_vector(11 downto 0);
          rptr_gray_sync : in    std_logic_vector(10 downto 0) := (others => 'U')
        );
  end component;

    signal \rptr[0]_net_1\, \rptr_s[0]\, \fifo_MEMRADDR[0]\, 
        \memraddr_r_s[0]\, \wptr[0]_net_1\, \wptr_s[0]\, 
        \wptr_gray[10]_net_1\, VCC_net_1, \wptr_gray_1[10]_net_1\, 
        GND_net_1, \wptr_gray[11]_net_1\, \wptr[11]_net_1\, 
        \rptr_gray[0]_net_1\, \rptr_gray_1[0]_net_1\, 
        \rptr_gray[1]_net_1\, \rptr_gray_1[1]_net_1\, 
        \rptr_gray[2]_net_1\, \rptr_gray_1[2]_net_1\, 
        \rptr_gray[3]_net_1\, \rptr_gray_1[3]_net_1\, 
        \rptr_gray[4]_net_1\, \rptr_gray_1[4]_net_1\, 
        \rptr_gray[5]_net_1\, \rptr_gray_1[5]_net_1\, 
        \rptr_gray[6]_net_1\, \rptr_gray_1[6]_net_1\, 
        \rptr_gray[7]_net_1\, \rptr_gray_1[7]_net_1\, 
        \rptr_gray[8]_net_1\, \rptr_gray_1[8]_net_1\, 
        \rptr_gray[9]_net_1\, \rptr_gray_1[9]_net_1\, 
        \rptr_gray[10]_net_1\, \rptr_gray_1[10]_net_1\, 
        \rptr_gray[11]_net_1\, \rptr[11]_net_1\, 
        \wptr_bin_sync2[7]_net_1\, \wptr_bin_sync[7]\, 
        \wptr_bin_sync2[8]_net_1\, \wptr_bin_sync[8]\, 
        \wptr_bin_sync2[9]_net_1\, \wptr_bin_sync[9]\, 
        \wptr_bin_sync2[10]_net_1\, \wptr_bin_sync[10]\, 
        \wptr_bin_sync2[11]_net_1\, \wptr_bin_sync[11]\, 
        \wptr_gray[0]_net_1\, \wptr_gray_1[0]_net_1\, 
        \wptr_gray[1]_net_1\, \wptr_gray_1[1]_net_1\, 
        \wptr_gray[2]_net_1\, \wptr_gray_1[2]_net_1\, 
        \wptr_gray[3]_net_1\, \wptr_gray_1[3]_net_1\, 
        \wptr_gray[4]_net_1\, \wptr_gray_1[4]_net_1\, 
        \wptr_gray[5]_net_1\, \wptr_gray_1[5]_net_1\, 
        \wptr_gray[6]_net_1\, \wptr_gray_1[6]_net_1\, 
        \wptr_gray[7]_net_1\, \wptr_gray_1[7]_net_1\, 
        \wptr_gray[8]_net_1\, \wptr_gray_1[8]_net_1\, 
        \wptr_gray[9]_net_1\, \wptr_gray_1[9]_net_1\, rdiff_bus, 
        \wptr_bin_sync[0]\, \wptr_bin_sync2[1]_net_1\, 
        \wptr_bin_sync[1]\, \wptr_bin_sync2[2]_net_1\, 
        \wptr_bin_sync[2]\, \wptr_bin_sync2[3]_net_1\, 
        \wptr_bin_sync[3]\, \wptr_bin_sync2[4]_net_1\, 
        \wptr_bin_sync[4]\, \wptr_bin_sync2[5]_net_1\, 
        \wptr_bin_sync[5]\, \wptr_bin_sync2[6]_net_1\, 
        \wptr_bin_sync[6]\, \rptr_bin_sync2[7]_net_1\, 
        \rptr_bin_sync[7]\, \rptr_bin_sync2[8]_net_1\, 
        \rptr_bin_sync[8]\, \rptr_bin_sync2[9]_net_1\, 
        \rptr_bin_sync[9]\, \rptr_bin_sync2[10]_net_1\, 
        \rptr_bin_sync[10]\, \rptr_bin_sync2[11]_net_1\, 
        \rptr_bin_sync[11]\, un1_we_p, \rptr_bin_sync2[0]_net_1\, 
        \rptr_bin_sync[0]\, \rptr_bin_sync2[1]_net_1\, 
        \rptr_bin_sync[1]\, \rptr_bin_sync2[2]_net_1\, 
        \rptr_bin_sync[2]\, \rptr_bin_sync2[3]_net_1\, 
        \rptr_bin_sync[3]\, \rptr_bin_sync2[4]_net_1\, 
        \rptr_bin_sync[4]\, \rptr_bin_sync2[5]_net_1\, 
        \rptr_bin_sync[5]\, \rptr_bin_sync2[6]_net_1\, 
        \rptr_bin_sync[6]\, \iRX_FIFO_Full_0\, fulli, 
        un2_re_p_i_i_a3_0, \iRX_FIFO_Empty_0\, empty_r_3, 
        \fifo_MEMWE\, \wptr[1]_net_1\, \wptr_s[1]\, 
        \wptr[2]_net_1\, \wptr_s[2]\, \wptr[3]_net_1\, 
        \wptr_s[3]\, \wptr[4]_net_1\, \wptr_s[4]\, 
        \wptr[5]_net_1\, \wptr_s[5]\, \wptr[6]_net_1\, 
        \wptr_s[6]\, \wptr[7]_net_1\, \wptr_s[7]\, 
        \wptr[8]_net_1\, \wptr_s[8]\, \wptr[9]_net_1\, 
        \wptr_s[9]\, \wptr[10]_net_1\, \wptr_s[10]\, 
        \wptr_s[11]_net_1\, \N_140_i\, \fifo_MEMRADDR[1]\, 
        \memraddr_r_s[1]\, \fifo_MEMRADDR[2]\, \memraddr_r_s[2]\, 
        \fifo_MEMRADDR[3]\, \memraddr_r_s[3]\, \fifo_MEMRADDR[4]\, 
        \memraddr_r_s[4]\, \fifo_MEMRADDR[5]\, \memraddr_r_s[5]\, 
        \fifo_MEMRADDR[6]\, \memraddr_r_s[6]\, \fifo_MEMRADDR[7]\, 
        \memraddr_r_s[7]\, \fifo_MEMRADDR[8]\, \memraddr_r_s[8]\, 
        \fifo_MEMRADDR[9]\, \memraddr_r_s[9]\, 
        \fifo_MEMRADDR[10]\, \memraddr_r_s[10]_net_1\, 
        \fifo_MEMWADDR[0]\, \memwaddr_r_s[0]\, N_862, 
        \fifo_MEMWADDR[1]\, \memwaddr_r_s[1]\, \fifo_MEMWADDR[2]\, 
        \memwaddr_r_s[2]\, \fifo_MEMWADDR[3]\, \memwaddr_r_s[3]\, 
        \fifo_MEMWADDR[4]\, \memwaddr_r_s[4]\, \fifo_MEMWADDR[5]\, 
        \memwaddr_r_s[5]\, \fifo_MEMWADDR[6]\, \memwaddr_r_s[6]\, 
        \fifo_MEMWADDR[7]\, \memwaddr_r_s[7]\, \fifo_MEMWADDR[8]\, 
        \memwaddr_r_s[8]\, \fifo_MEMWADDR[9]\, \memwaddr_r_s[9]\, 
        \fifo_MEMWADDR[10]\, \memwaddr_r_s[10]_net_1\, 
        \rptr[1]_net_1\, \rptr_s[1]\, \rptr[2]_net_1\, 
        \rptr_s[2]\, \rptr[3]_net_1\, \rptr_s[3]\, 
        \rptr[4]_net_1\, \rptr_s[4]\, \rptr[5]_net_1\, 
        \rptr_s[5]\, \rptr[6]_net_1\, \rptr_s[6]\, 
        \rptr[7]_net_1\, \rptr_s[7]\, \rptr[8]_net_1\, 
        \rptr_s[8]\, \rptr[9]_net_1\, \rptr_s[9]\, 
        \rptr[10]_net_1\, \rptr_s[10]\, \rptr_s[11]_net_1\, 
        memwaddr_r_cry_cy, \memwaddr_r_cry[0]_net_1\, 
        \memwaddr_r_cry[1]_net_1\, \memwaddr_r_cry[2]_net_1\, 
        \memwaddr_r_cry[3]_net_1\, \memwaddr_r_cry[4]_net_1\, 
        \memwaddr_r_cry[5]_net_1\, \memwaddr_r_cry[6]_net_1\, 
        \memwaddr_r_cry[7]_net_1\, \memwaddr_r_cry[8]_net_1\, 
        \memwaddr_r_cry[9]_net_1\, \rdiff_bus_cry_0\, 
        rdiff_bus_cry_0_Y_1, \rdiff_bus_cry_1\, \rdiff_bus[1]\, 
        \rdiff_bus_cry_2\, \rdiff_bus[2]\, \rdiff_bus_cry_3\, 
        \rdiff_bus[3]\, \rdiff_bus_cry_4\, \rdiff_bus[4]\, 
        \rdiff_bus_cry_5\, \rdiff_bus[5]\, \rdiff_bus_cry_6\, 
        \rdiff_bus[6]\, \rdiff_bus_cry_7\, \rdiff_bus[7]\, 
        \rdiff_bus_cry_8\, \rdiff_bus[8]\, \rdiff_bus_cry_9\, 
        \rdiff_bus[9]\, \rdiff_bus[11]\, \rdiff_bus_cry_10\, 
        \rdiff_bus[10]\, \wdiff_bus_cry_0\, wdiff_bus_cry_0_Y_1, 
        \wdiff_bus_cry_1\, \wdiff_bus[1]\, \wdiff_bus_cry_2\, 
        \wdiff_bus[2]\, \wdiff_bus_cry_3\, \wdiff_bus[3]\, 
        \wdiff_bus_cry_4\, \wdiff_bus[4]\, \wdiff_bus_cry_5\, 
        \wdiff_bus[5]\, \wdiff_bus_cry_6\, \wdiff_bus[6]\, 
        \wdiff_bus_cry_7\, \wdiff_bus[7]\, \wdiff_bus_cry_8\, 
        \wdiff_bus[8]\, \wdiff_bus_cry_9\, \wdiff_bus[9]\, 
        \wdiff_bus[11]\, \wdiff_bus_cry_10\, \wdiff_bus[10]\, 
        rptr_s_380_FCO, \rptr_cry[1]_net_1\, \rptr_cry[2]_net_1\, 
        \rptr_cry[3]_net_1\, \rptr_cry[4]_net_1\, 
        \rptr_cry[5]_net_1\, \rptr_cry[6]_net_1\, 
        \rptr_cry[7]_net_1\, \rptr_cry[8]_net_1\, 
        \rptr_cry[9]_net_1\, \rptr_cry[10]_net_1\, 
        memraddr_r_s_381_FCO, \memraddr_r_cry[1]_net_1\, 
        \memraddr_r_cry[2]_net_1\, \memraddr_r_cry[3]_net_1\, 
        \memraddr_r_cry[4]_net_1\, \memraddr_r_cry[5]_net_1\, 
        \memraddr_r_cry[6]_net_1\, \memraddr_r_cry[7]_net_1\, 
        \memraddr_r_cry[8]_net_1\, \memraddr_r_cry[9]_net_1\, 
        wptr_s_382_FCO, \wptr_cry[1]_net_1\, \wptr_cry[2]_net_1\, 
        \wptr_cry[3]_net_1\, \wptr_cry[4]_net_1\, 
        \wptr_cry[5]_net_1\, \wptr_cry[6]_net_1\, 
        \wptr_cry[7]_net_1\, \wptr_cry[8]_net_1\, 
        \wptr_cry[9]_net_1\, \wptr_cry[10]_net_1\, 
        empty_r_3_0_a2_1, \fulli_0_a2_7\, \fulli_0_a2_6\, 
        empty_r_3_0_a2_7, empty_r_3_0_a2_9, \fulli_0_a2_8\, 
        empty_r_3_0_a2_5, \wptr_gray_sync[0]\, 
        \wptr_gray_sync[1]\, \wptr_gray_sync[2]\, 
        \wptr_gray_sync[3]\, \wptr_gray_sync[4]\, 
        \wptr_gray_sync[5]\, \wptr_gray_sync[6]\, 
        \wptr_gray_sync[7]\, \wptr_gray_sync[8]\, 
        \wptr_gray_sync[9]\, \wptr_gray_sync[10]\, 
        \rptr_gray_sync[0]\, \rptr_gray_sync[1]\, 
        \rptr_gray_sync[2]\, \rptr_gray_sync[3]\, 
        \rptr_gray_sync[4]\, \rptr_gray_sync[5]\, 
        \rptr_gray_sync[6]\, \rptr_gray_sync[7]\, 
        \rptr_gray_sync[8]\, \rptr_gray_sync[9]\, 
        \rptr_gray_sync[10]\ : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_2
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_2(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_1
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_1(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_0
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_0(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_1
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_1(DEF_ARCH);
begin 

    fifo_MEMWADDR(10) <= \fifo_MEMWADDR[10]\;
    fifo_MEMWADDR(9) <= \fifo_MEMWADDR[9]\;
    fifo_MEMWADDR(8) <= \fifo_MEMWADDR[8]\;
    fifo_MEMWADDR(7) <= \fifo_MEMWADDR[7]\;
    fifo_MEMWADDR(6) <= \fifo_MEMWADDR[6]\;
    fifo_MEMWADDR(5) <= \fifo_MEMWADDR[5]\;
    fifo_MEMWADDR(4) <= \fifo_MEMWADDR[4]\;
    fifo_MEMWADDR(3) <= \fifo_MEMWADDR[3]\;
    fifo_MEMWADDR(2) <= \fifo_MEMWADDR[2]\;
    fifo_MEMWADDR(1) <= \fifo_MEMWADDR[1]\;
    fifo_MEMWADDR(0) <= \fifo_MEMWADDR[0]\;
    fifo_MEMRADDR(10) <= \fifo_MEMRADDR[10]\;
    fifo_MEMRADDR(9) <= \fifo_MEMRADDR[9]\;
    fifo_MEMRADDR(8) <= \fifo_MEMRADDR[8]\;
    fifo_MEMRADDR(7) <= \fifo_MEMRADDR[7]\;
    fifo_MEMRADDR(6) <= \fifo_MEMRADDR[6]\;
    fifo_MEMRADDR(5) <= \fifo_MEMRADDR[5]\;
    fifo_MEMRADDR(4) <= \fifo_MEMRADDR[4]\;
    fifo_MEMRADDR(3) <= \fifo_MEMRADDR[3]\;
    fifo_MEMRADDR(2) <= \fifo_MEMRADDR[2]\;
    fifo_MEMRADDR(1) <= \fifo_MEMRADDR[1]\;
    fifo_MEMRADDR(0) <= \fifo_MEMRADDR[0]\;
    iRX_FIFO_Empty_0 <= \iRX_FIFO_Empty_0\;
    iRX_FIFO_Full_0 <= \iRX_FIFO_Full_0\;
    N_140_i <= \N_140_i\;
    fifo_MEMWE <= \fifo_MEMWE\;

    \rptr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[4]_net_1\, S
         => \rptr_s[5]\, Y => OPEN, FCO => \rptr_cry[5]_net_1\);
    
    wdiff_bus_cry_8 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[8]_net_1\, B => 
        \rptr_bin_sync2[8]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_7\, S => \wdiff_bus[8]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_8\);
    
    \wptr_gray[4]\ : SLE
      port map(D => \wptr_gray_1[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[4]_net_1\);
    
    \rptr_gray_1[3]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[3]_net_1\, B => \rptr[4]_net_1\, Y => 
        \rptr_gray_1[3]_net_1\);
    
    \rptr_bin_sync2[6]\ : SLE
      port map(D => \rptr_bin_sync[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[6]_net_1\);
    
    fulli_0_a2_0_0_a2 : CFG3
      generic map(INIT => x"08")

      port map(A => ReadFIFO_Write_Ptr(0), B => N_1466, C => 
        ReadFIFO_Write_Ptr(1), Y => N_862);
    
    \rptr[1]\ : SLE
      port map(D => \rptr_s[1]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_140_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[1]_net_1\);
    
    \wptr_gray_1[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[9]_net_1\, B => \wptr[10]_net_1\, Y => 
        \wptr_gray_1[9]_net_1\);
    
    \rptr_gray_1[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[5]_net_1\, B => \rptr[6]_net_1\, Y => 
        \rptr_gray_1[5]_net_1\);
    
    \rptr_gray[9]\ : SLE
      port map(D => \rptr_gray_1[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[9]_net_1\);
    
    \rptr_gray[8]\ : SLE
      port map(D => \rptr_gray_1[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[8]_net_1\);
    
    \rptr_gray_1[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[2]_net_1\, B => \rptr[3]_net_1\, Y => 
        \rptr_gray_1[2]_net_1\);
    
    \rptr_bin_sync2[7]\ : SLE
      port map(D => \rptr_bin_sync[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[7]_net_1\);
    
    \memwaddr_r[1]\ : SLE
      port map(D => \memwaddr_r_s[1]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_862, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[1]\);
    
    \memwaddr_r_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[5]_net_1\, S => \memwaddr_r_s[6]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[6]_net_1\);
    
    \memwaddr_r_s[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[9]_net_1\, S => \memwaddr_r_s[10]_net_1\, 
        Y => OPEN, FCO => OPEN);
    
    \wptr_gray_1[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[7]_net_1\, B => \wptr[8]_net_1\, Y => 
        \wptr_gray_1[7]_net_1\);
    
    \memraddr_r[0]\ : SLE
      port map(D => \memraddr_r_s[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_140_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[0]\);
    
    \wptr[0]\ : SLE
      port map(D => \wptr_s[0]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[0]_net_1\);
    
    \rptr_bin_sync2[8]\ : SLE
      port map(D => \rptr_bin_sync[8]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[8]_net_1\);
    
    \rptr_gray_1[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[1]_net_1\, B => \rptr[2]_net_1\, Y => 
        \rptr_gray_1[1]_net_1\);
    
    \rptr_gray[10]\ : SLE
      port map(D => \rptr_gray_1[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[10]_net_1\);
    
    \wptr_gray_1[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[0]_net_1\, B => \wptr[1]_net_1\, Y => 
        \wptr_gray_1[0]_net_1\);
    
    wdiff_bus_cry_9 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[9]_net_1\, B => 
        \rptr_bin_sync2[9]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_8\, S => \wdiff_bus[9]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_9\);
    
    \rptr[5]\ : SLE
      port map(D => \rptr_s[5]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_140_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[5]_net_1\);
    
    \rptr_gray[3]\ : SLE
      port map(D => \rptr_gray_1[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[3]_net_1\);
    
    \rptr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[5]_net_1\, S
         => \rptr_s[6]\, Y => OPEN, FCO => \rptr_cry[6]_net_1\);
    
    \memwaddr_r_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[1]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[0]_net_1\, S => \memwaddr_r_s[1]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[1]_net_1\);
    
    fulli_0_a2_6 : CFG4
      generic map(INIT => x"8000")

      port map(A => \wdiff_bus[2]\, B => \wdiff_bus[3]\, C => 
        \wdiff_bus[5]\, D => \wdiff_bus[4]\, Y => \fulli_0_a2_6\);
    
    \wptr_gray[3]\ : SLE
      port map(D => \wptr_gray_1[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[3]_net_1\);
    
    \rptr_gray_1[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[11]_net_1\, B => \rptr[10]_net_1\, Y
         => \rptr_gray_1[10]_net_1\);
    
    wdiff_bus_s_11 : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \rptr_bin_sync2[11]_net_1\, C
         => \wptr[11]_net_1\, D => GND_net_1, FCI => 
        \wdiff_bus_cry_10\, S => \wdiff_bus[11]\, Y => OPEN, FCO
         => OPEN);
    
    \rptr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[7]_net_1\, S
         => \rptr_s[8]\, Y => OPEN, FCO => \rptr_cry[8]_net_1\);
    
    \rptr[7]\ : SLE
      port map(D => \rptr_s[7]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_140_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[7]_net_1\);
    
    rdiff_bus_cry_4 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[4]_net_1\, B => 
        \rptr[4]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_3\, S => \rdiff_bus[4]\, Y => OPEN, FCO
         => \rdiff_bus_cry_4\);
    
    \rptr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[9]_net_1\, S
         => \rptr_s[10]\, Y => OPEN, FCO => \rptr_cry[10]_net_1\);
    
    \rptr_bin_sync2[0]\ : SLE
      port map(D => \rptr_bin_sync[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[0]_net_1\);
    
    \L1.empty_r_3_0_a2_7\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \rdiff_bus[5]\, B => \rdiff_bus[6]\, C => 
        \rdiff_bus[7]\, D => \rdiff_bus[8]\, Y => 
        empty_r_3_0_a2_7);
    
    \wptr[11]\ : SLE
      port map(D => \wptr_s[11]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \wptr[11]_net_1\);
    
    rdiff_bus_cry_1 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[1]_net_1\, B => 
        \rptr[1]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_0\, S => \rdiff_bus[1]\, Y => OPEN, FCO
         => \rdiff_bus_cry_1\);
    
    \memraddr_r[1]\ : SLE
      port map(D => \memraddr_r_s[1]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_140_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[1]\);
    
    \L1.empty_r_3_0_a2_9\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \rdiff_bus[1]\, B => \rdiff_bus[2]\, C => 
        empty_r_3_0_a2_7, D => empty_r_3_0_a2_1, Y => 
        empty_r_3_0_a2_9);
    
    \rptr_bin_sync2[2]\ : SLE
      port map(D => \rptr_bin_sync[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[2]_net_1\);
    
    rdiff_bus_cry_6 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[6]_net_1\, B => 
        \rptr[6]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_5\, S => \rdiff_bus[6]\, Y => OPEN, FCO
         => \rdiff_bus_cry_6\);
    
    memraddr_r_s_381 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[0]\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => memraddr_r_s_381_FCO);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \memwaddr_r_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[3]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[2]_net_1\, S => \memwaddr_r_s[3]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[3]_net_1\);
    
    \rptr_gray[1]\ : SLE
      port map(D => \rptr_gray_1[1]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[1]_net_1\);
    
    \memwaddr_r[7]\ : SLE
      port map(D => \memwaddr_r_s[7]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_862, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[7]\);
    
    \memraddr_r_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[2]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[1]_net_1\, S => \memraddr_r_s[2]\, Y => 
        OPEN, FCO => \memraddr_r_cry[2]_net_1\);
    
    \wptr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[3]_net_1\, S
         => \wptr_s[4]\, Y => OPEN, FCO => \wptr_cry[4]_net_1\);
    
    empty_r_RNI0OFF1 : CFG3
      generic map(INIT => x"A6")

      port map(A => REN_d1, B => N_1003, C => \iRX_FIFO_Empty_0\, 
        Y => N_152_i_i);
    
    \memraddr_r_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[8]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[7]_net_1\, S => \memraddr_r_s[8]\, Y => 
        OPEN, FCO => \memraddr_r_cry[8]_net_1\);
    
    \wptr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[9]_net_1\, S
         => \wptr_s[10]\, Y => OPEN, FCO => \wptr_cry[10]_net_1\);
    
    wdiff_bus_cry_5 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[5]_net_1\, B => 
        \rptr_bin_sync2[5]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_4\, S => \wdiff_bus[5]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_5\);
    
    \memwaddr_r[4]\ : SLE
      port map(D => \memwaddr_r_s[4]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_862, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[4]\);
    
    \wptr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[1]_net_1\, S
         => \wptr_s[2]\, Y => OPEN, FCO => \wptr_cry[2]_net_1\);
    
    wdiff_bus_cry_0 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[0]_net_1\, B => 
        \rptr_bin_sync2[0]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => VCC_net_1, S => OPEN, Y => wdiff_bus_cry_0_Y_1, 
        FCO => \wdiff_bus_cry_0\);
    
    \wptr[1]\ : SLE
      port map(D => \wptr_s[1]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[1]_net_1\);
    
    \rptr_bin_sync2[4]\ : SLE
      port map(D => \rptr_bin_sync[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[4]_net_1\);
    
    \wptr_bin_sync2[6]\ : SLE
      port map(D => \wptr_bin_sync[6]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[6]_net_1\);
    
    \memwaddr_r_cry_cy[0]\ : ARI1
      generic map(INIT => x"45500")

      port map(A => VCC_net_1, B => \iRX_FIFO_Full_0\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => memwaddr_r_cry_cy);
    
    \rptr[3]\ : SLE
      port map(D => \rptr_s[3]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_140_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[3]_net_1\);
    
    \wptr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[2]_net_1\, S
         => \wptr_s[3]\, Y => OPEN, FCO => \wptr_cry[3]_net_1\);
    
    \memwaddr_r_cry[0]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[0]\, C => 
        GND_net_1, D => GND_net_1, FCI => memwaddr_r_cry_cy, S
         => \memwaddr_r_s[0]\, Y => OPEN, FCO => 
        \memwaddr_r_cry[0]_net_1\);
    
    \rptr[6]\ : SLE
      port map(D => \rptr_s[6]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_140_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[6]_net_1\);
    
    rdiff_bus_cry_8 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[8]_net_1\, B => 
        \rptr[8]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_7\, S => \rdiff_bus[8]\, Y => OPEN, FCO
         => \rdiff_bus_cry_8\);
    
    \wptr_gray[10]\ : SLE
      port map(D => \wptr_gray_1[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[10]_net_1\);
    
    rdiff_bus_cry_7 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[7]_net_1\, B => 
        \rptr[7]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_6\, S => \rdiff_bus[7]\, Y => OPEN, FCO
         => \rdiff_bus_cry_7\);
    
    \wptr_bin_sync2[7]\ : SLE
      port map(D => \wptr_bin_sync[7]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[7]_net_1\);
    
    \rptr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[8]_net_1\, S
         => \rptr_s[9]\, Y => OPEN, FCO => \rptr_cry[9]_net_1\);
    
    \rptr_gray[5]\ : SLE
      port map(D => \rptr_gray_1[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[5]_net_1\);
    
    \wptr_gray_1[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[2]_net_1\, B => \wptr[3]_net_1\, Y => 
        \wptr_gray_1[2]_net_1\);
    
    \wptr[5]\ : SLE
      port map(D => \wptr_s[5]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[5]_net_1\);
    
    rdiff_bus_cry_5 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[5]_net_1\, B => 
        \rptr[5]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_4\, S => \rdiff_bus[5]\, Y => OPEN, FCO
         => \rdiff_bus_cry_5\);
    
    \wptr_bin_sync2[8]\ : SLE
      port map(D => \wptr_bin_sync[8]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[8]_net_1\);
    
    \wptr[7]\ : SLE
      port map(D => \wptr_s[7]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[7]_net_1\);
    
    empty_r_RNI0OFF1_0 : CFG3
      generic map(INIT => x"A2")

      port map(A => REN_d1, B => N_1003, C => \iRX_FIFO_Empty_0\, 
        Y => N_89_i);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \wptr_gray[1]\ : SLE
      port map(D => \wptr_gray_1[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[1]_net_1\);
    
    \rptr_gray_1[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[9]_net_1\, B => \rptr[10]_net_1\, Y => 
        \rptr_gray_1[9]_net_1\);
    
    \rptr_bin_sync2[5]\ : SLE
      port map(D => \rptr_bin_sync[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[5]_net_1\);
    
    \rptr_bin_sync2[1]\ : SLE
      port map(D => \rptr_bin_sync[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[1]_net_1\);
    
    \memwaddr_r[10]\ : SLE
      port map(D => \memwaddr_r_s[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_862, ALn => irx_fifo_rst_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \fifo_MEMWADDR[10]\);
    
    wdiff_bus_cry_7 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[7]_net_1\, B => 
        \rptr_bin_sync2[7]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_6\, S => \wdiff_bus[7]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_7\);
    
    \wptr_bin_sync2[0]\ : SLE
      port map(D => \wptr_bin_sync[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rdiff_bus);
    
    \L1.un2_re_p_i_i_a3\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1003, B => \iRX_FIFO_Empty_0\, Y => 
        un2_re_p_i_i_a3_0);
    
    \L1.empty_r_3_0_a2_1\ : CFG2
      generic map(INIT => x"1")

      port map(A => \rdiff_bus[4]\, B => \rdiff_bus[3]\, Y => 
        empty_r_3_0_a2_1);
    
    \L1.un1_we_p_0_a2_0_a2\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_862, B => \iRX_FIFO_Full_0\, Y => un1_we_p);
    
    rdiff_bus_s_11 : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \rptr[11]_net_1\, C => 
        \wptr_bin_sync2[11]_net_1\, D => GND_net_1, FCI => 
        \rdiff_bus_cry_10\, S => \rdiff_bus[11]\, Y => OPEN, FCO
         => OPEN);
    
    \memwaddr_r_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[8]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[7]_net_1\, S => \memwaddr_r_s[8]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[8]_net_1\);
    
    \wptr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => wptr_s_382_FCO, S => 
        \wptr_s[1]\, Y => OPEN, FCO => \wptr_cry[1]_net_1\);
    
    \memraddr_r[8]\ : SLE
      port map(D => \memraddr_r_s[8]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_140_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[8]\);
    
    \rptr[9]\ : SLE
      port map(D => \rptr_s[9]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_140_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[9]_net_1\);
    
    \wptr_gray_1[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[6]_net_1\, B => \wptr[7]_net_1\, Y => 
        \wptr_gray_1[6]_net_1\);
    
    \wptr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[6]_net_1\, S
         => \wptr_s[7]\, Y => OPEN, FCO => \wptr_cry[7]_net_1\);
    
    \wptr_bin_sync2[2]\ : SLE
      port map(D => \wptr_bin_sync[2]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[2]_net_1\);
    
    \rptr_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \rptr[0]_net_1\, Y => \rptr_s[0]\);
    
    \rptr[4]\ : SLE
      port map(D => \rptr_s[4]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_140_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[4]_net_1\);
    
    \memwaddr_r_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[4]_net_1\, S => \memwaddr_r_s[5]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[5]_net_1\);
    
    \memraddr_r_s[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[9]_net_1\, S => \memraddr_r_s[10]_net_1\, 
        Y => OPEN, FCO => OPEN);
    
    \wptr_gray[6]\ : SLE
      port map(D => \wptr_gray_1[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[6]_net_1\);
    
    \wptr_gray_1[3]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[3]_net_1\, B => \wptr[4]_net_1\, Y => 
        \wptr_gray_1[3]_net_1\);
    
    \wptr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[4]_net_1\, S
         => \wptr_s[5]\, Y => OPEN, FCO => \wptr_cry[5]_net_1\);
    
    \memraddr_r_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[4]_net_1\, S => \memraddr_r_s[5]\, Y => 
        OPEN, FCO => \memraddr_r_cry[5]_net_1\);
    
    \memraddr_r_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[1]\, C => 
        GND_net_1, D => GND_net_1, FCI => memraddr_r_s_381_FCO, S
         => \memraddr_r_s[1]\, Y => OPEN, FCO => 
        \memraddr_r_cry[1]_net_1\);
    
    \rptr_gray[4]\ : SLE
      port map(D => \rptr_gray_1[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[4]_net_1\);
    
    \wptr_bin_sync2[4]\ : SLE
      port map(D => \wptr_bin_sync[4]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[4]_net_1\);
    
    \wptr[3]\ : SLE
      port map(D => \wptr_s[3]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[3]_net_1\);
    
    \memwaddr_r[6]\ : SLE
      port map(D => \memwaddr_r_s[6]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_862, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[6]\);
    
    \wptr_s[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[10]_net_1\, S
         => \wptr_s[11]_net_1\, Y => OPEN, FCO => OPEN);
    
    \wptr[6]\ : SLE
      port map(D => \wptr_s[6]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[6]_net_1\);
    
    rptr_s_380 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => rptr_s_380_FCO);
    
    \memwaddr_r[9]\ : SLE
      port map(D => \memwaddr_r_s[9]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_862, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[9]\);
    
    \memraddr_r_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[3]_net_1\, S => \memraddr_r_s[4]\, Y => 
        OPEN, FCO => \memraddr_r_cry[4]_net_1\);
    
    \memraddr_r[10]\ : SLE
      port map(D => \memraddr_r_s[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_140_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[10]\);
    
    \memwaddr_r[3]\ : SLE
      port map(D => \memwaddr_r_s[3]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_862, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[3]\);
    
    full_r : SLE
      port map(D => fulli, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \iRX_FIFO_Full_0\);
    
    \rptr_bin_sync2[3]\ : SLE
      port map(D => \rptr_bin_sync[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[3]_net_1\);
    
    \wptr_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \wptr[0]_net_1\, Y => \wptr_s[0]\);
    
    \rptr[2]\ : SLE
      port map(D => \rptr_s[2]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_140_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[2]_net_1\);
    
    \memraddr_r[3]\ : SLE
      port map(D => \memraddr_r_s[3]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_140_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[3]\);
    
    \rptr_bin_sync2[9]\ : SLE
      port map(D => \rptr_bin_sync[9]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[9]_net_1\);
    
    empty_r_RNI15131 : CFG2
      generic map(INIT => x"2")

      port map(A => N_1003, B => \iRX_FIFO_Empty_0\, Y => 
        \N_140_i\);
    
    \rptr[11]\ : SLE
      port map(D => \rptr_s[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_140_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rptr[11]_net_1\);
    
    \wptr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[5]_net_1\, S
         => \wptr_s[6]\, Y => OPEN, FCO => \wptr_cry[6]_net_1\);
    
    \rptr_bin_sync2[11]\ : SLE
      port map(D => \rptr_bin_sync[11]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[11]_net_1\);
    
    \wptr_bin_sync2[5]\ : SLE
      port map(D => \wptr_bin_sync[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[5]_net_1\);
    
    \wptr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[7]_net_1\, S
         => \wptr_s[8]\, Y => OPEN, FCO => \wptr_cry[8]_net_1\);
    
    \wptr_bin_sync2[1]\ : SLE
      port map(D => \wptr_bin_sync[1]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[1]_net_1\);
    
    Wr_corefifo_grayToBinConv : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_2
      port map(wptr_bin_sync(11) => \wptr_bin_sync[11]\, 
        wptr_bin_sync(10) => \wptr_bin_sync[10]\, 
        wptr_bin_sync(9) => \wptr_bin_sync[9]\, wptr_bin_sync(8)
         => \wptr_bin_sync[8]\, wptr_bin_sync(7) => 
        \wptr_bin_sync[7]\, wptr_bin_sync(6) => 
        \wptr_bin_sync[6]\, wptr_bin_sync(5) => 
        \wptr_bin_sync[5]\, wptr_bin_sync(4) => 
        \wptr_bin_sync[4]\, wptr_bin_sync(3) => 
        \wptr_bin_sync[3]\, wptr_bin_sync(2) => 
        \wptr_bin_sync[2]\, wptr_bin_sync(1) => 
        \wptr_bin_sync[1]\, wptr_bin_sync(0) => 
        \wptr_bin_sync[0]\, wptr_gray_sync(10) => 
        \wptr_gray_sync[10]\, wptr_gray_sync(9) => 
        \wptr_gray_sync[9]\, wptr_gray_sync(8) => 
        \wptr_gray_sync[8]\, wptr_gray_sync(7) => 
        \wptr_gray_sync[7]\, wptr_gray_sync(6) => 
        \wptr_gray_sync[6]\, wptr_gray_sync(5) => 
        \wptr_gray_sync[5]\, wptr_gray_sync(4) => 
        \wptr_gray_sync[4]\, wptr_gray_sync(3) => 
        \wptr_gray_sync[3]\, wptr_gray_sync(2) => 
        \wptr_gray_sync[2]\, wptr_gray_sync(1) => 
        \wptr_gray_sync[1]\, wptr_gray_sync(0) => 
        \wptr_gray_sync[0]\);
    
    \wptr_gray_1[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[4]_net_1\, B => \wptr[5]_net_1\, Y => 
        \wptr_gray_1[4]_net_1\);
    
    overflow_r : SLE
      port map(D => un1_we_p, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        iRX_FIFO_OVERFLOW_0);
    
    fulli_0 : CFG4
      generic map(INIT => x"EAAA")

      port map(A => \wdiff_bus[11]\, B => \fulli_0_a2_7\, C => 
        N_862, D => \fulli_0_a2_8\, Y => fulli);
    
    \memraddr_r_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \fifo_MEMRADDR[0]\, Y => \memraddr_r_s[0]\);
    
    \rptr_gray[11]\ : SLE
      port map(D => \rptr[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[11]_net_1\);
    
    \wptr_bin_sync2[10]\ : SLE
      port map(D => \wptr_bin_sync[10]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[10]_net_1\);
    
    \rptr[10]\ : SLE
      port map(D => \rptr_s[10]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_140_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rptr[10]_net_1\);
    
    \wptr[9]\ : SLE
      port map(D => \wptr_s[9]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[9]_net_1\);
    
    Wr_corefifo_doubleSync : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_1
      port map(wptr_gray(11) => \wptr_gray[11]_net_1\, 
        wptr_gray(10) => \wptr_gray[10]_net_1\, wptr_gray(9) => 
        \wptr_gray[9]_net_1\, wptr_gray(8) => 
        \wptr_gray[8]_net_1\, wptr_gray(7) => 
        \wptr_gray[7]_net_1\, wptr_gray(6) => 
        \wptr_gray[6]_net_1\, wptr_gray(5) => 
        \wptr_gray[5]_net_1\, wptr_gray(4) => 
        \wptr_gray[4]_net_1\, wptr_gray(3) => 
        \wptr_gray[3]_net_1\, wptr_gray(2) => 
        \wptr_gray[2]_net_1\, wptr_gray(1) => 
        \wptr_gray[1]_net_1\, wptr_gray(0) => 
        \wptr_gray[0]_net_1\, wptr_gray_sync(10) => 
        \wptr_gray_sync[10]\, wptr_gray_sync(9) => 
        \wptr_gray_sync[9]\, wptr_gray_sync(8) => 
        \wptr_gray_sync[8]\, wptr_gray_sync(7) => 
        \wptr_gray_sync[7]\, wptr_gray_sync(6) => 
        \wptr_gray_sync[6]\, wptr_gray_sync(5) => 
        \wptr_gray_sync[5]\, wptr_gray_sync(4) => 
        \wptr_gray_sync[4]\, wptr_gray_sync(3) => 
        \wptr_gray_sync[3]\, wptr_gray_sync(2) => 
        \wptr_gray_sync[2]\, wptr_gray_sync(1) => 
        \wptr_gray_sync[1]\, wptr_gray_sync(0) => 
        \wptr_gray_sync[0]\, wptr_bin_sync_0 => 
        \wptr_bin_sync[11]\, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, irx_fifo_rst_i => 
        irx_fifo_rst_i);
    
    \rptr_gray[0]\ : SLE
      port map(D => \rptr_gray_1[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[0]_net_1\);
    
    empty_r : SLE
      port map(D => empty_r_3, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \iRX_FIFO_Empty_0\);
    
    \rptr_gray_1[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[7]_net_1\, B => \rptr[8]_net_1\, Y => 
        \rptr_gray_1[7]_net_1\);
    
    \wptr[4]\ : SLE
      port map(D => \wptr_s[4]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[4]_net_1\);
    
    \memwaddr_r[8]\ : SLE
      port map(D => \memwaddr_r_s[8]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_862, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[8]\);
    
    \memwaddr_r[2]\ : SLE
      port map(D => \memwaddr_r_s[2]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_862, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[2]\);
    
    \L1.empty_r_3_0_a2_5\ : CFG3
      generic map(INIT => x"0E")

      port map(A => N_1003, B => rdiff_bus_cry_0_Y_1, C => 
        \rdiff_bus[11]\, Y => empty_r_3_0_a2_5);
    
    \wptr_bin_sync2[11]\ : SLE
      port map(D => \wptr_bin_sync[11]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[11]_net_1\);
    
    \wptr_gray_1[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[1]_net_1\, B => \wptr[2]_net_1\, Y => 
        \wptr_gray_1[1]_net_1\);
    
    underflow_r : SLE
      port map(D => un2_re_p_i_i_a3_0, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => iRX_FIFO_UNDERRUN_0);
    
    \memwaddr_r_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[6]_net_1\, S => \memwaddr_r_s[7]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[7]_net_1\);
    
    \wptr_gray[5]\ : SLE
      port map(D => \wptr_gray_1[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[5]_net_1\);
    
    \memraddr_r[7]\ : SLE
      port map(D => \memraddr_r_s[7]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_140_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[7]\);
    
    memwe_0_a2_0_a2 : CFG4
      generic map(INIT => x"1000")

      port map(A => ReadFIFO_Write_Ptr(1), B => \iRX_FIFO_Full_0\, 
        C => N_1466, D => ReadFIFO_Write_Ptr(0), Y => 
        \fifo_MEMWE\);
    
    \rptr_bin_sync2[10]\ : SLE
      port map(D => \rptr_bin_sync[10]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[10]_net_1\);
    
    wdiff_bus_cry_10 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[10]_net_1\, B => 
        \rptr_bin_sync2[10]_net_1\, C => GND_net_1, D => 
        GND_net_1, FCI => \wdiff_bus_cry_9\, S => \wdiff_bus[10]\, 
        Y => OPEN, FCO => \wdiff_bus_cry_10\);
    
    \memwaddr_r_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[9]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[8]_net_1\, S => \memwaddr_r_s[9]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[9]_net_1\);
    
    \wptr_gray[8]\ : SLE
      port map(D => \wptr_gray_1[8]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[8]_net_1\);
    
    \wptr_gray[7]\ : SLE
      port map(D => \wptr_gray_1[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[7]_net_1\);
    
    \wptr_gray_1[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[5]_net_1\, B => \wptr[6]_net_1\, Y => 
        \wptr_gray_1[5]_net_1\);
    
    \memwaddr_r[5]\ : SLE
      port map(D => \memwaddr_r_s[5]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_862, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[5]\);
    
    \L1.empty_r_3_0_a2\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \rdiff_bus[9]\, B => \rdiff_bus[10]\, C => 
        empty_r_3_0_a2_5, D => empty_r_3_0_a2_9, Y => empty_r_3);
    
    \rptr[8]\ : SLE
      port map(D => \rptr_s[8]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_140_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[8]_net_1\);
    
    Rd_corefifo_doubleSync : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_0
      port map(rptr_gray(11) => \rptr_gray[11]_net_1\, 
        rptr_gray(10) => \rptr_gray[10]_net_1\, rptr_gray(9) => 
        \rptr_gray[9]_net_1\, rptr_gray(8) => 
        \rptr_gray[8]_net_1\, rptr_gray(7) => 
        \rptr_gray[7]_net_1\, rptr_gray(6) => 
        \rptr_gray[6]_net_1\, rptr_gray(5) => 
        \rptr_gray[5]_net_1\, rptr_gray(4) => 
        \rptr_gray[4]_net_1\, rptr_gray(3) => 
        \rptr_gray[3]_net_1\, rptr_gray(2) => 
        \rptr_gray[2]_net_1\, rptr_gray(1) => 
        \rptr_gray[1]_net_1\, rptr_gray(0) => 
        \rptr_gray[0]_net_1\, rptr_gray_sync(10) => 
        \rptr_gray_sync[10]\, rptr_gray_sync(9) => 
        \rptr_gray_sync[9]\, rptr_gray_sync(8) => 
        \rptr_gray_sync[8]\, rptr_gray_sync(7) => 
        \rptr_gray_sync[7]\, rptr_gray_sync(6) => 
        \rptr_gray_sync[6]\, rptr_gray_sync(5) => 
        \rptr_gray_sync[5]\, rptr_gray_sync(4) => 
        \rptr_gray_sync[4]\, rptr_gray_sync(3) => 
        \rptr_gray_sync[3]\, rptr_gray_sync(2) => 
        \rptr_gray_sync[2]\, rptr_gray_sync(1) => 
        \rptr_gray_sync[1]\, rptr_gray_sync(0) => 
        \rptr_gray_sync[0]\, rptr_bin_sync_0 => 
        \rptr_bin_sync[11]\, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, irx_fifo_rst_i => irx_fifo_rst_i);
    
    \rptr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[3]_net_1\, S
         => \rptr_s[4]\, Y => OPEN, FCO => \rptr_cry[4]_net_1\);
    
    wdiff_bus_cry_2 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[2]_net_1\, B => 
        \rptr_bin_sync2[2]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_1\, S => \wdiff_bus[2]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_2\);
    
    \rptr_gray[2]\ : SLE
      port map(D => \rptr_gray_1[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[2]_net_1\);
    
    \wptr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[8]_net_1\, S
         => \wptr_s[9]\, Y => OPEN, FCO => \wptr_cry[9]_net_1\);
    
    \wptr_bin_sync2[3]\ : SLE
      port map(D => \wptr_bin_sync[3]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[3]_net_1\);
    
    \wptr[2]\ : SLE
      port map(D => \wptr_s[2]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[2]_net_1\);
    
    \rptr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[1]_net_1\, S
         => \rptr_s[2]\, Y => OPEN, FCO => \rptr_cry[2]_net_1\);
    
    rdiff_bus_cry_9 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[9]_net_1\, B => 
        \rptr[9]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_8\, S => \rdiff_bus[9]\, Y => OPEN, FCO
         => \rdiff_bus_cry_9\);
    
    \memwaddr_r[0]\ : SLE
      port map(D => \memwaddr_r_s[0]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_862, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[0]\);
    
    fulli_0_a2_7 : CFG4
      generic map(INIT => x"8000")

      port map(A => \wdiff_bus[6]\, B => \wdiff_bus[7]\, C => 
        \wdiff_bus[8]\, D => \wdiff_bus[9]\, Y => \fulli_0_a2_7\);
    
    \wptr_gray[2]\ : SLE
      port map(D => \wptr_gray_1[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[2]_net_1\);
    
    wdiff_bus_cry_4 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[4]_net_1\, B => 
        \rptr_bin_sync2[4]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_3\, S => \wdiff_bus[4]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_4\);
    
    \memwaddr_r_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[2]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[1]_net_1\, S => \memwaddr_r_s[2]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[2]_net_1\);
    
    \wptr_gray[11]\ : SLE
      port map(D => \wptr[11]_net_1\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr_gray[11]_net_1\);
    
    \wptr_bin_sync2[9]\ : SLE
      port map(D => \wptr_bin_sync[9]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[9]_net_1\);
    
    \rptr_gray_1[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[6]_net_1\, B => \rptr[7]_net_1\, Y => 
        \rptr_gray_1[6]_net_1\);
    
    \wptr_gray_1[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[11]_net_1\, B => \wptr[10]_net_1\, Y
         => \wptr_gray_1[10]_net_1\);
    
    wdiff_bus_cry_6 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[6]_net_1\, B => 
        \rptr_bin_sync2[6]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_5\, S => \wdiff_bus[6]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_6\);
    
    \rptr_s[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[10]_net_1\, S
         => \rptr_s[11]_net_1\, Y => OPEN, FCO => OPEN);
    
    \rptr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[2]_net_1\, S
         => \rptr_s[3]\, Y => OPEN, FCO => \rptr_cry[3]_net_1\);
    
    \memraddr_r[4]\ : SLE
      port map(D => \memraddr_r_s[4]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_140_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[4]\);
    
    \memraddr_r_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[6]_net_1\, S => \memraddr_r_s[7]\, Y => 
        OPEN, FCO => \memraddr_r_cry[7]_net_1\);
    
    fulli_0_a2_8 : CFG4
      generic map(INIT => x"4000")

      port map(A => wdiff_bus_cry_0_Y_1, B => \wdiff_bus[1]\, C
         => \wdiff_bus[10]\, D => \fulli_0_a2_6\, Y => 
        \fulli_0_a2_8\);
    
    \memraddr_r_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[9]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[8]_net_1\, S => \memraddr_r_s[9]\, Y => 
        OPEN, FCO => \memraddr_r_cry[9]_net_1\);
    
    \memraddr_r[5]\ : SLE
      port map(D => \memraddr_r_s[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_140_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[5]\);
    
    \rptr_gray[6]\ : SLE
      port map(D => \rptr_gray_1[6]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[6]_net_1\);
    
    \memraddr_r[9]\ : SLE
      port map(D => \memraddr_r_s[9]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_140_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[9]\);
    
    \rptr[0]\ : SLE
      port map(D => \rptr_s[0]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_140_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[0]_net_1\);
    
    \wptr[10]\ : SLE
      port map(D => \wptr_s[10]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[10]_net_1\);
    
    \memwaddr_r_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[3]_net_1\, S => \memwaddr_r_s[4]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[4]_net_1\);
    
    \memraddr_r_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[3]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[2]_net_1\, S => \memraddr_r_s[3]\, Y => 
        OPEN, FCO => \memraddr_r_cry[3]_net_1\);
    
    wdiff_bus_cry_1 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[1]_net_1\, B => 
        \rptr_bin_sync2[1]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_0\, S => \wdiff_bus[1]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_1\);
    
    rdiff_bus_cry_2 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[2]_net_1\, B => 
        \rptr[2]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_1\, S => \rdiff_bus[2]\, Y => OPEN, FCO
         => \rdiff_bus_cry_2\);
    
    \wptr_gray[9]\ : SLE
      port map(D => \wptr_gray_1[9]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[9]_net_1\);
    
    \rptr_gray_1[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[4]_net_1\, B => \rptr[5]_net_1\, Y => 
        \rptr_gray_1[4]_net_1\);
    
    \wptr_gray_1[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[8]_net_1\, B => \wptr[9]_net_1\, Y => 
        \wptr_gray_1[8]_net_1\);
    
    Rd_corefifo_grayToBinConv : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_1
      port map(rptr_bin_sync(11) => \rptr_bin_sync[11]\, 
        rptr_bin_sync(10) => \rptr_bin_sync[10]\, 
        rptr_bin_sync(9) => \rptr_bin_sync[9]\, rptr_bin_sync(8)
         => \rptr_bin_sync[8]\, rptr_bin_sync(7) => 
        \rptr_bin_sync[7]\, rptr_bin_sync(6) => 
        \rptr_bin_sync[6]\, rptr_bin_sync(5) => 
        \rptr_bin_sync[5]\, rptr_bin_sync(4) => 
        \rptr_bin_sync[4]\, rptr_bin_sync(3) => 
        \rptr_bin_sync[3]\, rptr_bin_sync(2) => 
        \rptr_bin_sync[2]\, rptr_bin_sync(1) => 
        \rptr_bin_sync[1]\, rptr_bin_sync(0) => 
        \rptr_bin_sync[0]\, rptr_gray_sync(10) => 
        \rptr_gray_sync[10]\, rptr_gray_sync(9) => 
        \rptr_gray_sync[9]\, rptr_gray_sync(8) => 
        \rptr_gray_sync[8]\, rptr_gray_sync(7) => 
        \rptr_gray_sync[7]\, rptr_gray_sync(6) => 
        \rptr_gray_sync[6]\, rptr_gray_sync(5) => 
        \rptr_gray_sync[5]\, rptr_gray_sync(4) => 
        \rptr_gray_sync[4]\, rptr_gray_sync(3) => 
        \rptr_gray_sync[3]\, rptr_gray_sync(2) => 
        \rptr_gray_sync[2]\, rptr_gray_sync(1) => 
        \rptr_gray_sync[1]\, rptr_gray_sync(0) => 
        \rptr_gray_sync[0]\);
    
    \rptr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => rptr_s_380_FCO, S => 
        \rptr_s[1]\, Y => OPEN, FCO => \rptr_cry[1]_net_1\);
    
    rdiff_bus_cry_3 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[3]_net_1\, B => 
        \rptr[3]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_2\, S => \rdiff_bus[3]\, Y => OPEN, FCO
         => \rdiff_bus_cry_3\);
    
    rdiff_bus_cry_10 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[10]_net_1\, B => 
        \rptr[10]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_9\, S => \rdiff_bus[10]\, Y => OPEN, FCO
         => \rdiff_bus_cry_10\);
    
    \memraddr_r_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[5]_net_1\, S => \memraddr_r_s[6]\, Y => 
        OPEN, FCO => \memraddr_r_cry[6]_net_1\);
    
    \memraddr_r[6]\ : SLE
      port map(D => \memraddr_r_s[6]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_140_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[6]\);
    
    \rptr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[6]_net_1\, S
         => \rptr_s[7]\, Y => OPEN, FCO => \rptr_cry[7]_net_1\);
    
    wptr_s_382 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => wptr_s_382_FCO);
    
    rdiff_bus_cry_0 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => rdiff_bus, B => \rptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => rdiff_bus_cry_0_Y_1, FCO => \rdiff_bus_cry_0\);
    
    \memraddr_r[2]\ : SLE
      port map(D => \memraddr_r_s[2]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_140_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[2]\);
    
    \wptr[8]\ : SLE
      port map(D => \wptr_s[8]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[8]_net_1\);
    
    wdiff_bus_cry_3 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[3]_net_1\, B => 
        \rptr_bin_sync2[3]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_2\, S => \wdiff_bus[3]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_3\);
    
    \rptr_gray[7]\ : SLE
      port map(D => \rptr_gray_1[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[7]_net_1\);
    
    \wptr_gray[0]\ : SLE
      port map(D => \wptr_gray_1[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[0]_net_1\);
    
    \rptr_gray_1[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[0]_net_1\, B => \rptr[1]_net_1\, Y => 
        \rptr_gray_1[0]_net_1\);
    
    \rptr_gray_1[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[8]_net_1\, B => \rptr[9]_net_1\, Y => 
        \rptr_gray_1[8]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_0 is

    port( RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          ReadFIFO_Write_Ptr        : in    std_logic_vector(1 downto 0);
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          RX_FIFO_DOUT_1_0          : out   std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          N_1466                    : in    std_logic;
          N_660                     : out   std_logic;
          N_662                     : out   std_logic;
          N_663                     : out   std_logic;
          N_717                     : out   std_logic;
          N_661                     : out   std_logic;
          N_659                     : out   std_logic;
          N_658                     : out   std_logic;
          N_657                     : out   std_logic;
          N_1003                    : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          irx_fifo_rst_i            : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_0;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_0
    port( RDATA_int                 : out   std_logic_vector(8 downto 0);
          fifo_MEMRADDR             : in    std_logic_vector(10 downto 0) := (others => 'U');
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          fifo_MEMWADDR             : in    std_logic_vector(10 downto 0) := (others => 'U');
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          N_140_i                   : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          fifo_MEMWE                : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_0
    port( ReadFIFO_Write_Ptr        : in    std_logic_vector(1 downto 0) := (others => 'U');
          fifo_MEMWADDR             : out   std_logic_vector(10 downto 0);
          fifo_MEMRADDR             : out   std_logic_vector(10 downto 0);
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          N_152_i_i                 : out   std_logic;
          N_89_i                    : out   std_logic;
          REN_d1                    : in    std_logic := 'U';
          N_1003                    : in    std_logic := 'U';
          N_1466                    : in    std_logic := 'U';
          N_140_i                   : out   std_logic;
          fifo_MEMWE                : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          irx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \RDATA_r[4]_net_1\, VCC_net_1, \RDATA_int[4]\, N_89_i, 
        GND_net_1, \RDATA_r[5]_net_1\, \RDATA_int[5]\, 
        \RDATA_r[6]_net_1\, \RDATA_int[6]\, \RDATA_r[7]_net_1\, 
        \RDATA_int[7]\, \RDATA_r[8]_net_1\, \RDATA_int[8]\, 
        \re_set\, \REN_d1\, N_152_i_i, \RDATA_r[0]_net_1\, 
        \RDATA_int[0]\, \RDATA_r[1]_net_1\, \RDATA_int[1]\, 
        \RDATA_r[2]_net_1\, \RDATA_int[2]\, \RDATA_r[3]_net_1\, 
        \RDATA_int[3]\, N_140_i, \RE_d1\, \re_pulse_d1\, 
        \re_pulse\, \iRX_FIFO_Empty_0\, \fifo_MEMWADDR[0]\, 
        \fifo_MEMWADDR[1]\, \fifo_MEMWADDR[2]\, 
        \fifo_MEMWADDR[3]\, \fifo_MEMWADDR[4]\, 
        \fifo_MEMWADDR[5]\, \fifo_MEMWADDR[6]\, 
        \fifo_MEMWADDR[7]\, \fifo_MEMWADDR[8]\, 
        \fifo_MEMWADDR[9]\, \fifo_MEMWADDR[10]\, 
        \fifo_MEMRADDR[0]\, \fifo_MEMRADDR[1]\, 
        \fifo_MEMRADDR[2]\, \fifo_MEMRADDR[3]\, 
        \fifo_MEMRADDR[4]\, \fifo_MEMRADDR[5]\, 
        \fifo_MEMRADDR[6]\, \fifo_MEMRADDR[7]\, 
        \fifo_MEMRADDR[8]\, \fifo_MEMRADDR[9]\, 
        \fifo_MEMRADDR[10]\, fifo_MEMWE : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_0
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_0(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_0
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_0(DEF_ARCH);
begin 

    iRX_FIFO_Empty_0 <= \iRX_FIFO_Empty_0\;

    re_pulse : CFG4
      generic map(INIT => x"FAF2")

      port map(A => \REN_d1\, B => N_1003, C => \re_set\, D => 
        \iRX_FIFO_Empty_0\, Y => \re_pulse\);
    
    \RDATA_r[3]\ : SLE
      port map(D => \RDATA_int[3]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[3]_net_1\);
    
    \Q_i_m2[2]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[2]_net_1\, C => 
        \RDATA_int[2]\, D => \RE_d1\, Y => N_658);
    
    re_pulse_d1 : SLE
      port map(D => \re_pulse\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \re_pulse_d1\);
    
    \RDATA_r[5]\ : SLE
      port map(D => \RDATA_int[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[5]_net_1\);
    
    \Q_i_m2[0]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[0]_net_1\, C => 
        \RDATA_int[0]\, D => \RE_d1\, Y => N_657);
    
    \Q_i_m2[3]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[3]_net_1\, C => 
        \RDATA_int[3]\, D => \RE_d1\, Y => N_659);
    
    \RDATA_r[8]\ : SLE
      port map(D => \RDATA_int[8]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[8]_net_1\);
    
    \Q_i_m2[7]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[7]_net_1\, C => 
        \RDATA_int[7]\, D => \RE_d1\, Y => N_663);
    
    \Q_i_m2[6]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[6]_net_1\, C => 
        \RDATA_int[6]\, D => \RE_d1\, Y => N_662);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \RW1.UI_ram_wrapper_1\ : FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_0
      port map(RDATA_int(8) => \RDATA_int[8]\, RDATA_int(7) => 
        \RDATA_int[7]\, RDATA_int(6) => \RDATA_int[6]\, 
        RDATA_int(5) => \RDATA_int[5]\, RDATA_int(4) => 
        \RDATA_int[4]\, RDATA_int(3) => \RDATA_int[3]\, 
        RDATA_int(2) => \RDATA_int[2]\, RDATA_int(1) => 
        \RDATA_int[1]\, RDATA_int(0) => \RDATA_int[0]\, 
        fifo_MEMRADDR(10) => \fifo_MEMRADDR[10]\, 
        fifo_MEMRADDR(9) => \fifo_MEMRADDR[9]\, fifo_MEMRADDR(8)
         => \fifo_MEMRADDR[8]\, fifo_MEMRADDR(7) => 
        \fifo_MEMRADDR[7]\, fifo_MEMRADDR(6) => 
        \fifo_MEMRADDR[6]\, fifo_MEMRADDR(5) => 
        \fifo_MEMRADDR[5]\, fifo_MEMRADDR(4) => 
        \fifo_MEMRADDR[4]\, fifo_MEMRADDR(3) => 
        \fifo_MEMRADDR[3]\, fifo_MEMRADDR(2) => 
        \fifo_MEMRADDR[2]\, fifo_MEMRADDR(1) => 
        \fifo_MEMRADDR[1]\, fifo_MEMRADDR(0) => 
        \fifo_MEMRADDR[0]\, RX_FIFO_DIN_pipe(8) => 
        RX_FIFO_DIN_pipe(8), RX_FIFO_DIN_pipe(7) => 
        RX_FIFO_DIN_pipe(7), RX_FIFO_DIN_pipe(6) => 
        RX_FIFO_DIN_pipe(6), RX_FIFO_DIN_pipe(5) => 
        RX_FIFO_DIN_pipe(5), RX_FIFO_DIN_pipe(4) => 
        RX_FIFO_DIN_pipe(4), RX_FIFO_DIN_pipe(3) => 
        RX_FIFO_DIN_pipe(3), RX_FIFO_DIN_pipe(2) => 
        RX_FIFO_DIN_pipe(2), RX_FIFO_DIN_pipe(1) => 
        RX_FIFO_DIN_pipe(1), RX_FIFO_DIN_pipe(0) => 
        RX_FIFO_DIN_pipe(0), fifo_MEMWADDR(10) => 
        \fifo_MEMWADDR[10]\, fifo_MEMWADDR(9) => 
        \fifo_MEMWADDR[9]\, fifo_MEMWADDR(8) => 
        \fifo_MEMWADDR[8]\, fifo_MEMWADDR(7) => 
        \fifo_MEMWADDR[7]\, fifo_MEMWADDR(6) => 
        \fifo_MEMWADDR[6]\, fifo_MEMWADDR(5) => 
        \fifo_MEMWADDR[5]\, fifo_MEMWADDR(4) => 
        \fifo_MEMWADDR[4]\, fifo_MEMWADDR(3) => 
        \fifo_MEMWADDR[3]\, fifo_MEMWADDR(2) => 
        \fifo_MEMWADDR[2]\, fifo_MEMWADDR(1) => 
        \fifo_MEMWADDR[1]\, fifo_MEMWADDR(0) => 
        \fifo_MEMWADDR[0]\, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, N_140_i => N_140_i, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, fifo_MEMWE
         => fifo_MEMWE);
    
    \RDATA_r[0]\ : SLE
      port map(D => \RDATA_int[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[0]_net_1\);
    
    \Q_i_m2[5]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[5]_net_1\, C => 
        \RDATA_int[5]\, D => \RE_d1\, Y => N_661);
    
    \RDATA_r[2]\ : SLE
      port map(D => \RDATA_int[2]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[2]_net_1\);
    
    \RDATA_r[6]\ : SLE
      port map(D => \RDATA_int[6]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[6]_net_1\);
    
    \L31.U_corefifo_async\ : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_0
      port map(ReadFIFO_Write_Ptr(1) => ReadFIFO_Write_Ptr(1), 
        ReadFIFO_Write_Ptr(0) => ReadFIFO_Write_Ptr(0), 
        fifo_MEMWADDR(10) => \fifo_MEMWADDR[10]\, 
        fifo_MEMWADDR(9) => \fifo_MEMWADDR[9]\, fifo_MEMWADDR(8)
         => \fifo_MEMWADDR[8]\, fifo_MEMWADDR(7) => 
        \fifo_MEMWADDR[7]\, fifo_MEMWADDR(6) => 
        \fifo_MEMWADDR[6]\, fifo_MEMWADDR(5) => 
        \fifo_MEMWADDR[5]\, fifo_MEMWADDR(4) => 
        \fifo_MEMWADDR[4]\, fifo_MEMWADDR(3) => 
        \fifo_MEMWADDR[3]\, fifo_MEMWADDR(2) => 
        \fifo_MEMWADDR[2]\, fifo_MEMWADDR(1) => 
        \fifo_MEMWADDR[1]\, fifo_MEMWADDR(0) => 
        \fifo_MEMWADDR[0]\, fifo_MEMRADDR(10) => 
        \fifo_MEMRADDR[10]\, fifo_MEMRADDR(9) => 
        \fifo_MEMRADDR[9]\, fifo_MEMRADDR(8) => 
        \fifo_MEMRADDR[8]\, fifo_MEMRADDR(7) => 
        \fifo_MEMRADDR[7]\, fifo_MEMRADDR(6) => 
        \fifo_MEMRADDR[6]\, fifo_MEMRADDR(5) => 
        \fifo_MEMRADDR[5]\, fifo_MEMRADDR(4) => 
        \fifo_MEMRADDR[4]\, fifo_MEMRADDR(3) => 
        \fifo_MEMRADDR[3]\, fifo_MEMRADDR(2) => 
        \fifo_MEMRADDR[2]\, fifo_MEMRADDR(1) => 
        \fifo_MEMRADDR[1]\, fifo_MEMRADDR(0) => 
        \fifo_MEMRADDR[0]\, iRX_FIFO_Empty_0 => 
        \iRX_FIFO_Empty_0\, iRX_FIFO_UNDERRUN_0 => 
        iRX_FIFO_UNDERRUN_0, iRX_FIFO_Full_0 => iRX_FIFO_Full_0, 
        iRX_FIFO_OVERFLOW_0 => iRX_FIFO_OVERFLOW_0, N_152_i_i => 
        N_152_i_i, N_89_i => N_89_i, REN_d1 => \REN_d1\, N_1003
         => N_1003, N_1466 => N_1466, N_140_i => N_140_i, 
        fifo_MEMWE => fifo_MEMWE, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, irx_fifo_rst_i => irx_fifo_rst_i);
    
    re_set : SLE
      port map(D => \REN_d1\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => N_152_i_i, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \re_set\);
    
    \Q_i_m2[8]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[8]_net_1\, C => 
        \RDATA_int[8]\, D => \RE_d1\, Y => N_717);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    RE_d1 : SLE
      port map(D => N_1003, CLK => m2s010_som_sb_0_CCC_71MHz, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \RE_d1\);
    
    \RDATA_r[7]\ : SLE
      port map(D => \RDATA_int[7]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[7]_net_1\);
    
    \RDATA_r[4]\ : SLE
      port map(D => \RDATA_int[4]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[4]_net_1\);
    
    \Q[1]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[1]_net_1\, C => 
        \RDATA_int[1]\, D => \RE_d1\, Y => RX_FIFO_DOUT_1_0);
    
    REN_d1 : SLE
      port map(D => N_140_i, CLK => m2s010_som_sb_0_CCC_71MHz, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \REN_d1\);
    
    \Q_i_m2[4]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[4]_net_1\, C => 
        \RDATA_int[4]\, D => \RE_d1\, Y => N_660);
    
    \RDATA_r[1]\ : SLE
      port map(D => \RDATA_int[1]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[1]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_0 is

    port( ReadFIFO_Write_Ptr        : in    std_logic_vector(1 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          RX_FIFO_DOUT_1_0          : out   std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          irx_fifo_rst_i            : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          N_1003                    : in    std_logic;
          N_657                     : out   std_logic;
          N_658                     : out   std_logic;
          N_659                     : out   std_logic;
          N_661                     : out   std_logic;
          N_717                     : out   std_logic;
          N_663                     : out   std_logic;
          N_662                     : out   std_logic;
          N_660                     : out   std_logic;
          N_1466                    : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic
        );

end FIFO_8Kx9_0;

architecture DEF_ARCH of FIFO_8Kx9_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_0
    port( RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          ReadFIFO_Write_Ptr        : in    std_logic_vector(1 downto 0) := (others => 'U');
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          RX_FIFO_DOUT_1_0          : out   std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          N_1466                    : in    std_logic := 'U';
          N_660                     : out   std_logic;
          N_662                     : out   std_logic;
          N_663                     : out   std_logic;
          N_717                     : out   std_logic;
          N_661                     : out   std_logic;
          N_659                     : out   std_logic;
          N_658                     : out   std_logic;
          N_657                     : out   std_logic;
          N_1003                    : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          irx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_0
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_0(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    FIFO_8Kx9_0 : FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_0
      port map(RX_FIFO_DIN_pipe(8) => RX_FIFO_DIN_pipe(8), 
        RX_FIFO_DIN_pipe(7) => RX_FIFO_DIN_pipe(7), 
        RX_FIFO_DIN_pipe(6) => RX_FIFO_DIN_pipe(6), 
        RX_FIFO_DIN_pipe(5) => RX_FIFO_DIN_pipe(5), 
        RX_FIFO_DIN_pipe(4) => RX_FIFO_DIN_pipe(4), 
        RX_FIFO_DIN_pipe(3) => RX_FIFO_DIN_pipe(3), 
        RX_FIFO_DIN_pipe(2) => RX_FIFO_DIN_pipe(2), 
        RX_FIFO_DIN_pipe(1) => RX_FIFO_DIN_pipe(1), 
        RX_FIFO_DIN_pipe(0) => RX_FIFO_DIN_pipe(0), 
        ReadFIFO_Write_Ptr(1) => ReadFIFO_Write_Ptr(1), 
        ReadFIFO_Write_Ptr(0) => ReadFIFO_Write_Ptr(0), 
        iRX_FIFO_OVERFLOW_0 => iRX_FIFO_OVERFLOW_0, 
        iRX_FIFO_Full_0 => iRX_FIFO_Full_0, iRX_FIFO_UNDERRUN_0
         => iRX_FIFO_UNDERRUN_0, iRX_FIFO_Empty_0 => 
        iRX_FIFO_Empty_0, RX_FIFO_DOUT_1_0 => RX_FIFO_DOUT_1_0, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, N_1466 => 
        N_1466, N_660 => N_660, N_662 => N_662, N_663 => N_663, 
        N_717 => N_717, N_661 => N_661, N_659 => N_659, N_658 => 
        N_658, N_657 => N_657, N_1003 => N_1003, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz, 
        irx_fifo_rst_i => irx_fifo_rst_i);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_1 is

    port( fifo_MEMWADDR             : in    std_logic_vector(10 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          fifo_MEMRADDR             : in    std_logic_vector(10 downto 0);
          RDATA_int                 : out   std_logic_vector(8 downto 0);
          fifo_MEMWE                : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          N_1005_i                  : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_1;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_1 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component RAM1K18
    generic (MEMORYFILE:string := "");

    port( A_DOUT        : out   std_logic_vector(17 downto 0);
          B_DOUT        : out   std_logic_vector(17 downto 0);
          BUSY          : out   std_logic;
          A_CLK         : in    std_logic := 'U';
          A_DOUT_CLK    : in    std_logic := 'U';
          A_ARST_N      : in    std_logic := 'U';
          A_DOUT_EN     : in    std_logic := 'U';
          A_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_DOUT_ARST_N : in    std_logic := 'U';
          A_DOUT_SRST_N : in    std_logic := 'U';
          A_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          A_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          A_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          B_CLK         : in    std_logic := 'U';
          B_DOUT_CLK    : in    std_logic := 'U';
          B_ARST_N      : in    std_logic := 'U';
          B_DOUT_EN     : in    std_logic := 'U';
          B_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_DOUT_ARST_N : in    std_logic := 'U';
          B_DOUT_SRST_N : in    std_logic := 'U';
          B_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          B_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          B_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          A_EN          : in    std_logic := 'U';
          A_DOUT_LAT    : in    std_logic := 'U';
          A_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_WMODE       : in    std_logic := 'U';
          B_EN          : in    std_logic := 'U';
          B_DOUT_LAT    : in    std_logic := 'U';
          B_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_WMODE       : in    std_logic := 'U';
          SII_LOCK      : in    std_logic := 'U'
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;
    signal nc24, nc1, nc8, nc13, nc16, nc19, nc25, nc20, nc27, 
        nc9, nc22, nc14, nc5, nc21, nc15, nc3, nc10, nc7, nc17, 
        nc4, nc12, nc2, nc23, nc18, nc26, nc6, nc11 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C0 : RAM1K18
      port map(A_DOUT(17) => nc24, A_DOUT(16) => nc1, A_DOUT(15)
         => nc8, A_DOUT(14) => nc13, A_DOUT(13) => nc16, 
        A_DOUT(12) => nc19, A_DOUT(11) => nc25, A_DOUT(10) => 
        nc20, A_DOUT(9) => nc27, A_DOUT(8) => RDATA_int(8), 
        A_DOUT(7) => RDATA_int(7), A_DOUT(6) => RDATA_int(6), 
        A_DOUT(5) => RDATA_int(5), A_DOUT(4) => RDATA_int(4), 
        A_DOUT(3) => RDATA_int(3), A_DOUT(2) => RDATA_int(2), 
        A_DOUT(1) => RDATA_int(1), A_DOUT(0) => RDATA_int(0), 
        B_DOUT(17) => nc9, B_DOUT(16) => nc22, B_DOUT(15) => nc14, 
        B_DOUT(14) => nc5, B_DOUT(13) => nc21, B_DOUT(12) => nc15, 
        B_DOUT(11) => nc3, B_DOUT(10) => nc10, B_DOUT(9) => nc7, 
        B_DOUT(8) => nc17, B_DOUT(7) => nc4, B_DOUT(6) => nc12, 
        B_DOUT(5) => nc2, B_DOUT(4) => nc23, B_DOUT(3) => nc18, 
        B_DOUT(2) => nc26, B_DOUT(1) => nc6, B_DOUT(0) => nc11, 
        BUSY => OPEN, A_CLK => m2s010_som_sb_0_CCC_71MHz, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => VCC_net_1, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_1005_i, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => GND_net_1, A_DIN(15) => GND_net_1, 
        A_DIN(14) => GND_net_1, A_DIN(13) => GND_net_1, A_DIN(12)
         => GND_net_1, A_DIN(11) => GND_net_1, A_DIN(10) => 
        GND_net_1, A_DIN(9) => GND_net_1, A_DIN(8) => GND_net_1, 
        A_DIN(7) => GND_net_1, A_DIN(6) => GND_net_1, A_DIN(5)
         => GND_net_1, A_DIN(4) => GND_net_1, A_DIN(3) => 
        GND_net_1, A_DIN(2) => GND_net_1, A_DIN(1) => GND_net_1, 
        A_DIN(0) => GND_net_1, A_ADDR(13) => fifo_MEMRADDR(10), 
        A_ADDR(12) => fifo_MEMRADDR(9), A_ADDR(11) => 
        fifo_MEMRADDR(8), A_ADDR(10) => fifo_MEMRADDR(7), 
        A_ADDR(9) => fifo_MEMRADDR(6), A_ADDR(8) => 
        fifo_MEMRADDR(5), A_ADDR(7) => fifo_MEMRADDR(4), 
        A_ADDR(6) => fifo_MEMRADDR(3), A_ADDR(5) => 
        fifo_MEMRADDR(2), A_ADDR(4) => fifo_MEMRADDR(1), 
        A_ADDR(3) => fifo_MEMRADDR(0), A_ADDR(2) => GND_net_1, 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => RX_FIFO_DIN_pipe(8), B_DIN(7) => RX_FIFO_DIN_pipe(7), 
        B_DIN(6) => RX_FIFO_DIN_pipe(6), B_DIN(5) => 
        RX_FIFO_DIN_pipe(5), B_DIN(4) => RX_FIFO_DIN_pipe(4), 
        B_DIN(3) => RX_FIFO_DIN_pipe(3), B_DIN(2) => 
        RX_FIFO_DIN_pipe(2), B_DIN(1) => RX_FIFO_DIN_pipe(1), 
        B_DIN(0) => RX_FIFO_DIN_pipe(0), B_ADDR(13) => 
        fifo_MEMWADDR(10), B_ADDR(12) => fifo_MEMWADDR(9), 
        B_ADDR(11) => fifo_MEMWADDR(8), B_ADDR(10) => 
        fifo_MEMWADDR(7), B_ADDR(9) => fifo_MEMWADDR(6), 
        B_ADDR(8) => fifo_MEMWADDR(5), B_ADDR(7) => 
        fifo_MEMWADDR(4), B_ADDR(6) => fifo_MEMWADDR(3), 
        B_ADDR(5) => fifo_MEMWADDR(2), B_ADDR(4) => 
        fifo_MEMWADDR(1), B_ADDR(3) => fifo_MEMWADDR(0), 
        B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, B_ADDR(0)
         => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0) => 
        VCC_net_1, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_1 is

    port( RDATA_int                 : out   std_logic_vector(8 downto 0);
          fifo_MEMRADDR             : in    std_logic_vector(10 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          fifo_MEMWADDR             : in    std_logic_vector(10 downto 0);
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          N_1005_i                  : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          fifo_MEMWE                : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_1;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_1 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_1
    port( fifo_MEMWADDR             : in    std_logic_vector(10 downto 0) := (others => 'U');
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          fifo_MEMRADDR             : in    std_logic_vector(10 downto 0) := (others => 'U');
          RDATA_int                 : out   std_logic_vector(8 downto 0);
          fifo_MEMWE                : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          N_1005_i                  : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_1
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_1(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    L1_asyncnonpipe : FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_1
      port map(fifo_MEMWADDR(10) => fifo_MEMWADDR(10), 
        fifo_MEMWADDR(9) => fifo_MEMWADDR(9), fifo_MEMWADDR(8)
         => fifo_MEMWADDR(8), fifo_MEMWADDR(7) => 
        fifo_MEMWADDR(7), fifo_MEMWADDR(6) => fifo_MEMWADDR(6), 
        fifo_MEMWADDR(5) => fifo_MEMWADDR(5), fifo_MEMWADDR(4)
         => fifo_MEMWADDR(4), fifo_MEMWADDR(3) => 
        fifo_MEMWADDR(3), fifo_MEMWADDR(2) => fifo_MEMWADDR(2), 
        fifo_MEMWADDR(1) => fifo_MEMWADDR(1), fifo_MEMWADDR(0)
         => fifo_MEMWADDR(0), RX_FIFO_DIN_pipe(8) => 
        RX_FIFO_DIN_pipe(8), RX_FIFO_DIN_pipe(7) => 
        RX_FIFO_DIN_pipe(7), RX_FIFO_DIN_pipe(6) => 
        RX_FIFO_DIN_pipe(6), RX_FIFO_DIN_pipe(5) => 
        RX_FIFO_DIN_pipe(5), RX_FIFO_DIN_pipe(4) => 
        RX_FIFO_DIN_pipe(4), RX_FIFO_DIN_pipe(3) => 
        RX_FIFO_DIN_pipe(3), RX_FIFO_DIN_pipe(2) => 
        RX_FIFO_DIN_pipe(2), RX_FIFO_DIN_pipe(1) => 
        RX_FIFO_DIN_pipe(1), RX_FIFO_DIN_pipe(0) => 
        RX_FIFO_DIN_pipe(0), fifo_MEMRADDR(10) => 
        fifo_MEMRADDR(10), fifo_MEMRADDR(9) => fifo_MEMRADDR(9), 
        fifo_MEMRADDR(8) => fifo_MEMRADDR(8), fifo_MEMRADDR(7)
         => fifo_MEMRADDR(7), fifo_MEMRADDR(6) => 
        fifo_MEMRADDR(6), fifo_MEMRADDR(5) => fifo_MEMRADDR(5), 
        fifo_MEMRADDR(4) => fifo_MEMRADDR(4), fifo_MEMRADDR(3)
         => fifo_MEMRADDR(3), fifo_MEMRADDR(2) => 
        fifo_MEMRADDR(2), fifo_MEMRADDR(1) => fifo_MEMRADDR(1), 
        fifo_MEMRADDR(0) => fifo_MEMRADDR(0), RDATA_int(8) => 
        RDATA_int(8), RDATA_int(7) => RDATA_int(7), RDATA_int(6)
         => RDATA_int(6), RDATA_int(5) => RDATA_int(5), 
        RDATA_int(4) => RDATA_int(4), RDATA_int(3) => 
        RDATA_int(3), RDATA_int(2) => RDATA_int(2), RDATA_int(1)
         => RDATA_int(1), RDATA_int(0) => RDATA_int(0), 
        fifo_MEMWE => fifo_MEMWE, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, N_1005_i => N_1005_i, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_4 is

    port( wptr_bin_sync  : inout std_logic_vector(11 downto 0) := (others => 'Z');
          wptr_gray_sync : in    std_logic_vector(10 downto 0)
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_4;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_4 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    \bin_out_xhdl1_0_a2[1]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(3), B => wptr_gray_sync(1), C
         => wptr_bin_sync(4), D => wptr_gray_sync(2), Y => 
        wptr_bin_sync(1));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \bin_out_xhdl1_0_a2[5]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(7), B => wptr_gray_sync(6), C
         => wptr_gray_sync(5), D => wptr_bin_sync(8), Y => 
        wptr_bin_sync(5));
    
    \bin_out_xhdl1_0_a2[2]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(4), B => wptr_gray_sync(3), C
         => wptr_gray_sync(2), D => wptr_bin_sync(5), Y => 
        wptr_bin_sync(2));
    
    \bin_out_xhdl1_0_a2[0]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(2), B => wptr_bin_sync(3), C
         => wptr_gray_sync(0), D => wptr_gray_sync(1), Y => 
        wptr_bin_sync(0));
    
    \bin_out_xhdl1_i_o2[9]\ : CFG3
      generic map(INIT => x"96")

      port map(A => wptr_gray_sync(10), B => wptr_gray_sync(9), C
         => wptr_bin_sync(11), Y => wptr_bin_sync(9));
    
    \bin_out_xhdl1_i_o2[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => wptr_bin_sync(11), B => wptr_gray_sync(10), Y
         => wptr_bin_sync(10));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \bin_out_xhdl1_0_a2[6]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(8), B => wptr_gray_sync(7), C
         => wptr_gray_sync(6), D => wptr_bin_sync(9), Y => 
        wptr_bin_sync(6));
    
    \bin_out_xhdl1_0_a2[4]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(6), B => wptr_gray_sync(5), C
         => wptr_gray_sync(4), D => wptr_bin_sync(7), Y => 
        wptr_bin_sync(4));
    
    \bin_out_xhdl1_0_a2[8]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(10), B => wptr_gray_sync(9), C
         => wptr_gray_sync(8), D => wptr_bin_sync(11), Y => 
        wptr_bin_sync(8));
    
    \bin_out_xhdl1_0_a2[7]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(9), B => wptr_gray_sync(8), C
         => wptr_gray_sync(7), D => wptr_bin_sync(10), Y => 
        wptr_bin_sync(7));
    
    \bin_out_xhdl1_0_a2[3]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(5), B => wptr_gray_sync(4), C
         => wptr_gray_sync(3), D => wptr_bin_sync(6), Y => 
        wptr_bin_sync(3));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_2 is

    port( wptr_gray                 : in    std_logic_vector(11 downto 0);
          wptr_gray_sync            : out   std_logic_vector(10 downto 0);
          wptr_bin_sync_0           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          irx_fifo_rst_i            : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_2;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_2 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \sync_int[10]_net_1\, VCC_net_1, GND_net_1, 
        \sync_int[11]_net_1\, \sync_int[0]_net_1\, 
        \sync_int[1]_net_1\, \sync_int[2]_net_1\, 
        \sync_int[3]_net_1\, \sync_int[4]_net_1\, 
        \sync_int[5]_net_1\, \sync_int[6]_net_1\, 
        \sync_int[7]_net_1\, \sync_int[8]_net_1\, 
        \sync_int[9]_net_1\ : std_logic;

begin 


    \sync_int[9]\ : SLE
      port map(D => wptr_gray(9), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[9]_net_1\);
    
    \sync_int[4]\ : SLE
      port map(D => wptr_gray(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[4]_net_1\);
    
    \sync_out_xhdl1[10]\ : SLE
      port map(D => \sync_int[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(10));
    
    \sync_int[1]\ : SLE
      port map(D => wptr_gray(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[1]_net_1\);
    
    \sync_int[11]\ : SLE
      port map(D => wptr_gray(11), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[11]_net_1\);
    
    \sync_out_xhdl1[6]\ : SLE
      port map(D => \sync_int[6]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(6));
    
    \sync_out_xhdl1[3]\ : SLE
      port map(D => \sync_int[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(3));
    
    \sync_int[6]\ : SLE
      port map(D => wptr_gray(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[6]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \sync_out_xhdl1[11]\ : SLE
      port map(D => \sync_int[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_bin_sync_0);
    
    \sync_int[3]\ : SLE
      port map(D => wptr_gray(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[3]_net_1\);
    
    \sync_out_xhdl1[4]\ : SLE
      port map(D => \sync_int[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(4));
    
    \sync_int[0]\ : SLE
      port map(D => wptr_gray(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[0]_net_1\);
    
    \sync_out_xhdl1[1]\ : SLE
      port map(D => \sync_int[1]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(1));
    
    \sync_int[5]\ : SLE
      port map(D => wptr_gray(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[5]_net_1\);
    
    \sync_int[2]\ : SLE
      port map(D => wptr_gray(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[2]_net_1\);
    
    \sync_out_xhdl1[9]\ : SLE
      port map(D => \sync_int[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(9));
    
    \sync_out_xhdl1[2]\ : SLE
      port map(D => \sync_int[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(2));
    
    \sync_int[8]\ : SLE
      port map(D => wptr_gray(8), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[8]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sync_out_xhdl1[7]\ : SLE
      port map(D => \sync_int[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(7));
    
    \sync_out_xhdl1[5]\ : SLE
      port map(D => \sync_int[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(5));
    
    \sync_out_xhdl1[0]\ : SLE
      port map(D => \sync_int[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(0));
    
    \sync_out_xhdl1[8]\ : SLE
      port map(D => \sync_int[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(8));
    
    \sync_int[7]\ : SLE
      port map(D => wptr_gray(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[7]_net_1\);
    
    \sync_int[10]\ : SLE
      port map(D => wptr_gray(10), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_1 is

    port( rptr_gray           : in    std_logic_vector(11 downto 0);
          rptr_gray_sync      : out   std_logic_vector(10 downto 0);
          rptr_bin_sync_0     : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          irx_fifo_rst_i      : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_1;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_1 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \sync_int[4]_net_1\, GND_net_1, 
        \sync_int[5]_net_1\, \sync_int[6]_net_1\, 
        \sync_int[7]_net_1\, \sync_int[8]_net_1\, 
        \sync_int[9]_net_1\, \sync_int[10]_net_1\, 
        \sync_int[11]_net_1\, \sync_int[1]_net_1\, 
        \sync_int[2]_net_1\, \sync_int[3]_net_1\, 
        \sync_int[0]_net_1\ : std_logic;

begin 


    \sync_int[9]\ : SLE
      port map(D => rptr_gray(9), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[9]_net_1\);
    
    \sync_int[4]\ : SLE
      port map(D => rptr_gray(4), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[4]_net_1\);
    
    \sync_out_xhdl1[10]\ : SLE
      port map(D => \sync_int[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(10));
    
    \sync_int[1]\ : SLE
      port map(D => rptr_gray(1), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[1]_net_1\);
    
    \sync_int[11]\ : SLE
      port map(D => rptr_gray(11), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[11]_net_1\);
    
    \sync_out_xhdl1[6]\ : SLE
      port map(D => \sync_int[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(6));
    
    \sync_out_xhdl1[3]\ : SLE
      port map(D => \sync_int[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(3));
    
    \sync_int[6]\ : SLE
      port map(D => rptr_gray(6), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[6]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \sync_out_xhdl1[11]\ : SLE
      port map(D => \sync_int[11]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_bin_sync_0);
    
    \sync_int[3]\ : SLE
      port map(D => rptr_gray(3), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[3]_net_1\);
    
    \sync_out_xhdl1[4]\ : SLE
      port map(D => \sync_int[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(4));
    
    \sync_int[0]\ : SLE
      port map(D => rptr_gray(0), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[0]_net_1\);
    
    \sync_out_xhdl1[1]\ : SLE
      port map(D => \sync_int[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(1));
    
    \sync_int[5]\ : SLE
      port map(D => rptr_gray(5), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[5]_net_1\);
    
    \sync_int[2]\ : SLE
      port map(D => rptr_gray(2), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[2]_net_1\);
    
    \sync_out_xhdl1[9]\ : SLE
      port map(D => \sync_int[9]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(9));
    
    \sync_out_xhdl1[2]\ : SLE
      port map(D => \sync_int[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(2));
    
    \sync_int[8]\ : SLE
      port map(D => rptr_gray(8), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[8]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sync_out_xhdl1[7]\ : SLE
      port map(D => \sync_int[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(7));
    
    \sync_out_xhdl1[5]\ : SLE
      port map(D => \sync_int[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(5));
    
    \sync_out_xhdl1[0]\ : SLE
      port map(D => \sync_int[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(0));
    
    \sync_out_xhdl1[8]\ : SLE
      port map(D => \sync_int[8]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(8));
    
    \sync_int[7]\ : SLE
      port map(D => rptr_gray(7), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[7]_net_1\);
    
    \sync_int[10]\ : SLE
      port map(D => rptr_gray(10), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_3 is

    port( rptr_bin_sync  : inout std_logic_vector(11 downto 0) := (others => 'Z');
          rptr_gray_sync : in    std_logic_vector(10 downto 0)
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_3;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_3 is 

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    \bin_out_xhdl1_0_a2[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(2), B => rptr_gray_sync(1), Y
         => rptr_bin_sync(1));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \bin_out_xhdl1_0_a2[5]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(5), B => rptr_gray_sync(6), C
         => rptr_bin_sync(7), Y => rptr_bin_sync(5));
    
    \bin_out_xhdl1_0_a2[2]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(2), B => rptr_gray_sync(3), C
         => rptr_gray_sync(4), D => rptr_bin_sync(5), Y => 
        rptr_bin_sync(2));
    
    \bin_out_xhdl1_0_a2[0]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(1), B => rptr_bin_sync(2), C
         => rptr_gray_sync(0), Y => rptr_bin_sync(0));
    
    \bin_out_xhdl1_i_o2[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(10), B => rptr_gray_sync(9), Y
         => rptr_bin_sync(9));
    
    \bin_out_xhdl1_i_o2[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(11), B => rptr_gray_sync(10), Y
         => rptr_bin_sync(10));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \bin_out_xhdl1_0_a2[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(7), B => rptr_gray_sync(6), Y
         => rptr_bin_sync(6));
    
    \bin_out_xhdl1_0_a2[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(5), B => rptr_gray_sync(4), Y
         => rptr_bin_sync(4));
    
    \bin_out_xhdl1_0_a2[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(9), B => rptr_gray_sync(8), Y
         => rptr_bin_sync(8));
    
    \bin_out_xhdl1_0_a2[7]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(9), B => rptr_gray_sync(7), C
         => rptr_bin_sync(10), D => rptr_gray_sync(8), Y => 
        rptr_bin_sync(7));
    
    \bin_out_xhdl1_0_a2[3]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(4), B => rptr_bin_sync(5), C
         => rptr_gray_sync(3), Y => rptr_bin_sync(3));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_1 is

    port( ReadFIFO_Write_Ptr        : in    std_logic_vector(1 downto 0);
          fifo_MEMWADDR             : out   std_logic_vector(10 downto 0);
          fifo_MEMRADDR             : out   std_logic_vector(10 downto 0);
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          N_155_i_i                 : out   std_logic;
          N_89_i                    : out   std_logic;
          REN_d1                    : in    std_logic;
          N_134                     : in    std_logic;
          N_1466                    : in    std_logic;
          N_1005_i                  : out   std_logic;
          fifo_MEMWE                : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          irx_fifo_rst_i            : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_1;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_1 is 

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_4
    port( wptr_bin_sync  : inout   std_logic_vector(11 downto 0);
          wptr_gray_sync : in    std_logic_vector(10 downto 0) := (others => 'U')
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_2
    port( wptr_gray                 : in    std_logic_vector(11 downto 0) := (others => 'U');
          wptr_gray_sync            : out   std_logic_vector(10 downto 0);
          wptr_bin_sync_0           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          irx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_1
    port( rptr_gray           : in    std_logic_vector(11 downto 0) := (others => 'U');
          rptr_gray_sync      : out   std_logic_vector(10 downto 0);
          rptr_bin_sync_0     : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          irx_fifo_rst_i      : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_3
    port( rptr_bin_sync  : inout   std_logic_vector(11 downto 0);
          rptr_gray_sync : in    std_logic_vector(10 downto 0) := (others => 'U')
        );
  end component;

    signal \rptr[0]_net_1\, \rptr_s[0]\, \fifo_MEMRADDR[0]\, 
        \memraddr_r_s[0]\, \wptr[0]_net_1\, \wptr_s[0]\, 
        \wptr_gray[10]_net_1\, VCC_net_1, \wptr_gray_1[10]_net_1\, 
        GND_net_1, \wptr_gray[11]_net_1\, \wptr[11]_net_1\, 
        \rptr_gray[0]_net_1\, \rptr_gray_1[0]_net_1\, 
        \rptr_gray[1]_net_1\, \rptr_gray_1[1]_net_1\, 
        \rptr_gray[2]_net_1\, \rptr_gray_1[2]_net_1\, 
        \rptr_gray[3]_net_1\, \rptr_gray_1[3]_net_1\, 
        \rptr_gray[4]_net_1\, \rptr_gray_1[4]_net_1\, 
        \rptr_gray[5]_net_1\, \rptr_gray_1[5]_net_1\, 
        \rptr_gray[6]_net_1\, \rptr_gray_1[6]_net_1\, 
        \rptr_gray[7]_net_1\, \rptr_gray_1[7]_net_1\, 
        \rptr_gray[8]_net_1\, \rptr_gray_1[8]_net_1\, 
        \rptr_gray[9]_net_1\, \rptr_gray_1[9]_net_1\, 
        \rptr_gray[10]_net_1\, \rptr_gray_1[10]_net_1\, 
        \rptr_gray[11]_net_1\, \rptr[11]_net_1\, 
        \wptr_bin_sync2[7]_net_1\, \wptr_bin_sync[7]\, 
        \wptr_bin_sync2[8]_net_1\, \wptr_bin_sync[8]\, 
        \wptr_bin_sync2[9]_net_1\, \wptr_bin_sync[9]\, 
        \wptr_bin_sync2[10]_net_1\, \wptr_bin_sync[10]\, 
        \wptr_bin_sync2[11]_net_1\, \wptr_bin_sync[11]\, 
        \wptr_gray[0]_net_1\, \wptr_gray_1[0]_net_1\, 
        \wptr_gray[1]_net_1\, \wptr_gray_1[1]_net_1\, 
        \wptr_gray[2]_net_1\, \wptr_gray_1[2]_net_1\, 
        \wptr_gray[3]_net_1\, \wptr_gray_1[3]_net_1\, 
        \wptr_gray[4]_net_1\, \wptr_gray_1[4]_net_1\, 
        \wptr_gray[5]_net_1\, \wptr_gray_1[5]_net_1\, 
        \wptr_gray[6]_net_1\, \wptr_gray_1[6]_net_1\, 
        \wptr_gray[7]_net_1\, \wptr_gray_1[7]_net_1\, 
        \wptr_gray[8]_net_1\, \wptr_gray_1[8]_net_1\, 
        \wptr_gray[9]_net_1\, \wptr_gray_1[9]_net_1\, rdiff_bus, 
        \wptr_bin_sync[0]\, \wptr_bin_sync2[1]_net_1\, 
        \wptr_bin_sync[1]\, \wptr_bin_sync2[2]_net_1\, 
        \wptr_bin_sync[2]\, \wptr_bin_sync2[3]_net_1\, 
        \wptr_bin_sync[3]\, \wptr_bin_sync2[4]_net_1\, 
        \wptr_bin_sync[4]\, \wptr_bin_sync2[5]_net_1\, 
        \wptr_bin_sync[5]\, \wptr_bin_sync2[6]_net_1\, 
        \wptr_bin_sync[6]\, \rptr_bin_sync2[7]_net_1\, 
        \rptr_bin_sync[7]\, \rptr_bin_sync2[8]_net_1\, 
        \rptr_bin_sync[8]\, \rptr_bin_sync2[9]_net_1\, 
        \rptr_bin_sync[9]\, \rptr_bin_sync2[10]_net_1\, 
        \rptr_bin_sync[10]\, \rptr_bin_sync2[11]_net_1\, 
        \rptr_bin_sync[11]\, un1_we_p, \rptr_bin_sync2[0]_net_1\, 
        \rptr_bin_sync[0]\, \rptr_bin_sync2[1]_net_1\, 
        \rptr_bin_sync[1]\, \rptr_bin_sync2[2]_net_1\, 
        \rptr_bin_sync[2]\, \rptr_bin_sync2[3]_net_1\, 
        \rptr_bin_sync[3]\, \rptr_bin_sync2[4]_net_1\, 
        \rptr_bin_sync[4]\, \rptr_bin_sync2[5]_net_1\, 
        \rptr_bin_sync[5]\, \rptr_bin_sync2[6]_net_1\, 
        \rptr_bin_sync[6]\, \iRX_FIFO_Full_0\, fulli, 
        un2_re_p_i_i_a3_1, \iRX_FIFO_Empty_0\, empty_r_3, 
        \fifo_MEMWE\, \wptr[1]_net_1\, \wptr_s[1]\, 
        \wptr[2]_net_1\, \wptr_s[2]\, \wptr[3]_net_1\, 
        \wptr_s[3]\, \wptr[4]_net_1\, \wptr_s[4]\, 
        \wptr[5]_net_1\, \wptr_s[5]\, \wptr[6]_net_1\, 
        \wptr_s[6]\, \wptr[7]_net_1\, \wptr_s[7]\, 
        \wptr[8]_net_1\, \wptr_s[8]\, \wptr[9]_net_1\, 
        \wptr_s[9]\, \wptr[10]_net_1\, \wptr_s[10]\, 
        \wptr_s[11]_net_1\, \N_1005_i\, \fifo_MEMRADDR[1]\, 
        \memraddr_r_s[1]\, \fifo_MEMRADDR[2]\, \memraddr_r_s[2]\, 
        \fifo_MEMRADDR[3]\, \memraddr_r_s[3]\, \fifo_MEMRADDR[4]\, 
        \memraddr_r_s[4]\, \fifo_MEMRADDR[5]\, \memraddr_r_s[5]\, 
        \fifo_MEMRADDR[6]\, \memraddr_r_s[6]\, \fifo_MEMRADDR[7]\, 
        \memraddr_r_s[7]\, \fifo_MEMRADDR[8]\, \memraddr_r_s[8]\, 
        \fifo_MEMRADDR[9]\, \memraddr_r_s[9]\, 
        \fifo_MEMRADDR[10]\, \memraddr_r_s[10]_net_1\, 
        \fifo_MEMWADDR[0]\, \memwaddr_r_s[0]\, N_269, 
        \fifo_MEMWADDR[1]\, \memwaddr_r_s[1]\, \fifo_MEMWADDR[2]\, 
        \memwaddr_r_s[2]\, \fifo_MEMWADDR[3]\, \memwaddr_r_s[3]\, 
        \fifo_MEMWADDR[4]\, \memwaddr_r_s[4]\, \fifo_MEMWADDR[5]\, 
        \memwaddr_r_s[5]\, \fifo_MEMWADDR[6]\, \memwaddr_r_s[6]\, 
        \fifo_MEMWADDR[7]\, \memwaddr_r_s[7]\, \fifo_MEMWADDR[8]\, 
        \memwaddr_r_s[8]\, \fifo_MEMWADDR[9]\, \memwaddr_r_s[9]\, 
        \fifo_MEMWADDR[10]\, \memwaddr_r_s[10]_net_1\, 
        \rptr[1]_net_1\, \rptr_s[1]\, \rptr[2]_net_1\, 
        \rptr_s[2]\, \rptr[3]_net_1\, \rptr_s[3]\, 
        \rptr[4]_net_1\, \rptr_s[4]\, \rptr[5]_net_1\, 
        \rptr_s[5]\, \rptr[6]_net_1\, \rptr_s[6]\, 
        \rptr[7]_net_1\, \rptr_s[7]\, \rptr[8]_net_1\, 
        \rptr_s[8]\, \rptr[9]_net_1\, \rptr_s[9]\, 
        \rptr[10]_net_1\, \rptr_s[10]\, \rptr_s[11]_net_1\, 
        memwaddr_r_cry_cy, \memwaddr_r_cry[0]_net_1\, 
        \memwaddr_r_cry[1]_net_1\, \memwaddr_r_cry[2]_net_1\, 
        \memwaddr_r_cry[3]_net_1\, \memwaddr_r_cry[4]_net_1\, 
        \memwaddr_r_cry[5]_net_1\, \memwaddr_r_cry[6]_net_1\, 
        \memwaddr_r_cry[7]_net_1\, \memwaddr_r_cry[8]_net_1\, 
        \memwaddr_r_cry[9]_net_1\, \rdiff_bus_cry_0\, 
        rdiff_bus_cry_0_Y_2, \rdiff_bus_cry_1\, \rdiff_bus[1]\, 
        \rdiff_bus_cry_2\, \rdiff_bus[2]\, \rdiff_bus_cry_3\, 
        \rdiff_bus[3]\, \rdiff_bus_cry_4\, \rdiff_bus[4]\, 
        \rdiff_bus_cry_5\, \rdiff_bus[5]\, \rdiff_bus_cry_6\, 
        \rdiff_bus[6]\, \rdiff_bus_cry_7\, \rdiff_bus[7]\, 
        \rdiff_bus_cry_8\, \rdiff_bus[8]\, \rdiff_bus_cry_9\, 
        \rdiff_bus[9]\, \rdiff_bus[11]\, \rdiff_bus_cry_10\, 
        \rdiff_bus[10]\, \wdiff_bus_cry_0\, wdiff_bus_cry_0_Y_2, 
        \wdiff_bus_cry_1\, \wdiff_bus[1]\, \wdiff_bus_cry_2\, 
        \wdiff_bus[2]\, \wdiff_bus_cry_3\, \wdiff_bus[3]\, 
        \wdiff_bus_cry_4\, \wdiff_bus[4]\, \wdiff_bus_cry_5\, 
        \wdiff_bus[5]\, \wdiff_bus_cry_6\, \wdiff_bus[6]\, 
        \wdiff_bus_cry_7\, \wdiff_bus[7]\, \wdiff_bus_cry_8\, 
        \wdiff_bus[8]\, \wdiff_bus_cry_9\, \wdiff_bus[9]\, 
        \wdiff_bus[11]\, \wdiff_bus_cry_10\, \wdiff_bus[10]\, 
        rptr_s_377_FCO, \rptr_cry[1]_net_1\, \rptr_cry[2]_net_1\, 
        \rptr_cry[3]_net_1\, \rptr_cry[4]_net_1\, 
        \rptr_cry[5]_net_1\, \rptr_cry[6]_net_1\, 
        \rptr_cry[7]_net_1\, \rptr_cry[8]_net_1\, 
        \rptr_cry[9]_net_1\, \rptr_cry[10]_net_1\, 
        memraddr_r_s_378_FCO, \memraddr_r_cry[1]_net_1\, 
        \memraddr_r_cry[2]_net_1\, \memraddr_r_cry[3]_net_1\, 
        \memraddr_r_cry[4]_net_1\, \memraddr_r_cry[5]_net_1\, 
        \memraddr_r_cry[6]_net_1\, \memraddr_r_cry[7]_net_1\, 
        \memraddr_r_cry[8]_net_1\, \memraddr_r_cry[9]_net_1\, 
        wptr_s_379_FCO, \wptr_cry[1]_net_1\, \wptr_cry[2]_net_1\, 
        \wptr_cry[3]_net_1\, \wptr_cry[4]_net_1\, 
        \wptr_cry[5]_net_1\, \wptr_cry[6]_net_1\, 
        \wptr_cry[7]_net_1\, \wptr_cry[8]_net_1\, 
        \wptr_cry[9]_net_1\, \wptr_cry[10]_net_1\, 
        empty_r_3_0_a2_1, \fulli_0_a3_7\, \fulli_0_a3_6\, 
        empty_r_3_0_a2_7, empty_r_3_0_a2_9, \fulli_0_a3_8\, 
        empty_r_3_0_a2_5, \wptr_gray_sync[0]\, 
        \wptr_gray_sync[1]\, \wptr_gray_sync[2]\, 
        \wptr_gray_sync[3]\, \wptr_gray_sync[4]\, 
        \wptr_gray_sync[5]\, \wptr_gray_sync[6]\, 
        \wptr_gray_sync[7]\, \wptr_gray_sync[8]\, 
        \wptr_gray_sync[9]\, \wptr_gray_sync[10]\, 
        \rptr_gray_sync[0]\, \rptr_gray_sync[1]\, 
        \rptr_gray_sync[2]\, \rptr_gray_sync[3]\, 
        \rptr_gray_sync[4]\, \rptr_gray_sync[5]\, 
        \rptr_gray_sync[6]\, \rptr_gray_sync[7]\, 
        \rptr_gray_sync[8]\, \rptr_gray_sync[9]\, 
        \rptr_gray_sync[10]\ : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_4
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_4(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_2
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_2(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_1
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_1(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_3
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_3(DEF_ARCH);
begin 

    fifo_MEMWADDR(10) <= \fifo_MEMWADDR[10]\;
    fifo_MEMWADDR(9) <= \fifo_MEMWADDR[9]\;
    fifo_MEMWADDR(8) <= \fifo_MEMWADDR[8]\;
    fifo_MEMWADDR(7) <= \fifo_MEMWADDR[7]\;
    fifo_MEMWADDR(6) <= \fifo_MEMWADDR[6]\;
    fifo_MEMWADDR(5) <= \fifo_MEMWADDR[5]\;
    fifo_MEMWADDR(4) <= \fifo_MEMWADDR[4]\;
    fifo_MEMWADDR(3) <= \fifo_MEMWADDR[3]\;
    fifo_MEMWADDR(2) <= \fifo_MEMWADDR[2]\;
    fifo_MEMWADDR(1) <= \fifo_MEMWADDR[1]\;
    fifo_MEMWADDR(0) <= \fifo_MEMWADDR[0]\;
    fifo_MEMRADDR(10) <= \fifo_MEMRADDR[10]\;
    fifo_MEMRADDR(9) <= \fifo_MEMRADDR[9]\;
    fifo_MEMRADDR(8) <= \fifo_MEMRADDR[8]\;
    fifo_MEMRADDR(7) <= \fifo_MEMRADDR[7]\;
    fifo_MEMRADDR(6) <= \fifo_MEMRADDR[6]\;
    fifo_MEMRADDR(5) <= \fifo_MEMRADDR[5]\;
    fifo_MEMRADDR(4) <= \fifo_MEMRADDR[4]\;
    fifo_MEMRADDR(3) <= \fifo_MEMRADDR[3]\;
    fifo_MEMRADDR(2) <= \fifo_MEMRADDR[2]\;
    fifo_MEMRADDR(1) <= \fifo_MEMRADDR[1]\;
    fifo_MEMRADDR(0) <= \fifo_MEMRADDR[0]\;
    iRX_FIFO_Empty_0 <= \iRX_FIFO_Empty_0\;
    iRX_FIFO_Full_0 <= \iRX_FIFO_Full_0\;
    N_1005_i <= \N_1005_i\;
    fifo_MEMWE <= \fifo_MEMWE\;

    \rptr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[4]_net_1\, S
         => \rptr_s[5]\, Y => OPEN, FCO => \rptr_cry[5]_net_1\);
    
    wdiff_bus_cry_8 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[8]_net_1\, B => 
        \rptr_bin_sync2[8]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_7\, S => \wdiff_bus[8]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_8\);
    
    \wptr_gray[4]\ : SLE
      port map(D => \wptr_gray_1[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[4]_net_1\);
    
    \rptr_gray_1[3]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[3]_net_1\, B => \rptr[4]_net_1\, Y => 
        \rptr_gray_1[3]_net_1\);
    
    \rptr_bin_sync2[6]\ : SLE
      port map(D => \rptr_bin_sync[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[6]_net_1\);
    
    \rptr[1]\ : SLE
      port map(D => \rptr_s[1]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1005_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[1]_net_1\);
    
    \wptr_gray_1[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[9]_net_1\, B => \wptr[10]_net_1\, Y => 
        \wptr_gray_1[9]_net_1\);
    
    \rptr_gray_1[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[5]_net_1\, B => \rptr[6]_net_1\, Y => 
        \rptr_gray_1[5]_net_1\);
    
    \rptr_gray[9]\ : SLE
      port map(D => \rptr_gray_1[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[9]_net_1\);
    
    \rptr_gray[8]\ : SLE
      port map(D => \rptr_gray_1[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[8]_net_1\);
    
    \rptr_gray_1[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[2]_net_1\, B => \rptr[3]_net_1\, Y => 
        \rptr_gray_1[2]_net_1\);
    
    \rptr_bin_sync2[7]\ : SLE
      port map(D => \rptr_bin_sync[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[7]_net_1\);
    
    \memwaddr_r[1]\ : SLE
      port map(D => \memwaddr_r_s[1]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_269, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[1]\);
    
    \memwaddr_r_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[5]_net_1\, S => \memwaddr_r_s[6]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[6]_net_1\);
    
    \memwaddr_r_s[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[9]_net_1\, S => \memwaddr_r_s[10]_net_1\, 
        Y => OPEN, FCO => OPEN);
    
    \wptr_gray_1[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[7]_net_1\, B => \wptr[8]_net_1\, Y => 
        \wptr_gray_1[7]_net_1\);
    
    \memraddr_r[0]\ : SLE
      port map(D => \memraddr_r_s[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1005_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[0]\);
    
    \wptr[0]\ : SLE
      port map(D => \wptr_s[0]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[0]_net_1\);
    
    \rptr_bin_sync2[8]\ : SLE
      port map(D => \rptr_bin_sync[8]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[8]_net_1\);
    
    \rptr_gray_1[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[1]_net_1\, B => \rptr[2]_net_1\, Y => 
        \rptr_gray_1[1]_net_1\);
    
    \rptr_gray[10]\ : SLE
      port map(D => \rptr_gray_1[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[10]_net_1\);
    
    \wptr_gray_1[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[0]_net_1\, B => \wptr[1]_net_1\, Y => 
        \wptr_gray_1[0]_net_1\);
    
    wdiff_bus_cry_9 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[9]_net_1\, B => 
        \rptr_bin_sync2[9]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_8\, S => \wdiff_bus[9]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_9\);
    
    \rptr[5]\ : SLE
      port map(D => \rptr_s[5]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1005_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[5]_net_1\);
    
    \rptr_gray[3]\ : SLE
      port map(D => \rptr_gray_1[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[3]_net_1\);
    
    \rptr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[5]_net_1\, S
         => \rptr_s[6]\, Y => OPEN, FCO => \rptr_cry[6]_net_1\);
    
    \memwaddr_r_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[1]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[0]_net_1\, S => \memwaddr_r_s[1]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[1]_net_1\);
    
    \wptr_gray[3]\ : SLE
      port map(D => \wptr_gray_1[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[3]_net_1\);
    
    \rptr_gray_1[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[11]_net_1\, B => \rptr[10]_net_1\, Y
         => \rptr_gray_1[10]_net_1\);
    
    wdiff_bus_s_11 : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \rptr_bin_sync2[11]_net_1\, C
         => \wptr[11]_net_1\, D => GND_net_1, FCI => 
        \wdiff_bus_cry_10\, S => \wdiff_bus[11]\, Y => OPEN, FCO
         => OPEN);
    
    \rptr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[7]_net_1\, S
         => \rptr_s[8]\, Y => OPEN, FCO => \rptr_cry[8]_net_1\);
    
    \rptr[7]\ : SLE
      port map(D => \rptr_s[7]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1005_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[7]_net_1\);
    
    rdiff_bus_cry_4 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[4]_net_1\, B => 
        \rptr[4]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_3\, S => \rdiff_bus[4]\, Y => OPEN, FCO
         => \rdiff_bus_cry_4\);
    
    \rptr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[9]_net_1\, S
         => \rptr_s[10]\, Y => OPEN, FCO => \rptr_cry[10]_net_1\);
    
    fulli_0_a2_0_a2 : CFG3
      generic map(INIT => x"40")

      port map(A => ReadFIFO_Write_Ptr(0), B => N_1466, C => 
        ReadFIFO_Write_Ptr(1), Y => N_269);
    
    \rptr_bin_sync2[0]\ : SLE
      port map(D => \rptr_bin_sync[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[0]_net_1\);
    
    \L1.empty_r_3_0_a2_7\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \rdiff_bus[5]\, B => \rdiff_bus[6]\, C => 
        \rdiff_bus[7]\, D => \rdiff_bus[8]\, Y => 
        empty_r_3_0_a2_7);
    
    \wptr[11]\ : SLE
      port map(D => \wptr_s[11]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \wptr[11]_net_1\);
    
    rdiff_bus_cry_1 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[1]_net_1\, B => 
        \rptr[1]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_0\, S => \rdiff_bus[1]\, Y => OPEN, FCO
         => \rdiff_bus_cry_1\);
    
    \memraddr_r[1]\ : SLE
      port map(D => \memraddr_r_s[1]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1005_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[1]\);
    
    \L1.empty_r_3_0_a2_9\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \rdiff_bus[1]\, B => \rdiff_bus[2]\, C => 
        empty_r_3_0_a2_7, D => empty_r_3_0_a2_1, Y => 
        empty_r_3_0_a2_9);
    
    \rptr_bin_sync2[2]\ : SLE
      port map(D => \rptr_bin_sync[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[2]_net_1\);
    
    rdiff_bus_cry_6 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[6]_net_1\, B => 
        \rptr[6]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_5\, S => \rdiff_bus[6]\, Y => OPEN, FCO
         => \rdiff_bus_cry_6\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \memwaddr_r_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[3]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[2]_net_1\, S => \memwaddr_r_s[3]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[3]_net_1\);
    
    \rptr_gray[1]\ : SLE
      port map(D => \rptr_gray_1[1]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[1]_net_1\);
    
    \memwaddr_r[7]\ : SLE
      port map(D => \memwaddr_r_s[7]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_269, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[7]\);
    
    \memraddr_r_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[2]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[1]_net_1\, S => \memraddr_r_s[2]\, Y => 
        OPEN, FCO => \memraddr_r_cry[2]_net_1\);
    
    \wptr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[3]_net_1\, S
         => \wptr_s[4]\, Y => OPEN, FCO => \wptr_cry[4]_net_1\);
    
    empty_r_RNI2EM01 : CFG2
      generic map(INIT => x"2")

      port map(A => N_134, B => \iRX_FIFO_Empty_0\, Y => 
        \N_1005_i\);
    
    \memraddr_r_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[8]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[7]_net_1\, S => \memraddr_r_s[8]\, Y => 
        OPEN, FCO => \memraddr_r_cry[8]_net_1\);
    
    \wptr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[9]_net_1\, S
         => \wptr_s[10]\, Y => OPEN, FCO => \wptr_cry[10]_net_1\);
    
    wdiff_bus_cry_5 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[5]_net_1\, B => 
        \rptr_bin_sync2[5]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_4\, S => \wdiff_bus[5]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_5\);
    
    \memwaddr_r[4]\ : SLE
      port map(D => \memwaddr_r_s[4]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_269, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[4]\);
    
    memraddr_r_s_378 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[0]\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => memraddr_r_s_378_FCO);
    
    \wptr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[1]_net_1\, S
         => \wptr_s[2]\, Y => OPEN, FCO => \wptr_cry[2]_net_1\);
    
    wdiff_bus_cry_0 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[0]_net_1\, B => 
        \rptr_bin_sync2[0]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => VCC_net_1, S => OPEN, Y => wdiff_bus_cry_0_Y_2, 
        FCO => \wdiff_bus_cry_0\);
    
    \wptr[1]\ : SLE
      port map(D => \wptr_s[1]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[1]_net_1\);
    
    \rptr_bin_sync2[4]\ : SLE
      port map(D => \rptr_bin_sync[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[4]_net_1\);
    
    \wptr_bin_sync2[6]\ : SLE
      port map(D => \wptr_bin_sync[6]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[6]_net_1\);
    
    \memwaddr_r_cry_cy[0]\ : ARI1
      generic map(INIT => x"45500")

      port map(A => VCC_net_1, B => \iRX_FIFO_Full_0\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => memwaddr_r_cry_cy);
    
    \rptr[3]\ : SLE
      port map(D => \rptr_s[3]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1005_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[3]_net_1\);
    
    \wptr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[2]_net_1\, S
         => \wptr_s[3]\, Y => OPEN, FCO => \wptr_cry[3]_net_1\);
    
    \memwaddr_r_cry[0]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[0]\, C => 
        GND_net_1, D => GND_net_1, FCI => memwaddr_r_cry_cy, S
         => \memwaddr_r_s[0]\, Y => OPEN, FCO => 
        \memwaddr_r_cry[0]_net_1\);
    
    \rptr[6]\ : SLE
      port map(D => \rptr_s[6]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1005_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[6]_net_1\);
    
    rdiff_bus_cry_8 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[8]_net_1\, B => 
        \rptr[8]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_7\, S => \rdiff_bus[8]\, Y => OPEN, FCO
         => \rdiff_bus_cry_8\);
    
    \wptr_gray[10]\ : SLE
      port map(D => \wptr_gray_1[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[10]_net_1\);
    
    rdiff_bus_cry_7 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[7]_net_1\, B => 
        \rptr[7]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_6\, S => \rdiff_bus[7]\, Y => OPEN, FCO
         => \rdiff_bus_cry_7\);
    
    \wptr_bin_sync2[7]\ : SLE
      port map(D => \wptr_bin_sync[7]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[7]_net_1\);
    
    \rptr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[8]_net_1\, S
         => \rptr_s[9]\, Y => OPEN, FCO => \rptr_cry[9]_net_1\);
    
    \rptr_gray[5]\ : SLE
      port map(D => \rptr_gray_1[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[5]_net_1\);
    
    empty_r_RNI2KGB1_0 : CFG3
      generic map(INIT => x"A2")

      port map(A => REN_d1, B => N_134, C => \iRX_FIFO_Empty_0\, 
        Y => N_89_i);
    
    \wptr_gray_1[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[2]_net_1\, B => \wptr[3]_net_1\, Y => 
        \wptr_gray_1[2]_net_1\);
    
    \wptr[5]\ : SLE
      port map(D => \wptr_s[5]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[5]_net_1\);
    
    rdiff_bus_cry_5 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[5]_net_1\, B => 
        \rptr[5]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_4\, S => \rdiff_bus[5]\, Y => OPEN, FCO
         => \rdiff_bus_cry_5\);
    
    \wptr_bin_sync2[8]\ : SLE
      port map(D => \wptr_bin_sync[8]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[8]_net_1\);
    
    \wptr[7]\ : SLE
      port map(D => \wptr_s[7]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[7]_net_1\);
    
    empty_r_RNI2KGB1 : CFG3
      generic map(INIT => x"A6")

      port map(A => REN_d1, B => N_134, C => \iRX_FIFO_Empty_0\, 
        Y => N_155_i_i);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \wptr_gray[1]\ : SLE
      port map(D => \wptr_gray_1[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[1]_net_1\);
    
    \rptr_gray_1[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[9]_net_1\, B => \rptr[10]_net_1\, Y => 
        \rptr_gray_1[9]_net_1\);
    
    \rptr_bin_sync2[5]\ : SLE
      port map(D => \rptr_bin_sync[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[5]_net_1\);
    
    \rptr_bin_sync2[1]\ : SLE
      port map(D => \rptr_bin_sync[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[1]_net_1\);
    
    \memwaddr_r[10]\ : SLE
      port map(D => \memwaddr_r_s[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_269, ALn => irx_fifo_rst_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \fifo_MEMWADDR[10]\);
    
    wdiff_bus_cry_7 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[7]_net_1\, B => 
        \rptr_bin_sync2[7]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_6\, S => \wdiff_bus[7]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_7\);
    
    \wptr_bin_sync2[0]\ : SLE
      port map(D => \wptr_bin_sync[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rdiff_bus);
    
    \L1.un2_re_p_i_i_a3\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_134, B => \iRX_FIFO_Empty_0\, Y => 
        un2_re_p_i_i_a3_1);
    
    \L1.empty_r_3_0_a2_1\ : CFG2
      generic map(INIT => x"1")

      port map(A => \rdiff_bus[4]\, B => \rdiff_bus[3]\, Y => 
        empty_r_3_0_a2_1);
    
    rdiff_bus_s_11 : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \rptr[11]_net_1\, C => 
        \wptr_bin_sync2[11]_net_1\, D => GND_net_1, FCI => 
        \rdiff_bus_cry_10\, S => \rdiff_bus[11]\, Y => OPEN, FCO
         => OPEN);
    
    \memwaddr_r_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[8]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[7]_net_1\, S => \memwaddr_r_s[8]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[8]_net_1\);
    
    \wptr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => wptr_s_379_FCO, S => 
        \wptr_s[1]\, Y => OPEN, FCO => \wptr_cry[1]_net_1\);
    
    \memraddr_r[8]\ : SLE
      port map(D => \memraddr_r_s[8]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1005_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[8]\);
    
    \rptr[9]\ : SLE
      port map(D => \rptr_s[9]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1005_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[9]_net_1\);
    
    \wptr_gray_1[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[6]_net_1\, B => \wptr[7]_net_1\, Y => 
        \wptr_gray_1[6]_net_1\);
    
    \wptr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[6]_net_1\, S
         => \wptr_s[7]\, Y => OPEN, FCO => \wptr_cry[7]_net_1\);
    
    \wptr_bin_sync2[2]\ : SLE
      port map(D => \wptr_bin_sync[2]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[2]_net_1\);
    
    \rptr_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \rptr[0]_net_1\, Y => \rptr_s[0]\);
    
    \rptr[4]\ : SLE
      port map(D => \rptr_s[4]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1005_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[4]_net_1\);
    
    \memwaddr_r_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[4]_net_1\, S => \memwaddr_r_s[5]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[5]_net_1\);
    
    \memraddr_r_s[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[9]_net_1\, S => \memraddr_r_s[10]_net_1\, 
        Y => OPEN, FCO => OPEN);
    
    \wptr_gray[6]\ : SLE
      port map(D => \wptr_gray_1[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[6]_net_1\);
    
    \wptr_gray_1[3]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[3]_net_1\, B => \wptr[4]_net_1\, Y => 
        \wptr_gray_1[3]_net_1\);
    
    \wptr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[4]_net_1\, S
         => \wptr_s[5]\, Y => OPEN, FCO => \wptr_cry[5]_net_1\);
    
    \memraddr_r_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[4]_net_1\, S => \memraddr_r_s[5]\, Y => 
        OPEN, FCO => \memraddr_r_cry[5]_net_1\);
    
    \memraddr_r_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[1]\, C => 
        GND_net_1, D => GND_net_1, FCI => memraddr_r_s_378_FCO, S
         => \memraddr_r_s[1]\, Y => OPEN, FCO => 
        \memraddr_r_cry[1]_net_1\);
    
    \rptr_gray[4]\ : SLE
      port map(D => \rptr_gray_1[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[4]_net_1\);
    
    \wptr_bin_sync2[4]\ : SLE
      port map(D => \wptr_bin_sync[4]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[4]_net_1\);
    
    \wptr[3]\ : SLE
      port map(D => \wptr_s[3]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[3]_net_1\);
    
    \memwaddr_r[6]\ : SLE
      port map(D => \memwaddr_r_s[6]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_269, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[6]\);
    
    \wptr_s[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[10]_net_1\, S
         => \wptr_s[11]_net_1\, Y => OPEN, FCO => OPEN);
    
    \wptr[6]\ : SLE
      port map(D => \wptr_s[6]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[6]_net_1\);
    
    \memwaddr_r[9]\ : SLE
      port map(D => \memwaddr_r_s[9]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_269, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[9]\);
    
    \memraddr_r_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[3]_net_1\, S => \memraddr_r_s[4]\, Y => 
        OPEN, FCO => \memraddr_r_cry[4]_net_1\);
    
    \memraddr_r[10]\ : SLE
      port map(D => \memraddr_r_s[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1005_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[10]\);
    
    \memwaddr_r[3]\ : SLE
      port map(D => \memwaddr_r_s[3]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_269, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[3]\);
    
    full_r : SLE
      port map(D => fulli, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \iRX_FIFO_Full_0\);
    
    \rptr_bin_sync2[3]\ : SLE
      port map(D => \rptr_bin_sync[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[3]_net_1\);
    
    \wptr_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \wptr[0]_net_1\, Y => \wptr_s[0]\);
    
    \rptr[2]\ : SLE
      port map(D => \rptr_s[2]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1005_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[2]_net_1\);
    
    \memraddr_r[3]\ : SLE
      port map(D => \memraddr_r_s[3]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1005_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[3]\);
    
    \rptr_bin_sync2[9]\ : SLE
      port map(D => \rptr_bin_sync[9]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[9]_net_1\);
    
    \rptr[11]\ : SLE
      port map(D => \rptr_s[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1005_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rptr[11]_net_1\);
    
    \wptr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[5]_net_1\, S
         => \wptr_s[6]\, Y => OPEN, FCO => \wptr_cry[6]_net_1\);
    
    \rptr_bin_sync2[11]\ : SLE
      port map(D => \rptr_bin_sync[11]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[11]_net_1\);
    
    \wptr_bin_sync2[5]\ : SLE
      port map(D => \wptr_bin_sync[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[5]_net_1\);
    
    \wptr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[7]_net_1\, S
         => \wptr_s[8]\, Y => OPEN, FCO => \wptr_cry[8]_net_1\);
    
    \wptr_bin_sync2[1]\ : SLE
      port map(D => \wptr_bin_sync[1]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[1]_net_1\);
    
    \L1.un1_we_p_0_a3_0_a2\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_269, B => \iRX_FIFO_Full_0\, Y => un1_we_p);
    
    Wr_corefifo_grayToBinConv : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_4
      port map(wptr_bin_sync(11) => \wptr_bin_sync[11]\, 
        wptr_bin_sync(10) => \wptr_bin_sync[10]\, 
        wptr_bin_sync(9) => \wptr_bin_sync[9]\, wptr_bin_sync(8)
         => \wptr_bin_sync[8]\, wptr_bin_sync(7) => 
        \wptr_bin_sync[7]\, wptr_bin_sync(6) => 
        \wptr_bin_sync[6]\, wptr_bin_sync(5) => 
        \wptr_bin_sync[5]\, wptr_bin_sync(4) => 
        \wptr_bin_sync[4]\, wptr_bin_sync(3) => 
        \wptr_bin_sync[3]\, wptr_bin_sync(2) => 
        \wptr_bin_sync[2]\, wptr_bin_sync(1) => 
        \wptr_bin_sync[1]\, wptr_bin_sync(0) => 
        \wptr_bin_sync[0]\, wptr_gray_sync(10) => 
        \wptr_gray_sync[10]\, wptr_gray_sync(9) => 
        \wptr_gray_sync[9]\, wptr_gray_sync(8) => 
        \wptr_gray_sync[8]\, wptr_gray_sync(7) => 
        \wptr_gray_sync[7]\, wptr_gray_sync(6) => 
        \wptr_gray_sync[6]\, wptr_gray_sync(5) => 
        \wptr_gray_sync[5]\, wptr_gray_sync(4) => 
        \wptr_gray_sync[4]\, wptr_gray_sync(3) => 
        \wptr_gray_sync[3]\, wptr_gray_sync(2) => 
        \wptr_gray_sync[2]\, wptr_gray_sync(1) => 
        \wptr_gray_sync[1]\, wptr_gray_sync(0) => 
        \wptr_gray_sync[0]\);
    
    \wptr_gray_1[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[4]_net_1\, B => \wptr[5]_net_1\, Y => 
        \wptr_gray_1[4]_net_1\);
    
    wptr_s_379 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => wptr_s_379_FCO);
    
    overflow_r : SLE
      port map(D => un1_we_p, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        iRX_FIFO_OVERFLOW_0);
    
    fulli_0 : CFG4
      generic map(INIT => x"EAAA")

      port map(A => \wdiff_bus[11]\, B => \fulli_0_a3_7\, C => 
        N_269, D => \fulli_0_a3_8\, Y => fulli);
    
    \memraddr_r_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \fifo_MEMRADDR[0]\, Y => \memraddr_r_s[0]\);
    
    \rptr_gray[11]\ : SLE
      port map(D => \rptr[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[11]_net_1\);
    
    \wptr_bin_sync2[10]\ : SLE
      port map(D => \wptr_bin_sync[10]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[10]_net_1\);
    
    \rptr[10]\ : SLE
      port map(D => \rptr_s[10]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1005_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rptr[10]_net_1\);
    
    \wptr[9]\ : SLE
      port map(D => \wptr_s[9]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[9]_net_1\);
    
    Wr_corefifo_doubleSync : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_2
      port map(wptr_gray(11) => \wptr_gray[11]_net_1\, 
        wptr_gray(10) => \wptr_gray[10]_net_1\, wptr_gray(9) => 
        \wptr_gray[9]_net_1\, wptr_gray(8) => 
        \wptr_gray[8]_net_1\, wptr_gray(7) => 
        \wptr_gray[7]_net_1\, wptr_gray(6) => 
        \wptr_gray[6]_net_1\, wptr_gray(5) => 
        \wptr_gray[5]_net_1\, wptr_gray(4) => 
        \wptr_gray[4]_net_1\, wptr_gray(3) => 
        \wptr_gray[3]_net_1\, wptr_gray(2) => 
        \wptr_gray[2]_net_1\, wptr_gray(1) => 
        \wptr_gray[1]_net_1\, wptr_gray(0) => 
        \wptr_gray[0]_net_1\, wptr_gray_sync(10) => 
        \wptr_gray_sync[10]\, wptr_gray_sync(9) => 
        \wptr_gray_sync[9]\, wptr_gray_sync(8) => 
        \wptr_gray_sync[8]\, wptr_gray_sync(7) => 
        \wptr_gray_sync[7]\, wptr_gray_sync(6) => 
        \wptr_gray_sync[6]\, wptr_gray_sync(5) => 
        \wptr_gray_sync[5]\, wptr_gray_sync(4) => 
        \wptr_gray_sync[4]\, wptr_gray_sync(3) => 
        \wptr_gray_sync[3]\, wptr_gray_sync(2) => 
        \wptr_gray_sync[2]\, wptr_gray_sync(1) => 
        \wptr_gray_sync[1]\, wptr_gray_sync(0) => 
        \wptr_gray_sync[0]\, wptr_bin_sync_0 => 
        \wptr_bin_sync[11]\, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, irx_fifo_rst_i => 
        irx_fifo_rst_i);
    
    \rptr_gray[0]\ : SLE
      port map(D => \rptr_gray_1[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[0]_net_1\);
    
    empty_r : SLE
      port map(D => empty_r_3, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \iRX_FIFO_Empty_0\);
    
    \rptr_gray_1[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[7]_net_1\, B => \rptr[8]_net_1\, Y => 
        \rptr_gray_1[7]_net_1\);
    
    \wptr[4]\ : SLE
      port map(D => \wptr_s[4]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[4]_net_1\);
    
    \memwaddr_r[8]\ : SLE
      port map(D => \memwaddr_r_s[8]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_269, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[8]\);
    
    \memwaddr_r[2]\ : SLE
      port map(D => \memwaddr_r_s[2]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_269, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[2]\);
    
    \L1.empty_r_3_0_a2_5\ : CFG3
      generic map(INIT => x"0E")

      port map(A => N_134, B => rdiff_bus_cry_0_Y_2, C => 
        \rdiff_bus[11]\, Y => empty_r_3_0_a2_5);
    
    \wptr_bin_sync2[11]\ : SLE
      port map(D => \wptr_bin_sync[11]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[11]_net_1\);
    
    \wptr_gray_1[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[1]_net_1\, B => \wptr[2]_net_1\, Y => 
        \wptr_gray_1[1]_net_1\);
    
    underflow_r : SLE
      port map(D => un2_re_p_i_i_a3_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => iRX_FIFO_UNDERRUN_0);
    
    fulli_0_a3_7 : CFG4
      generic map(INIT => x"8000")

      port map(A => \wdiff_bus[6]\, B => \wdiff_bus[7]\, C => 
        \wdiff_bus[8]\, D => \wdiff_bus[9]\, Y => \fulli_0_a3_7\);
    
    \memwaddr_r_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[6]_net_1\, S => \memwaddr_r_s[7]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[7]_net_1\);
    
    \wptr_gray[5]\ : SLE
      port map(D => \wptr_gray_1[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[5]_net_1\);
    
    \memraddr_r[7]\ : SLE
      port map(D => \memraddr_r_s[7]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1005_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[7]\);
    
    \rptr_bin_sync2[10]\ : SLE
      port map(D => \rptr_bin_sync[10]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[10]_net_1\);
    
    wdiff_bus_cry_10 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[10]_net_1\, B => 
        \rptr_bin_sync2[10]_net_1\, C => GND_net_1, D => 
        GND_net_1, FCI => \wdiff_bus_cry_9\, S => \wdiff_bus[10]\, 
        Y => OPEN, FCO => \wdiff_bus_cry_10\);
    
    \memwaddr_r_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[9]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[8]_net_1\, S => \memwaddr_r_s[9]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[9]_net_1\);
    
    \wptr_gray[8]\ : SLE
      port map(D => \wptr_gray_1[8]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[8]_net_1\);
    
    \wptr_gray[7]\ : SLE
      port map(D => \wptr_gray_1[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[7]_net_1\);
    
    \wptr_gray_1[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[5]_net_1\, B => \wptr[6]_net_1\, Y => 
        \wptr_gray_1[5]_net_1\);
    
    \memwaddr_r[5]\ : SLE
      port map(D => \memwaddr_r_s[5]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_269, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[5]\);
    
    \L1.empty_r_3_0_a2\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \rdiff_bus[9]\, B => \rdiff_bus[10]\, C => 
        empty_r_3_0_a2_5, D => empty_r_3_0_a2_9, Y => empty_r_3);
    
    \rptr[8]\ : SLE
      port map(D => \rptr_s[8]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1005_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[8]_net_1\);
    
    Rd_corefifo_doubleSync : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_1
      port map(rptr_gray(11) => \rptr_gray[11]_net_1\, 
        rptr_gray(10) => \rptr_gray[10]_net_1\, rptr_gray(9) => 
        \rptr_gray[9]_net_1\, rptr_gray(8) => 
        \rptr_gray[8]_net_1\, rptr_gray(7) => 
        \rptr_gray[7]_net_1\, rptr_gray(6) => 
        \rptr_gray[6]_net_1\, rptr_gray(5) => 
        \rptr_gray[5]_net_1\, rptr_gray(4) => 
        \rptr_gray[4]_net_1\, rptr_gray(3) => 
        \rptr_gray[3]_net_1\, rptr_gray(2) => 
        \rptr_gray[2]_net_1\, rptr_gray(1) => 
        \rptr_gray[1]_net_1\, rptr_gray(0) => 
        \rptr_gray[0]_net_1\, rptr_gray_sync(10) => 
        \rptr_gray_sync[10]\, rptr_gray_sync(9) => 
        \rptr_gray_sync[9]\, rptr_gray_sync(8) => 
        \rptr_gray_sync[8]\, rptr_gray_sync(7) => 
        \rptr_gray_sync[7]\, rptr_gray_sync(6) => 
        \rptr_gray_sync[6]\, rptr_gray_sync(5) => 
        \rptr_gray_sync[5]\, rptr_gray_sync(4) => 
        \rptr_gray_sync[4]\, rptr_gray_sync(3) => 
        \rptr_gray_sync[3]\, rptr_gray_sync(2) => 
        \rptr_gray_sync[2]\, rptr_gray_sync(1) => 
        \rptr_gray_sync[1]\, rptr_gray_sync(0) => 
        \rptr_gray_sync[0]\, rptr_bin_sync_0 => 
        \rptr_bin_sync[11]\, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, irx_fifo_rst_i => irx_fifo_rst_i);
    
    \rptr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[3]_net_1\, S
         => \rptr_s[4]\, Y => OPEN, FCO => \rptr_cry[4]_net_1\);
    
    wdiff_bus_cry_2 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[2]_net_1\, B => 
        \rptr_bin_sync2[2]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_1\, S => \wdiff_bus[2]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_2\);
    
    \rptr_gray[2]\ : SLE
      port map(D => \rptr_gray_1[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[2]_net_1\);
    
    \wptr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[8]_net_1\, S
         => \wptr_s[9]\, Y => OPEN, FCO => \wptr_cry[9]_net_1\);
    
    \wptr_bin_sync2[3]\ : SLE
      port map(D => \wptr_bin_sync[3]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[3]_net_1\);
    
    \wptr[2]\ : SLE
      port map(D => \wptr_s[2]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[2]_net_1\);
    
    \rptr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[1]_net_1\, S
         => \rptr_s[2]\, Y => OPEN, FCO => \rptr_cry[2]_net_1\);
    
    rdiff_bus_cry_9 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[9]_net_1\, B => 
        \rptr[9]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_8\, S => \rdiff_bus[9]\, Y => OPEN, FCO
         => \rdiff_bus_cry_9\);
    
    \memwaddr_r[0]\ : SLE
      port map(D => \memwaddr_r_s[0]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_269, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[0]\);
    
    \wptr_gray[2]\ : SLE
      port map(D => \wptr_gray_1[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[2]_net_1\);
    
    wdiff_bus_cry_4 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[4]_net_1\, B => 
        \rptr_bin_sync2[4]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_3\, S => \wdiff_bus[4]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_4\);
    
    \memwaddr_r_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[2]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[1]_net_1\, S => \memwaddr_r_s[2]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[2]_net_1\);
    
    \wptr_gray[11]\ : SLE
      port map(D => \wptr[11]_net_1\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr_gray[11]_net_1\);
    
    \wptr_bin_sync2[9]\ : SLE
      port map(D => \wptr_bin_sync[9]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[9]_net_1\);
    
    rptr_s_377 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => rptr_s_377_FCO);
    
    \rptr_gray_1[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[6]_net_1\, B => \rptr[7]_net_1\, Y => 
        \rptr_gray_1[6]_net_1\);
    
    \wptr_gray_1[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[11]_net_1\, B => \wptr[10]_net_1\, Y
         => \wptr_gray_1[10]_net_1\);
    
    wdiff_bus_cry_6 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[6]_net_1\, B => 
        \rptr_bin_sync2[6]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_5\, S => \wdiff_bus[6]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_6\);
    
    \rptr_s[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[10]_net_1\, S
         => \rptr_s[11]_net_1\, Y => OPEN, FCO => OPEN);
    
    \rptr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[2]_net_1\, S
         => \rptr_s[3]\, Y => OPEN, FCO => \rptr_cry[3]_net_1\);
    
    \memraddr_r[4]\ : SLE
      port map(D => \memraddr_r_s[4]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1005_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[4]\);
    
    \memraddr_r_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[6]_net_1\, S => \memraddr_r_s[7]\, Y => 
        OPEN, FCO => \memraddr_r_cry[7]_net_1\);
    
    memwe_0_a3_0_a2 : CFG4
      generic map(INIT => x"0020")

      port map(A => ReadFIFO_Write_Ptr(1), B => \iRX_FIFO_Full_0\, 
        C => N_1466, D => ReadFIFO_Write_Ptr(0), Y => 
        \fifo_MEMWE\);
    
    \memraddr_r_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[9]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[8]_net_1\, S => \memraddr_r_s[9]\, Y => 
        OPEN, FCO => \memraddr_r_cry[9]_net_1\);
    
    \memraddr_r[5]\ : SLE
      port map(D => \memraddr_r_s[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1005_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[5]\);
    
    \rptr_gray[6]\ : SLE
      port map(D => \rptr_gray_1[6]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[6]_net_1\);
    
    \memraddr_r[9]\ : SLE
      port map(D => \memraddr_r_s[9]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1005_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[9]\);
    
    \rptr[0]\ : SLE
      port map(D => \rptr_s[0]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1005_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[0]_net_1\);
    
    fulli_0_a3_6 : CFG4
      generic map(INIT => x"8000")

      port map(A => \wdiff_bus[2]\, B => \wdiff_bus[3]\, C => 
        \wdiff_bus[5]\, D => \wdiff_bus[4]\, Y => \fulli_0_a3_6\);
    
    \wptr[10]\ : SLE
      port map(D => \wptr_s[10]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[10]_net_1\);
    
    \memwaddr_r_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[3]_net_1\, S => \memwaddr_r_s[4]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[4]_net_1\);
    
    \memraddr_r_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[3]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[2]_net_1\, S => \memraddr_r_s[3]\, Y => 
        OPEN, FCO => \memraddr_r_cry[3]_net_1\);
    
    wdiff_bus_cry_1 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[1]_net_1\, B => 
        \rptr_bin_sync2[1]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_0\, S => \wdiff_bus[1]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_1\);
    
    rdiff_bus_cry_2 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[2]_net_1\, B => 
        \rptr[2]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_1\, S => \rdiff_bus[2]\, Y => OPEN, FCO
         => \rdiff_bus_cry_2\);
    
    \wptr_gray[9]\ : SLE
      port map(D => \wptr_gray_1[9]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[9]_net_1\);
    
    \rptr_gray_1[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[4]_net_1\, B => \rptr[5]_net_1\, Y => 
        \rptr_gray_1[4]_net_1\);
    
    \wptr_gray_1[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[8]_net_1\, B => \wptr[9]_net_1\, Y => 
        \wptr_gray_1[8]_net_1\);
    
    Rd_corefifo_grayToBinConv : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_3
      port map(rptr_bin_sync(11) => \rptr_bin_sync[11]\, 
        rptr_bin_sync(10) => \rptr_bin_sync[10]\, 
        rptr_bin_sync(9) => \rptr_bin_sync[9]\, rptr_bin_sync(8)
         => \rptr_bin_sync[8]\, rptr_bin_sync(7) => 
        \rptr_bin_sync[7]\, rptr_bin_sync(6) => 
        \rptr_bin_sync[6]\, rptr_bin_sync(5) => 
        \rptr_bin_sync[5]\, rptr_bin_sync(4) => 
        \rptr_bin_sync[4]\, rptr_bin_sync(3) => 
        \rptr_bin_sync[3]\, rptr_bin_sync(2) => 
        \rptr_bin_sync[2]\, rptr_bin_sync(1) => 
        \rptr_bin_sync[1]\, rptr_bin_sync(0) => 
        \rptr_bin_sync[0]\, rptr_gray_sync(10) => 
        \rptr_gray_sync[10]\, rptr_gray_sync(9) => 
        \rptr_gray_sync[9]\, rptr_gray_sync(8) => 
        \rptr_gray_sync[8]\, rptr_gray_sync(7) => 
        \rptr_gray_sync[7]\, rptr_gray_sync(6) => 
        \rptr_gray_sync[6]\, rptr_gray_sync(5) => 
        \rptr_gray_sync[5]\, rptr_gray_sync(4) => 
        \rptr_gray_sync[4]\, rptr_gray_sync(3) => 
        \rptr_gray_sync[3]\, rptr_gray_sync(2) => 
        \rptr_gray_sync[2]\, rptr_gray_sync(1) => 
        \rptr_gray_sync[1]\, rptr_gray_sync(0) => 
        \rptr_gray_sync[0]\);
    
    \rptr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => rptr_s_377_FCO, S => 
        \rptr_s[1]\, Y => OPEN, FCO => \rptr_cry[1]_net_1\);
    
    rdiff_bus_cry_3 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[3]_net_1\, B => 
        \rptr[3]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_2\, S => \rdiff_bus[3]\, Y => OPEN, FCO
         => \rdiff_bus_cry_3\);
    
    rdiff_bus_cry_10 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[10]_net_1\, B => 
        \rptr[10]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_9\, S => \rdiff_bus[10]\, Y => OPEN, FCO
         => \rdiff_bus_cry_10\);
    
    \memraddr_r_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[5]_net_1\, S => \memraddr_r_s[6]\, Y => 
        OPEN, FCO => \memraddr_r_cry[6]_net_1\);
    
    \memraddr_r[6]\ : SLE
      port map(D => \memraddr_r_s[6]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1005_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[6]\);
    
    \rptr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[6]_net_1\, S
         => \rptr_s[7]\, Y => OPEN, FCO => \rptr_cry[7]_net_1\);
    
    rdiff_bus_cry_0 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => rdiff_bus, B => \rptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => rdiff_bus_cry_0_Y_2, FCO => \rdiff_bus_cry_0\);
    
    \memraddr_r[2]\ : SLE
      port map(D => \memraddr_r_s[2]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1005_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[2]\);
    
    \wptr[8]\ : SLE
      port map(D => \wptr_s[8]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[8]_net_1\);
    
    wdiff_bus_cry_3 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[3]_net_1\, B => 
        \rptr_bin_sync2[3]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_2\, S => \wdiff_bus[3]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_3\);
    
    fulli_0_a3_8 : CFG4
      generic map(INIT => x"4000")

      port map(A => wdiff_bus_cry_0_Y_2, B => \wdiff_bus[1]\, C
         => \wdiff_bus[10]\, D => \fulli_0_a3_6\, Y => 
        \fulli_0_a3_8\);
    
    \rptr_gray[7]\ : SLE
      port map(D => \rptr_gray_1[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[7]_net_1\);
    
    \wptr_gray[0]\ : SLE
      port map(D => \wptr_gray_1[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[0]_net_1\);
    
    \rptr_gray_1[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[0]_net_1\, B => \rptr[1]_net_1\, Y => 
        \rptr_gray_1[0]_net_1\);
    
    \rptr_gray_1[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[8]_net_1\, B => \rptr[9]_net_1\, Y => 
        \rptr_gray_1[8]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_1 is

    port( RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          ReadFIFO_Write_Ptr        : in    std_logic_vector(1 downto 0);
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          RX_FIFO_DOUT_2_0          : out   std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          N_1466                    : in    std_logic;
          N_667                     : out   std_logic;
          N_669                     : out   std_logic;
          N_716                     : out   std_logic;
          N_670                     : out   std_logic;
          N_668                     : out   std_logic;
          N_666                     : out   std_logic;
          N_665                     : out   std_logic;
          N_664                     : out   std_logic;
          N_134                     : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          irx_fifo_rst_i            : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_1;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_1 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_1
    port( RDATA_int                 : out   std_logic_vector(8 downto 0);
          fifo_MEMRADDR             : in    std_logic_vector(10 downto 0) := (others => 'U');
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          fifo_MEMWADDR             : in    std_logic_vector(10 downto 0) := (others => 'U');
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          N_1005_i                  : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          fifo_MEMWE                : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_1
    port( ReadFIFO_Write_Ptr        : in    std_logic_vector(1 downto 0) := (others => 'U');
          fifo_MEMWADDR             : out   std_logic_vector(10 downto 0);
          fifo_MEMRADDR             : out   std_logic_vector(10 downto 0);
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          N_155_i_i                 : out   std_logic;
          N_89_i                    : out   std_logic;
          REN_d1                    : in    std_logic := 'U';
          N_134                     : in    std_logic := 'U';
          N_1466                    : in    std_logic := 'U';
          N_1005_i                  : out   std_logic;
          fifo_MEMWE                : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          irx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \RDATA_r[4]_net_1\, VCC_net_1, \RDATA_int[4]\, N_89_i, 
        GND_net_1, \RDATA_r[5]_net_1\, \RDATA_int[5]\, 
        \RDATA_r[6]_net_1\, \RDATA_int[6]\, \RDATA_r[7]_net_1\, 
        \RDATA_int[7]\, \RDATA_r[8]_net_1\, \RDATA_int[8]\, 
        \re_set\, \REN_d1\, N_155_i_i, \RDATA_r[0]_net_1\, 
        \RDATA_int[0]\, \RDATA_r[1]_net_1\, \RDATA_int[1]\, 
        \RDATA_r[2]_net_1\, \RDATA_int[2]\, \RDATA_r[3]_net_1\, 
        \RDATA_int[3]\, N_1005_i, \RE_d1\, \re_pulse_d1\, 
        \re_pulse\, \iRX_FIFO_Empty_0\, \fifo_MEMWADDR[0]\, 
        \fifo_MEMWADDR[1]\, \fifo_MEMWADDR[2]\, 
        \fifo_MEMWADDR[3]\, \fifo_MEMWADDR[4]\, 
        \fifo_MEMWADDR[5]\, \fifo_MEMWADDR[6]\, 
        \fifo_MEMWADDR[7]\, \fifo_MEMWADDR[8]\, 
        \fifo_MEMWADDR[9]\, \fifo_MEMWADDR[10]\, 
        \fifo_MEMRADDR[0]\, \fifo_MEMRADDR[1]\, 
        \fifo_MEMRADDR[2]\, \fifo_MEMRADDR[3]\, 
        \fifo_MEMRADDR[4]\, \fifo_MEMRADDR[5]\, 
        \fifo_MEMRADDR[6]\, \fifo_MEMRADDR[7]\, 
        \fifo_MEMRADDR[8]\, \fifo_MEMRADDR[9]\, 
        \fifo_MEMRADDR[10]\, fifo_MEMWE : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_1
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_1(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_1
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_1(DEF_ARCH);
begin 

    iRX_FIFO_Empty_0 <= \iRX_FIFO_Empty_0\;

    re_pulse : CFG4
      generic map(INIT => x"FAF2")

      port map(A => \REN_d1\, B => N_134, C => \re_set\, D => 
        \iRX_FIFO_Empty_0\, Y => \re_pulse\);
    
    \RDATA_r[3]\ : SLE
      port map(D => \RDATA_int[3]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[3]_net_1\);
    
    \Q_i_m2[2]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[2]_net_1\, C => 
        \RDATA_int[2]\, D => \RE_d1\, Y => N_665);
    
    re_pulse_d1 : SLE
      port map(D => \re_pulse\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \re_pulse_d1\);
    
    \RDATA_r[5]\ : SLE
      port map(D => \RDATA_int[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[5]_net_1\);
    
    \Q_i_m2[0]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[0]_net_1\, C => 
        \RDATA_int[0]\, D => \RE_d1\, Y => N_664);
    
    \Q_i_m2[3]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[3]_net_1\, C => 
        \RDATA_int[3]\, D => \RE_d1\, Y => N_666);
    
    \RDATA_r[8]\ : SLE
      port map(D => \RDATA_int[8]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[8]_net_1\);
    
    \Q_i_m2[7]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[7]_net_1\, C => 
        \RDATA_int[7]\, D => \RE_d1\, Y => N_670);
    
    \Q_i_m2[6]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[6]_net_1\, C => 
        \RDATA_int[6]\, D => \RE_d1\, Y => N_669);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \RW1.UI_ram_wrapper_1\ : FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_1
      port map(RDATA_int(8) => \RDATA_int[8]\, RDATA_int(7) => 
        \RDATA_int[7]\, RDATA_int(6) => \RDATA_int[6]\, 
        RDATA_int(5) => \RDATA_int[5]\, RDATA_int(4) => 
        \RDATA_int[4]\, RDATA_int(3) => \RDATA_int[3]\, 
        RDATA_int(2) => \RDATA_int[2]\, RDATA_int(1) => 
        \RDATA_int[1]\, RDATA_int(0) => \RDATA_int[0]\, 
        fifo_MEMRADDR(10) => \fifo_MEMRADDR[10]\, 
        fifo_MEMRADDR(9) => \fifo_MEMRADDR[9]\, fifo_MEMRADDR(8)
         => \fifo_MEMRADDR[8]\, fifo_MEMRADDR(7) => 
        \fifo_MEMRADDR[7]\, fifo_MEMRADDR(6) => 
        \fifo_MEMRADDR[6]\, fifo_MEMRADDR(5) => 
        \fifo_MEMRADDR[5]\, fifo_MEMRADDR(4) => 
        \fifo_MEMRADDR[4]\, fifo_MEMRADDR(3) => 
        \fifo_MEMRADDR[3]\, fifo_MEMRADDR(2) => 
        \fifo_MEMRADDR[2]\, fifo_MEMRADDR(1) => 
        \fifo_MEMRADDR[1]\, fifo_MEMRADDR(0) => 
        \fifo_MEMRADDR[0]\, RX_FIFO_DIN_pipe(8) => 
        RX_FIFO_DIN_pipe(8), RX_FIFO_DIN_pipe(7) => 
        RX_FIFO_DIN_pipe(7), RX_FIFO_DIN_pipe(6) => 
        RX_FIFO_DIN_pipe(6), RX_FIFO_DIN_pipe(5) => 
        RX_FIFO_DIN_pipe(5), RX_FIFO_DIN_pipe(4) => 
        RX_FIFO_DIN_pipe(4), RX_FIFO_DIN_pipe(3) => 
        RX_FIFO_DIN_pipe(3), RX_FIFO_DIN_pipe(2) => 
        RX_FIFO_DIN_pipe(2), RX_FIFO_DIN_pipe(1) => 
        RX_FIFO_DIN_pipe(1), RX_FIFO_DIN_pipe(0) => 
        RX_FIFO_DIN_pipe(0), fifo_MEMWADDR(10) => 
        \fifo_MEMWADDR[10]\, fifo_MEMWADDR(9) => 
        \fifo_MEMWADDR[9]\, fifo_MEMWADDR(8) => 
        \fifo_MEMWADDR[8]\, fifo_MEMWADDR(7) => 
        \fifo_MEMWADDR[7]\, fifo_MEMWADDR(6) => 
        \fifo_MEMWADDR[6]\, fifo_MEMWADDR(5) => 
        \fifo_MEMWADDR[5]\, fifo_MEMWADDR(4) => 
        \fifo_MEMWADDR[4]\, fifo_MEMWADDR(3) => 
        \fifo_MEMWADDR[3]\, fifo_MEMWADDR(2) => 
        \fifo_MEMWADDR[2]\, fifo_MEMWADDR(1) => 
        \fifo_MEMWADDR[1]\, fifo_MEMWADDR(0) => 
        \fifo_MEMWADDR[0]\, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, N_1005_i => N_1005_i, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, fifo_MEMWE
         => fifo_MEMWE);
    
    \RDATA_r[0]\ : SLE
      port map(D => \RDATA_int[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[0]_net_1\);
    
    \Q_i_m2[5]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[5]_net_1\, C => 
        \RDATA_int[5]\, D => \RE_d1\, Y => N_668);
    
    \RDATA_r[2]\ : SLE
      port map(D => \RDATA_int[2]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[2]_net_1\);
    
    \RDATA_r[6]\ : SLE
      port map(D => \RDATA_int[6]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[6]_net_1\);
    
    \L31.U_corefifo_async\ : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_1
      port map(ReadFIFO_Write_Ptr(1) => ReadFIFO_Write_Ptr(1), 
        ReadFIFO_Write_Ptr(0) => ReadFIFO_Write_Ptr(0), 
        fifo_MEMWADDR(10) => \fifo_MEMWADDR[10]\, 
        fifo_MEMWADDR(9) => \fifo_MEMWADDR[9]\, fifo_MEMWADDR(8)
         => \fifo_MEMWADDR[8]\, fifo_MEMWADDR(7) => 
        \fifo_MEMWADDR[7]\, fifo_MEMWADDR(6) => 
        \fifo_MEMWADDR[6]\, fifo_MEMWADDR(5) => 
        \fifo_MEMWADDR[5]\, fifo_MEMWADDR(4) => 
        \fifo_MEMWADDR[4]\, fifo_MEMWADDR(3) => 
        \fifo_MEMWADDR[3]\, fifo_MEMWADDR(2) => 
        \fifo_MEMWADDR[2]\, fifo_MEMWADDR(1) => 
        \fifo_MEMWADDR[1]\, fifo_MEMWADDR(0) => 
        \fifo_MEMWADDR[0]\, fifo_MEMRADDR(10) => 
        \fifo_MEMRADDR[10]\, fifo_MEMRADDR(9) => 
        \fifo_MEMRADDR[9]\, fifo_MEMRADDR(8) => 
        \fifo_MEMRADDR[8]\, fifo_MEMRADDR(7) => 
        \fifo_MEMRADDR[7]\, fifo_MEMRADDR(6) => 
        \fifo_MEMRADDR[6]\, fifo_MEMRADDR(5) => 
        \fifo_MEMRADDR[5]\, fifo_MEMRADDR(4) => 
        \fifo_MEMRADDR[4]\, fifo_MEMRADDR(3) => 
        \fifo_MEMRADDR[3]\, fifo_MEMRADDR(2) => 
        \fifo_MEMRADDR[2]\, fifo_MEMRADDR(1) => 
        \fifo_MEMRADDR[1]\, fifo_MEMRADDR(0) => 
        \fifo_MEMRADDR[0]\, iRX_FIFO_Empty_0 => 
        \iRX_FIFO_Empty_0\, iRX_FIFO_UNDERRUN_0 => 
        iRX_FIFO_UNDERRUN_0, iRX_FIFO_Full_0 => iRX_FIFO_Full_0, 
        iRX_FIFO_OVERFLOW_0 => iRX_FIFO_OVERFLOW_0, N_155_i_i => 
        N_155_i_i, N_89_i => N_89_i, REN_d1 => \REN_d1\, N_134
         => N_134, N_1466 => N_1466, N_1005_i => N_1005_i, 
        fifo_MEMWE => fifo_MEMWE, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, irx_fifo_rst_i => irx_fifo_rst_i);
    
    re_set : SLE
      port map(D => \REN_d1\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => N_155_i_i, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \re_set\);
    
    \Q_i_m2[8]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[8]_net_1\, C => 
        \RDATA_int[8]\, D => \RE_d1\, Y => N_716);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    RE_d1 : SLE
      port map(D => N_134, CLK => m2s010_som_sb_0_CCC_71MHz, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \RE_d1\);
    
    \RDATA_r[7]\ : SLE
      port map(D => \RDATA_int[7]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[7]_net_1\);
    
    \RDATA_r[4]\ : SLE
      port map(D => \RDATA_int[4]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[4]_net_1\);
    
    \Q[1]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[1]_net_1\, C => 
        \RDATA_int[1]\, D => \RE_d1\, Y => RX_FIFO_DOUT_2_0);
    
    REN_d1 : SLE
      port map(D => N_1005_i, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \REN_d1\);
    
    \Q_i_m2[4]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[4]_net_1\, C => 
        \RDATA_int[4]\, D => \RE_d1\, Y => N_667);
    
    \RDATA_r[1]\ : SLE
      port map(D => \RDATA_int[1]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[1]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_1 is

    port( ReadFIFO_Write_Ptr        : in    std_logic_vector(1 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          RX_FIFO_DOUT_2_0          : out   std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          irx_fifo_rst_i            : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          N_134                     : in    std_logic;
          N_664                     : out   std_logic;
          N_665                     : out   std_logic;
          N_666                     : out   std_logic;
          N_668                     : out   std_logic;
          N_670                     : out   std_logic;
          N_716                     : out   std_logic;
          N_669                     : out   std_logic;
          N_667                     : out   std_logic;
          N_1466                    : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic
        );

end FIFO_8Kx9_1;

architecture DEF_ARCH of FIFO_8Kx9_1 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_1
    port( RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          ReadFIFO_Write_Ptr        : in    std_logic_vector(1 downto 0) := (others => 'U');
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          RX_FIFO_DOUT_2_0          : out   std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          N_1466                    : in    std_logic := 'U';
          N_667                     : out   std_logic;
          N_669                     : out   std_logic;
          N_716                     : out   std_logic;
          N_670                     : out   std_logic;
          N_668                     : out   std_logic;
          N_666                     : out   std_logic;
          N_665                     : out   std_logic;
          N_664                     : out   std_logic;
          N_134                     : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          irx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_1
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_1(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    FIFO_8Kx9_0 : FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_1
      port map(RX_FIFO_DIN_pipe(8) => RX_FIFO_DIN_pipe(8), 
        RX_FIFO_DIN_pipe(7) => RX_FIFO_DIN_pipe(7), 
        RX_FIFO_DIN_pipe(6) => RX_FIFO_DIN_pipe(6), 
        RX_FIFO_DIN_pipe(5) => RX_FIFO_DIN_pipe(5), 
        RX_FIFO_DIN_pipe(4) => RX_FIFO_DIN_pipe(4), 
        RX_FIFO_DIN_pipe(3) => RX_FIFO_DIN_pipe(3), 
        RX_FIFO_DIN_pipe(2) => RX_FIFO_DIN_pipe(2), 
        RX_FIFO_DIN_pipe(1) => RX_FIFO_DIN_pipe(1), 
        RX_FIFO_DIN_pipe(0) => RX_FIFO_DIN_pipe(0), 
        ReadFIFO_Write_Ptr(1) => ReadFIFO_Write_Ptr(1), 
        ReadFIFO_Write_Ptr(0) => ReadFIFO_Write_Ptr(0), 
        iRX_FIFO_OVERFLOW_0 => iRX_FIFO_OVERFLOW_0, 
        iRX_FIFO_Full_0 => iRX_FIFO_Full_0, iRX_FIFO_UNDERRUN_0
         => iRX_FIFO_UNDERRUN_0, iRX_FIFO_Empty_0 => 
        iRX_FIFO_Empty_0, RX_FIFO_DOUT_2_0 => RX_FIFO_DOUT_2_0, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, N_1466 => 
        N_1466, N_667 => N_667, N_669 => N_669, N_716 => N_716, 
        N_670 => N_670, N_668 => N_668, N_666 => N_666, N_665 => 
        N_665, N_664 => N_664, N_134 => N_134, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz, 
        irx_fifo_rst_i => irx_fifo_rst_i);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_2 is

    port( fifo_MEMWADDR             : in    std_logic_vector(10 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          fifo_MEMRADDR             : in    std_logic_vector(10 downto 0);
          RDATA_int                 : out   std_logic_vector(8 downto 0);
          fifo_MEMWE                : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          N_1006_i                  : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_2;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_2 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component RAM1K18
    generic (MEMORYFILE:string := "");

    port( A_DOUT        : out   std_logic_vector(17 downto 0);
          B_DOUT        : out   std_logic_vector(17 downto 0);
          BUSY          : out   std_logic;
          A_CLK         : in    std_logic := 'U';
          A_DOUT_CLK    : in    std_logic := 'U';
          A_ARST_N      : in    std_logic := 'U';
          A_DOUT_EN     : in    std_logic := 'U';
          A_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_DOUT_ARST_N : in    std_logic := 'U';
          A_DOUT_SRST_N : in    std_logic := 'U';
          A_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          A_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          A_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          B_CLK         : in    std_logic := 'U';
          B_DOUT_CLK    : in    std_logic := 'U';
          B_ARST_N      : in    std_logic := 'U';
          B_DOUT_EN     : in    std_logic := 'U';
          B_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_DOUT_ARST_N : in    std_logic := 'U';
          B_DOUT_SRST_N : in    std_logic := 'U';
          B_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          B_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          B_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          A_EN          : in    std_logic := 'U';
          A_DOUT_LAT    : in    std_logic := 'U';
          A_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_WMODE       : in    std_logic := 'U';
          B_EN          : in    std_logic := 'U';
          B_DOUT_LAT    : in    std_logic := 'U';
          B_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_WMODE       : in    std_logic := 'U';
          SII_LOCK      : in    std_logic := 'U'
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;
    signal nc24, nc1, nc8, nc13, nc16, nc19, nc25, nc20, nc27, 
        nc9, nc22, nc14, nc5, nc21, nc15, nc3, nc10, nc7, nc17, 
        nc4, nc12, nc2, nc23, nc18, nc26, nc6, nc11 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C0 : RAM1K18
      port map(A_DOUT(17) => nc24, A_DOUT(16) => nc1, A_DOUT(15)
         => nc8, A_DOUT(14) => nc13, A_DOUT(13) => nc16, 
        A_DOUT(12) => nc19, A_DOUT(11) => nc25, A_DOUT(10) => 
        nc20, A_DOUT(9) => nc27, A_DOUT(8) => RDATA_int(8), 
        A_DOUT(7) => RDATA_int(7), A_DOUT(6) => RDATA_int(6), 
        A_DOUT(5) => RDATA_int(5), A_DOUT(4) => RDATA_int(4), 
        A_DOUT(3) => RDATA_int(3), A_DOUT(2) => RDATA_int(2), 
        A_DOUT(1) => RDATA_int(1), A_DOUT(0) => RDATA_int(0), 
        B_DOUT(17) => nc9, B_DOUT(16) => nc22, B_DOUT(15) => nc14, 
        B_DOUT(14) => nc5, B_DOUT(13) => nc21, B_DOUT(12) => nc15, 
        B_DOUT(11) => nc3, B_DOUT(10) => nc10, B_DOUT(9) => nc7, 
        B_DOUT(8) => nc17, B_DOUT(7) => nc4, B_DOUT(6) => nc12, 
        B_DOUT(5) => nc2, B_DOUT(4) => nc23, B_DOUT(3) => nc18, 
        B_DOUT(2) => nc26, B_DOUT(1) => nc6, B_DOUT(0) => nc11, 
        BUSY => OPEN, A_CLK => m2s010_som_sb_0_CCC_71MHz, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => VCC_net_1, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_1006_i, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => GND_net_1, A_DIN(15) => GND_net_1, 
        A_DIN(14) => GND_net_1, A_DIN(13) => GND_net_1, A_DIN(12)
         => GND_net_1, A_DIN(11) => GND_net_1, A_DIN(10) => 
        GND_net_1, A_DIN(9) => GND_net_1, A_DIN(8) => GND_net_1, 
        A_DIN(7) => GND_net_1, A_DIN(6) => GND_net_1, A_DIN(5)
         => GND_net_1, A_DIN(4) => GND_net_1, A_DIN(3) => 
        GND_net_1, A_DIN(2) => GND_net_1, A_DIN(1) => GND_net_1, 
        A_DIN(0) => GND_net_1, A_ADDR(13) => fifo_MEMRADDR(10), 
        A_ADDR(12) => fifo_MEMRADDR(9), A_ADDR(11) => 
        fifo_MEMRADDR(8), A_ADDR(10) => fifo_MEMRADDR(7), 
        A_ADDR(9) => fifo_MEMRADDR(6), A_ADDR(8) => 
        fifo_MEMRADDR(5), A_ADDR(7) => fifo_MEMRADDR(4), 
        A_ADDR(6) => fifo_MEMRADDR(3), A_ADDR(5) => 
        fifo_MEMRADDR(2), A_ADDR(4) => fifo_MEMRADDR(1), 
        A_ADDR(3) => fifo_MEMRADDR(0), A_ADDR(2) => GND_net_1, 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => RX_FIFO_DIN_pipe(8), B_DIN(7) => RX_FIFO_DIN_pipe(7), 
        B_DIN(6) => RX_FIFO_DIN_pipe(6), B_DIN(5) => 
        RX_FIFO_DIN_pipe(5), B_DIN(4) => RX_FIFO_DIN_pipe(4), 
        B_DIN(3) => RX_FIFO_DIN_pipe(3), B_DIN(2) => 
        RX_FIFO_DIN_pipe(2), B_DIN(1) => RX_FIFO_DIN_pipe(1), 
        B_DIN(0) => RX_FIFO_DIN_pipe(0), B_ADDR(13) => 
        fifo_MEMWADDR(10), B_ADDR(12) => fifo_MEMWADDR(9), 
        B_ADDR(11) => fifo_MEMWADDR(8), B_ADDR(10) => 
        fifo_MEMWADDR(7), B_ADDR(9) => fifo_MEMWADDR(6), 
        B_ADDR(8) => fifo_MEMWADDR(5), B_ADDR(7) => 
        fifo_MEMWADDR(4), B_ADDR(6) => fifo_MEMWADDR(3), 
        B_ADDR(5) => fifo_MEMWADDR(2), B_ADDR(4) => 
        fifo_MEMWADDR(1), B_ADDR(3) => fifo_MEMWADDR(0), 
        B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, B_ADDR(0)
         => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0) => 
        VCC_net_1, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_2 is

    port( RDATA_int                 : out   std_logic_vector(8 downto 0);
          fifo_MEMRADDR             : in    std_logic_vector(10 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          fifo_MEMWADDR             : in    std_logic_vector(10 downto 0);
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          N_1006_i                  : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          fifo_MEMWE                : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_2;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_2 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_2
    port( fifo_MEMWADDR             : in    std_logic_vector(10 downto 0) := (others => 'U');
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          fifo_MEMRADDR             : in    std_logic_vector(10 downto 0) := (others => 'U');
          RDATA_int                 : out   std_logic_vector(8 downto 0);
          fifo_MEMWE                : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          N_1006_i                  : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_2
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_2(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    L1_asyncnonpipe : FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_2
      port map(fifo_MEMWADDR(10) => fifo_MEMWADDR(10), 
        fifo_MEMWADDR(9) => fifo_MEMWADDR(9), fifo_MEMWADDR(8)
         => fifo_MEMWADDR(8), fifo_MEMWADDR(7) => 
        fifo_MEMWADDR(7), fifo_MEMWADDR(6) => fifo_MEMWADDR(6), 
        fifo_MEMWADDR(5) => fifo_MEMWADDR(5), fifo_MEMWADDR(4)
         => fifo_MEMWADDR(4), fifo_MEMWADDR(3) => 
        fifo_MEMWADDR(3), fifo_MEMWADDR(2) => fifo_MEMWADDR(2), 
        fifo_MEMWADDR(1) => fifo_MEMWADDR(1), fifo_MEMWADDR(0)
         => fifo_MEMWADDR(0), RX_FIFO_DIN_pipe(8) => 
        RX_FIFO_DIN_pipe(8), RX_FIFO_DIN_pipe(7) => 
        RX_FIFO_DIN_pipe(7), RX_FIFO_DIN_pipe(6) => 
        RX_FIFO_DIN_pipe(6), RX_FIFO_DIN_pipe(5) => 
        RX_FIFO_DIN_pipe(5), RX_FIFO_DIN_pipe(4) => 
        RX_FIFO_DIN_pipe(4), RX_FIFO_DIN_pipe(3) => 
        RX_FIFO_DIN_pipe(3), RX_FIFO_DIN_pipe(2) => 
        RX_FIFO_DIN_pipe(2), RX_FIFO_DIN_pipe(1) => 
        RX_FIFO_DIN_pipe(1), RX_FIFO_DIN_pipe(0) => 
        RX_FIFO_DIN_pipe(0), fifo_MEMRADDR(10) => 
        fifo_MEMRADDR(10), fifo_MEMRADDR(9) => fifo_MEMRADDR(9), 
        fifo_MEMRADDR(8) => fifo_MEMRADDR(8), fifo_MEMRADDR(7)
         => fifo_MEMRADDR(7), fifo_MEMRADDR(6) => 
        fifo_MEMRADDR(6), fifo_MEMRADDR(5) => fifo_MEMRADDR(5), 
        fifo_MEMRADDR(4) => fifo_MEMRADDR(4), fifo_MEMRADDR(3)
         => fifo_MEMRADDR(3), fifo_MEMRADDR(2) => 
        fifo_MEMRADDR(2), fifo_MEMRADDR(1) => fifo_MEMRADDR(1), 
        fifo_MEMRADDR(0) => fifo_MEMRADDR(0), RDATA_int(8) => 
        RDATA_int(8), RDATA_int(7) => RDATA_int(7), RDATA_int(6)
         => RDATA_int(6), RDATA_int(5) => RDATA_int(5), 
        RDATA_int(4) => RDATA_int(4), RDATA_int(3) => 
        RDATA_int(3), RDATA_int(2) => RDATA_int(2), RDATA_int(1)
         => RDATA_int(1), RDATA_int(0) => RDATA_int(0), 
        fifo_MEMWE => fifo_MEMWE, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, N_1006_i => N_1006_i, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_6 is

    port( wptr_bin_sync  : inout std_logic_vector(11 downto 0) := (others => 'Z');
          wptr_gray_sync : in    std_logic_vector(10 downto 0)
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_6;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_6 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    \bin_out_xhdl1_0_a2[1]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(3), B => wptr_gray_sync(1), C
         => wptr_bin_sync(4), D => wptr_gray_sync(2), Y => 
        wptr_bin_sync(1));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \bin_out_xhdl1_0_a2[5]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(7), B => wptr_gray_sync(6), C
         => wptr_gray_sync(5), D => wptr_bin_sync(8), Y => 
        wptr_bin_sync(5));
    
    \bin_out_xhdl1_0_a2[2]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(4), B => wptr_gray_sync(3), C
         => wptr_gray_sync(2), D => wptr_bin_sync(5), Y => 
        wptr_bin_sync(2));
    
    \bin_out_xhdl1_0_a2[0]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(2), B => wptr_bin_sync(3), C
         => wptr_gray_sync(0), D => wptr_gray_sync(1), Y => 
        wptr_bin_sync(0));
    
    \bin_out_xhdl1_i_o2[9]\ : CFG3
      generic map(INIT => x"96")

      port map(A => wptr_gray_sync(10), B => wptr_gray_sync(9), C
         => wptr_bin_sync(11), Y => wptr_bin_sync(9));
    
    \bin_out_xhdl1_i_o2[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => wptr_bin_sync(11), B => wptr_gray_sync(10), Y
         => wptr_bin_sync(10));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \bin_out_xhdl1_0_a2[6]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(8), B => wptr_gray_sync(7), C
         => wptr_gray_sync(6), D => wptr_bin_sync(9), Y => 
        wptr_bin_sync(6));
    
    \bin_out_xhdl1_0_a2[4]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(6), B => wptr_gray_sync(5), C
         => wptr_gray_sync(4), D => wptr_bin_sync(7), Y => 
        wptr_bin_sync(4));
    
    \bin_out_xhdl1_0_a2[8]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(10), B => wptr_gray_sync(9), C
         => wptr_gray_sync(8), D => wptr_bin_sync(11), Y => 
        wptr_bin_sync(8));
    
    \bin_out_xhdl1_0_a2[7]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(9), B => wptr_gray_sync(8), C
         => wptr_gray_sync(7), D => wptr_bin_sync(10), Y => 
        wptr_bin_sync(7));
    
    \bin_out_xhdl1_0_a2[3]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(5), B => wptr_gray_sync(4), C
         => wptr_gray_sync(3), D => wptr_bin_sync(6), Y => 
        wptr_bin_sync(3));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_3 is

    port( wptr_gray                 : in    std_logic_vector(11 downto 0);
          wptr_gray_sync            : out   std_logic_vector(10 downto 0);
          wptr_bin_sync_0           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          irx_fifo_rst_i            : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_3;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_3 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \sync_int[10]_net_1\, VCC_net_1, GND_net_1, 
        \sync_int[11]_net_1\, \sync_int[0]_net_1\, 
        \sync_int[1]_net_1\, \sync_int[2]_net_1\, 
        \sync_int[3]_net_1\, \sync_int[4]_net_1\, 
        \sync_int[5]_net_1\, \sync_int[6]_net_1\, 
        \sync_int[7]_net_1\, \sync_int[8]_net_1\, 
        \sync_int[9]_net_1\ : std_logic;

begin 


    \sync_int[9]\ : SLE
      port map(D => wptr_gray(9), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[9]_net_1\);
    
    \sync_int[4]\ : SLE
      port map(D => wptr_gray(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[4]_net_1\);
    
    \sync_out_xhdl1[10]\ : SLE
      port map(D => \sync_int[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(10));
    
    \sync_int[1]\ : SLE
      port map(D => wptr_gray(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[1]_net_1\);
    
    \sync_int[11]\ : SLE
      port map(D => wptr_gray(11), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[11]_net_1\);
    
    \sync_out_xhdl1[6]\ : SLE
      port map(D => \sync_int[6]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(6));
    
    \sync_out_xhdl1[3]\ : SLE
      port map(D => \sync_int[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(3));
    
    \sync_int[6]\ : SLE
      port map(D => wptr_gray(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[6]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \sync_out_xhdl1[11]\ : SLE
      port map(D => \sync_int[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_bin_sync_0);
    
    \sync_int[3]\ : SLE
      port map(D => wptr_gray(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[3]_net_1\);
    
    \sync_out_xhdl1[4]\ : SLE
      port map(D => \sync_int[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(4));
    
    \sync_int[0]\ : SLE
      port map(D => wptr_gray(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[0]_net_1\);
    
    \sync_out_xhdl1[1]\ : SLE
      port map(D => \sync_int[1]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(1));
    
    \sync_int[5]\ : SLE
      port map(D => wptr_gray(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[5]_net_1\);
    
    \sync_int[2]\ : SLE
      port map(D => wptr_gray(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[2]_net_1\);
    
    \sync_out_xhdl1[9]\ : SLE
      port map(D => \sync_int[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(9));
    
    \sync_out_xhdl1[2]\ : SLE
      port map(D => \sync_int[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(2));
    
    \sync_int[8]\ : SLE
      port map(D => wptr_gray(8), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[8]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sync_out_xhdl1[7]\ : SLE
      port map(D => \sync_int[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(7));
    
    \sync_out_xhdl1[5]\ : SLE
      port map(D => \sync_int[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(5));
    
    \sync_out_xhdl1[0]\ : SLE
      port map(D => \sync_int[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(0));
    
    \sync_out_xhdl1[8]\ : SLE
      port map(D => \sync_int[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(8));
    
    \sync_int[7]\ : SLE
      port map(D => wptr_gray(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[7]_net_1\);
    
    \sync_int[10]\ : SLE
      port map(D => wptr_gray(10), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_2 is

    port( rptr_gray           : in    std_logic_vector(11 downto 0);
          rptr_gray_sync      : out   std_logic_vector(10 downto 0);
          rptr_bin_sync_0     : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          irx_fifo_rst_i      : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_2;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_2 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \sync_int[4]_net_1\, GND_net_1, 
        \sync_int[5]_net_1\, \sync_int[6]_net_1\, 
        \sync_int[7]_net_1\, \sync_int[8]_net_1\, 
        \sync_int[9]_net_1\, \sync_int[10]_net_1\, 
        \sync_int[11]_net_1\, \sync_int[1]_net_1\, 
        \sync_int[2]_net_1\, \sync_int[3]_net_1\, 
        \sync_int[0]_net_1\ : std_logic;

begin 


    \sync_int[9]\ : SLE
      port map(D => rptr_gray(9), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[9]_net_1\);
    
    \sync_int[4]\ : SLE
      port map(D => rptr_gray(4), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[4]_net_1\);
    
    \sync_out_xhdl1[10]\ : SLE
      port map(D => \sync_int[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(10));
    
    \sync_int[1]\ : SLE
      port map(D => rptr_gray(1), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[1]_net_1\);
    
    \sync_int[11]\ : SLE
      port map(D => rptr_gray(11), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[11]_net_1\);
    
    \sync_out_xhdl1[6]\ : SLE
      port map(D => \sync_int[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(6));
    
    \sync_out_xhdl1[3]\ : SLE
      port map(D => \sync_int[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(3));
    
    \sync_int[6]\ : SLE
      port map(D => rptr_gray(6), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[6]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \sync_out_xhdl1[11]\ : SLE
      port map(D => \sync_int[11]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_bin_sync_0);
    
    \sync_int[3]\ : SLE
      port map(D => rptr_gray(3), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[3]_net_1\);
    
    \sync_out_xhdl1[4]\ : SLE
      port map(D => \sync_int[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(4));
    
    \sync_int[0]\ : SLE
      port map(D => rptr_gray(0), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[0]_net_1\);
    
    \sync_out_xhdl1[1]\ : SLE
      port map(D => \sync_int[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(1));
    
    \sync_int[5]\ : SLE
      port map(D => rptr_gray(5), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[5]_net_1\);
    
    \sync_int[2]\ : SLE
      port map(D => rptr_gray(2), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[2]_net_1\);
    
    \sync_out_xhdl1[9]\ : SLE
      port map(D => \sync_int[9]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(9));
    
    \sync_out_xhdl1[2]\ : SLE
      port map(D => \sync_int[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(2));
    
    \sync_int[8]\ : SLE
      port map(D => rptr_gray(8), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[8]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sync_out_xhdl1[7]\ : SLE
      port map(D => \sync_int[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(7));
    
    \sync_out_xhdl1[5]\ : SLE
      port map(D => \sync_int[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(5));
    
    \sync_out_xhdl1[0]\ : SLE
      port map(D => \sync_int[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(0));
    
    \sync_out_xhdl1[8]\ : SLE
      port map(D => \sync_int[8]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(8));
    
    \sync_int[7]\ : SLE
      port map(D => rptr_gray(7), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[7]_net_1\);
    
    \sync_int[10]\ : SLE
      port map(D => rptr_gray(10), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_5 is

    port( rptr_bin_sync  : inout std_logic_vector(11 downto 0) := (others => 'Z');
          rptr_gray_sync : in    std_logic_vector(10 downto 0)
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_5;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_5 is 

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    \bin_out_xhdl1_0_a2[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(2), B => rptr_gray_sync(1), Y
         => rptr_bin_sync(1));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \bin_out_xhdl1_0_a2[5]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(6), B => rptr_bin_sync(7), C
         => rptr_gray_sync(5), Y => rptr_bin_sync(5));
    
    \bin_out_xhdl1_0_a2[2]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(2), B => rptr_gray_sync(3), C
         => rptr_gray_sync(4), D => rptr_bin_sync(5), Y => 
        rptr_bin_sync(2));
    
    \bin_out_xhdl1_0_a2[0]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(1), B => rptr_bin_sync(2), C
         => rptr_gray_sync(0), Y => rptr_bin_sync(0));
    
    \bin_out_xhdl1_i_o2[9]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(9), B => rptr_gray_sync(10), C
         => rptr_bin_sync(11), Y => rptr_bin_sync(9));
    
    \bin_out_xhdl1_i_o2[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(11), B => rptr_gray_sync(10), Y
         => rptr_bin_sync(10));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \bin_out_xhdl1_0_a2[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(7), B => rptr_gray_sync(6), Y
         => rptr_bin_sync(6));
    
    \bin_out_xhdl1_0_a2[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(5), B => rptr_gray_sync(4), Y
         => rptr_bin_sync(4));
    
    \bin_out_xhdl1_0_a2[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(9), B => rptr_gray_sync(8), Y
         => rptr_bin_sync(8));
    
    \bin_out_xhdl1_0_a2[7]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(8), B => rptr_bin_sync(9), C
         => rptr_gray_sync(7), Y => rptr_bin_sync(7));
    
    \bin_out_xhdl1_0_a2[3]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(4), B => rptr_bin_sync(5), C
         => rptr_gray_sync(3), Y => rptr_bin_sync(3));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_2 is

    port( ReadFIFO_Write_Ptr        : in    std_logic_vector(1 downto 0);
          fifo_MEMWADDR             : out   std_logic_vector(10 downto 0);
          fifo_MEMRADDR             : out   std_logic_vector(10 downto 0);
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          N_154_i_i                 : out   std_logic;
          N_89_i                    : out   std_logic;
          REN_d1                    : in    std_logic;
          N_133                     : in    std_logic;
          N_1466                    : in    std_logic;
          N_1006_i                  : out   std_logic;
          fifo_MEMWE                : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          irx_fifo_rst_i            : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_2;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_2 is 

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_6
    port( wptr_bin_sync  : inout   std_logic_vector(11 downto 0);
          wptr_gray_sync : in    std_logic_vector(10 downto 0) := (others => 'U')
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_3
    port( wptr_gray                 : in    std_logic_vector(11 downto 0) := (others => 'U');
          wptr_gray_sync            : out   std_logic_vector(10 downto 0);
          wptr_bin_sync_0           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          irx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_2
    port( rptr_gray           : in    std_logic_vector(11 downto 0) := (others => 'U');
          rptr_gray_sync      : out   std_logic_vector(10 downto 0);
          rptr_bin_sync_0     : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          irx_fifo_rst_i      : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_5
    port( rptr_bin_sync  : inout   std_logic_vector(11 downto 0);
          rptr_gray_sync : in    std_logic_vector(10 downto 0) := (others => 'U')
        );
  end component;

    signal \rptr[0]_net_1\, \rptr_s[0]\, \fifo_MEMRADDR[0]\, 
        \memraddr_r_s[0]\, \wptr[0]_net_1\, \wptr_s[0]\, 
        \wptr_gray[10]_net_1\, VCC_net_1, \wptr_gray_1[10]_net_1\, 
        GND_net_1, \wptr_gray[11]_net_1\, \wptr[11]_net_1\, 
        \rptr_gray[0]_net_1\, \rptr_gray_1[0]_net_1\, 
        \rptr_gray[1]_net_1\, \rptr_gray_1[1]_net_1\, 
        \rptr_gray[2]_net_1\, \rptr_gray_1[2]_net_1\, 
        \rptr_gray[3]_net_1\, \rptr_gray_1[3]_net_1\, 
        \rptr_gray[4]_net_1\, \rptr_gray_1[4]_net_1\, 
        \rptr_gray[5]_net_1\, \rptr_gray_1[5]_net_1\, 
        \rptr_gray[6]_net_1\, \rptr_gray_1[6]_net_1\, 
        \rptr_gray[7]_net_1\, \rptr_gray_1[7]_net_1\, 
        \rptr_gray[8]_net_1\, \rptr_gray_1[8]_net_1\, 
        \rptr_gray[9]_net_1\, \rptr_gray_1[9]_net_1\, 
        \rptr_gray[10]_net_1\, \rptr_gray_1[10]_net_1\, 
        \rptr_gray[11]_net_1\, \rptr[11]_net_1\, 
        \wptr_bin_sync2[7]_net_1\, \wptr_bin_sync[7]\, 
        \wptr_bin_sync2[8]_net_1\, \wptr_bin_sync[8]\, 
        \wptr_bin_sync2[9]_net_1\, \wptr_bin_sync[9]\, 
        \wptr_bin_sync2[10]_net_1\, \wptr_bin_sync[10]\, 
        \wptr_bin_sync2[11]_net_1\, \wptr_bin_sync[11]\, 
        \wptr_gray[0]_net_1\, \wptr_gray_1[0]_net_1\, 
        \wptr_gray[1]_net_1\, \wptr_gray_1[1]_net_1\, 
        \wptr_gray[2]_net_1\, \wptr_gray_1[2]_net_1\, 
        \wptr_gray[3]_net_1\, \wptr_gray_1[3]_net_1\, 
        \wptr_gray[4]_net_1\, \wptr_gray_1[4]_net_1\, 
        \wptr_gray[5]_net_1\, \wptr_gray_1[5]_net_1\, 
        \wptr_gray[6]_net_1\, \wptr_gray_1[6]_net_1\, 
        \wptr_gray[7]_net_1\, \wptr_gray_1[7]_net_1\, 
        \wptr_gray[8]_net_1\, \wptr_gray_1[8]_net_1\, 
        \wptr_gray[9]_net_1\, \wptr_gray_1[9]_net_1\, rdiff_bus, 
        \wptr_bin_sync[0]\, \wptr_bin_sync2[1]_net_1\, 
        \wptr_bin_sync[1]\, \wptr_bin_sync2[2]_net_1\, 
        \wptr_bin_sync[2]\, \wptr_bin_sync2[3]_net_1\, 
        \wptr_bin_sync[3]\, \wptr_bin_sync2[4]_net_1\, 
        \wptr_bin_sync[4]\, \wptr_bin_sync2[5]_net_1\, 
        \wptr_bin_sync[5]\, \wptr_bin_sync2[6]_net_1\, 
        \wptr_bin_sync[6]\, \rptr_bin_sync2[7]_net_1\, 
        \rptr_bin_sync[7]\, \rptr_bin_sync2[8]_net_1\, 
        \rptr_bin_sync[8]\, \rptr_bin_sync2[9]_net_1\, 
        \rptr_bin_sync[9]\, \rptr_bin_sync2[10]_net_1\, 
        \rptr_bin_sync[10]\, \rptr_bin_sync2[11]_net_1\, 
        \rptr_bin_sync[11]\, un1_we_p, \rptr_bin_sync2[0]_net_1\, 
        \rptr_bin_sync[0]\, \rptr_bin_sync2[1]_net_1\, 
        \rptr_bin_sync[1]\, \rptr_bin_sync2[2]_net_1\, 
        \rptr_bin_sync[2]\, \rptr_bin_sync2[3]_net_1\, 
        \rptr_bin_sync[3]\, \rptr_bin_sync2[4]_net_1\, 
        \rptr_bin_sync[4]\, \rptr_bin_sync2[5]_net_1\, 
        \rptr_bin_sync[5]\, \rptr_bin_sync2[6]_net_1\, 
        \rptr_bin_sync[6]\, \iRX_FIFO_Full_0\, fulli, 
        un2_re_p_i_i_a3_2, \iRX_FIFO_Empty_0\, empty_r_3, 
        \fifo_MEMWE\, \wptr[1]_net_1\, \wptr_s[1]\, 
        \wptr[2]_net_1\, \wptr_s[2]\, \wptr[3]_net_1\, 
        \wptr_s[3]\, \wptr[4]_net_1\, \wptr_s[4]\, 
        \wptr[5]_net_1\, \wptr_s[5]\, \wptr[6]_net_1\, 
        \wptr_s[6]\, \wptr[7]_net_1\, \wptr_s[7]\, 
        \wptr[8]_net_1\, \wptr_s[8]\, \wptr[9]_net_1\, 
        \wptr_s[9]\, \wptr[10]_net_1\, \wptr_s[10]\, 
        \wptr_s[11]_net_1\, \N_1006_i\, \fifo_MEMRADDR[1]\, 
        \memraddr_r_s[1]\, \fifo_MEMRADDR[2]\, \memraddr_r_s[2]\, 
        \fifo_MEMRADDR[3]\, \memraddr_r_s[3]\, \fifo_MEMRADDR[4]\, 
        \memraddr_r_s[4]\, \fifo_MEMRADDR[5]\, \memraddr_r_s[5]\, 
        \fifo_MEMRADDR[6]\, \memraddr_r_s[6]\, \fifo_MEMRADDR[7]\, 
        \memraddr_r_s[7]\, \fifo_MEMRADDR[8]\, \memraddr_r_s[8]\, 
        \fifo_MEMRADDR[9]\, \memraddr_r_s[9]\, 
        \fifo_MEMRADDR[10]\, \memraddr_r_s[10]_net_1\, 
        \fifo_MEMWADDR[0]\, \memwaddr_r_s[0]\, N_249, 
        \fifo_MEMWADDR[1]\, \memwaddr_r_s[1]\, \fifo_MEMWADDR[2]\, 
        \memwaddr_r_s[2]\, \fifo_MEMWADDR[3]\, \memwaddr_r_s[3]\, 
        \fifo_MEMWADDR[4]\, \memwaddr_r_s[4]\, \fifo_MEMWADDR[5]\, 
        \memwaddr_r_s[5]\, \fifo_MEMWADDR[6]\, \memwaddr_r_s[6]\, 
        \fifo_MEMWADDR[7]\, \memwaddr_r_s[7]\, \fifo_MEMWADDR[8]\, 
        \memwaddr_r_s[8]\, \fifo_MEMWADDR[9]\, \memwaddr_r_s[9]\, 
        \fifo_MEMWADDR[10]\, \memwaddr_r_s[10]_net_1\, 
        \rptr[1]_net_1\, \rptr_s[1]\, \rptr[2]_net_1\, 
        \rptr_s[2]\, \rptr[3]_net_1\, \rptr_s[3]\, 
        \rptr[4]_net_1\, \rptr_s[4]\, \rptr[5]_net_1\, 
        \rptr_s[5]\, \rptr[6]_net_1\, \rptr_s[6]\, 
        \rptr[7]_net_1\, \rptr_s[7]\, \rptr[8]_net_1\, 
        \rptr_s[8]\, \rptr[9]_net_1\, \rptr_s[9]\, 
        \rptr[10]_net_1\, \rptr_s[10]\, \rptr_s[11]_net_1\, 
        memwaddr_r_cry_cy, \memwaddr_r_cry[0]_net_1\, 
        \memwaddr_r_cry[1]_net_1\, \memwaddr_r_cry[2]_net_1\, 
        \memwaddr_r_cry[3]_net_1\, \memwaddr_r_cry[4]_net_1\, 
        \memwaddr_r_cry[5]_net_1\, \memwaddr_r_cry[6]_net_1\, 
        \memwaddr_r_cry[7]_net_1\, \memwaddr_r_cry[8]_net_1\, 
        \memwaddr_r_cry[9]_net_1\, \rdiff_bus_cry_0\, 
        rdiff_bus_cry_0_Y_3, \rdiff_bus_cry_1\, \rdiff_bus[1]\, 
        \rdiff_bus_cry_2\, \rdiff_bus[2]\, \rdiff_bus_cry_3\, 
        \rdiff_bus[3]\, \rdiff_bus_cry_4\, \rdiff_bus[4]\, 
        \rdiff_bus_cry_5\, \rdiff_bus[5]\, \rdiff_bus_cry_6\, 
        \rdiff_bus[6]\, \rdiff_bus_cry_7\, \rdiff_bus[7]\, 
        \rdiff_bus_cry_8\, \rdiff_bus[8]\, \rdiff_bus_cry_9\, 
        \rdiff_bus[9]\, \rdiff_bus[11]\, \rdiff_bus_cry_10\, 
        \rdiff_bus[10]\, \wdiff_bus_cry_0\, wdiff_bus_cry_0_Y_3, 
        \wdiff_bus_cry_1\, \wdiff_bus[1]\, \wdiff_bus_cry_2\, 
        \wdiff_bus[2]\, \wdiff_bus_cry_3\, \wdiff_bus[3]\, 
        \wdiff_bus_cry_4\, \wdiff_bus[4]\, \wdiff_bus_cry_5\, 
        \wdiff_bus[5]\, \wdiff_bus_cry_6\, \wdiff_bus[6]\, 
        \wdiff_bus_cry_7\, \wdiff_bus[7]\, \wdiff_bus_cry_8\, 
        \wdiff_bus[8]\, \wdiff_bus_cry_9\, \wdiff_bus[9]\, 
        \wdiff_bus[11]\, \wdiff_bus_cry_10\, \wdiff_bus[10]\, 
        rptr_s_374_FCO, \rptr_cry[1]_net_1\, \rptr_cry[2]_net_1\, 
        \rptr_cry[3]_net_1\, \rptr_cry[4]_net_1\, 
        \rptr_cry[5]_net_1\, \rptr_cry[6]_net_1\, 
        \rptr_cry[7]_net_1\, \rptr_cry[8]_net_1\, 
        \rptr_cry[9]_net_1\, \rptr_cry[10]_net_1\, 
        memraddr_r_s_375_FCO, \memraddr_r_cry[1]_net_1\, 
        \memraddr_r_cry[2]_net_1\, \memraddr_r_cry[3]_net_1\, 
        \memraddr_r_cry[4]_net_1\, \memraddr_r_cry[5]_net_1\, 
        \memraddr_r_cry[6]_net_1\, \memraddr_r_cry[7]_net_1\, 
        \memraddr_r_cry[8]_net_1\, \memraddr_r_cry[9]_net_1\, 
        wptr_s_376_FCO, \wptr_cry[1]_net_1\, \wptr_cry[2]_net_1\, 
        \wptr_cry[3]_net_1\, \wptr_cry[4]_net_1\, 
        \wptr_cry[5]_net_1\, \wptr_cry[6]_net_1\, 
        \wptr_cry[7]_net_1\, \wptr_cry[8]_net_1\, 
        \wptr_cry[9]_net_1\, \wptr_cry[10]_net_1\, 
        empty_r_3_0_a2_1, \fulli_0_a2_7\, \fulli_0_a2_6\, 
        empty_r_3_0_a2_7, empty_r_3_0_a2_9, \fulli_0_a2_8\, 
        empty_r_3_0_a2_5, \wptr_gray_sync[0]\, 
        \wptr_gray_sync[1]\, \wptr_gray_sync[2]\, 
        \wptr_gray_sync[3]\, \wptr_gray_sync[4]\, 
        \wptr_gray_sync[5]\, \wptr_gray_sync[6]\, 
        \wptr_gray_sync[7]\, \wptr_gray_sync[8]\, 
        \wptr_gray_sync[9]\, \wptr_gray_sync[10]\, 
        \rptr_gray_sync[0]\, \rptr_gray_sync[1]\, 
        \rptr_gray_sync[2]\, \rptr_gray_sync[3]\, 
        \rptr_gray_sync[4]\, \rptr_gray_sync[5]\, 
        \rptr_gray_sync[6]\, \rptr_gray_sync[7]\, 
        \rptr_gray_sync[8]\, \rptr_gray_sync[9]\, 
        \rptr_gray_sync[10]\ : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_6
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_6(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_3
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_3(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_2
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_2(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_5
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_5(DEF_ARCH);
begin 

    fifo_MEMWADDR(10) <= \fifo_MEMWADDR[10]\;
    fifo_MEMWADDR(9) <= \fifo_MEMWADDR[9]\;
    fifo_MEMWADDR(8) <= \fifo_MEMWADDR[8]\;
    fifo_MEMWADDR(7) <= \fifo_MEMWADDR[7]\;
    fifo_MEMWADDR(6) <= \fifo_MEMWADDR[6]\;
    fifo_MEMWADDR(5) <= \fifo_MEMWADDR[5]\;
    fifo_MEMWADDR(4) <= \fifo_MEMWADDR[4]\;
    fifo_MEMWADDR(3) <= \fifo_MEMWADDR[3]\;
    fifo_MEMWADDR(2) <= \fifo_MEMWADDR[2]\;
    fifo_MEMWADDR(1) <= \fifo_MEMWADDR[1]\;
    fifo_MEMWADDR(0) <= \fifo_MEMWADDR[0]\;
    fifo_MEMRADDR(10) <= \fifo_MEMRADDR[10]\;
    fifo_MEMRADDR(9) <= \fifo_MEMRADDR[9]\;
    fifo_MEMRADDR(8) <= \fifo_MEMRADDR[8]\;
    fifo_MEMRADDR(7) <= \fifo_MEMRADDR[7]\;
    fifo_MEMRADDR(6) <= \fifo_MEMRADDR[6]\;
    fifo_MEMRADDR(5) <= \fifo_MEMRADDR[5]\;
    fifo_MEMRADDR(4) <= \fifo_MEMRADDR[4]\;
    fifo_MEMRADDR(3) <= \fifo_MEMRADDR[3]\;
    fifo_MEMRADDR(2) <= \fifo_MEMRADDR[2]\;
    fifo_MEMRADDR(1) <= \fifo_MEMRADDR[1]\;
    fifo_MEMRADDR(0) <= \fifo_MEMRADDR[0]\;
    iRX_FIFO_Empty_0 <= \iRX_FIFO_Empty_0\;
    iRX_FIFO_Full_0 <= \iRX_FIFO_Full_0\;
    N_1006_i <= \N_1006_i\;
    fifo_MEMWE <= \fifo_MEMWE\;

    \rptr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[4]_net_1\, S
         => \rptr_s[5]\, Y => OPEN, FCO => \rptr_cry[5]_net_1\);
    
    wdiff_bus_cry_8 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[8]_net_1\, B => 
        \rptr_bin_sync2[8]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_7\, S => \wdiff_bus[8]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_8\);
    
    \wptr_gray[4]\ : SLE
      port map(D => \wptr_gray_1[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[4]_net_1\);
    
    \rptr_gray_1[3]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[3]_net_1\, B => \rptr[4]_net_1\, Y => 
        \rptr_gray_1[3]_net_1\);
    
    \rptr_bin_sync2[6]\ : SLE
      port map(D => \rptr_bin_sync[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[6]_net_1\);
    
    fulli_0_a2_0_0_a2 : CFG3
      generic map(INIT => x"80")

      port map(A => ReadFIFO_Write_Ptr(0), B => N_1466, C => 
        ReadFIFO_Write_Ptr(1), Y => N_249);
    
    empty_r_RNI4GH71_0 : CFG3
      generic map(INIT => x"A2")

      port map(A => REN_d1, B => N_133, C => \iRX_FIFO_Empty_0\, 
        Y => N_89_i);
    
    \rptr[1]\ : SLE
      port map(D => \rptr_s[1]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1006_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[1]_net_1\);
    
    \wptr_gray_1[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[9]_net_1\, B => \wptr[10]_net_1\, Y => 
        \wptr_gray_1[9]_net_1\);
    
    \rptr_gray_1[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[5]_net_1\, B => \rptr[6]_net_1\, Y => 
        \rptr_gray_1[5]_net_1\);
    
    \rptr_gray[9]\ : SLE
      port map(D => \rptr_gray_1[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[9]_net_1\);
    
    \rptr_gray[8]\ : SLE
      port map(D => \rptr_gray_1[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[8]_net_1\);
    
    \rptr_gray_1[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[2]_net_1\, B => \rptr[3]_net_1\, Y => 
        \rptr_gray_1[2]_net_1\);
    
    \rptr_bin_sync2[7]\ : SLE
      port map(D => \rptr_bin_sync[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[7]_net_1\);
    
    \memwaddr_r[1]\ : SLE
      port map(D => \memwaddr_r_s[1]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_249, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[1]\);
    
    \memwaddr_r_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[5]_net_1\, S => \memwaddr_r_s[6]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[6]_net_1\);
    
    \memwaddr_r_s[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[9]_net_1\, S => \memwaddr_r_s[10]_net_1\, 
        Y => OPEN, FCO => OPEN);
    
    \wptr_gray_1[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[7]_net_1\, B => \wptr[8]_net_1\, Y => 
        \wptr_gray_1[7]_net_1\);
    
    \memraddr_r[0]\ : SLE
      port map(D => \memraddr_r_s[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1006_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[0]\);
    
    \wptr[0]\ : SLE
      port map(D => \wptr_s[0]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[0]_net_1\);
    
    \rptr_bin_sync2[8]\ : SLE
      port map(D => \rptr_bin_sync[8]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[8]_net_1\);
    
    \rptr_gray_1[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[1]_net_1\, B => \rptr[2]_net_1\, Y => 
        \rptr_gray_1[1]_net_1\);
    
    \rptr_gray[10]\ : SLE
      port map(D => \rptr_gray_1[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[10]_net_1\);
    
    \wptr_gray_1[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[0]_net_1\, B => \wptr[1]_net_1\, Y => 
        \wptr_gray_1[0]_net_1\);
    
    wdiff_bus_cry_9 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[9]_net_1\, B => 
        \rptr_bin_sync2[9]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_8\, S => \wdiff_bus[9]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_9\);
    
    \rptr[5]\ : SLE
      port map(D => \rptr_s[5]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1006_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[5]_net_1\);
    
    \rptr_gray[3]\ : SLE
      port map(D => \rptr_gray_1[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[3]_net_1\);
    
    \rptr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[5]_net_1\, S
         => \rptr_s[6]\, Y => OPEN, FCO => \rptr_cry[6]_net_1\);
    
    \memwaddr_r_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[1]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[0]_net_1\, S => \memwaddr_r_s[1]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[1]_net_1\);
    
    fulli_0_a2_6 : CFG4
      generic map(INIT => x"8000")

      port map(A => \wdiff_bus[2]\, B => \wdiff_bus[3]\, C => 
        \wdiff_bus[5]\, D => \wdiff_bus[4]\, Y => \fulli_0_a2_6\);
    
    \wptr_gray[3]\ : SLE
      port map(D => \wptr_gray_1[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[3]_net_1\);
    
    \rptr_gray_1[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[11]_net_1\, B => \rptr[10]_net_1\, Y
         => \rptr_gray_1[10]_net_1\);
    
    wdiff_bus_s_11 : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \rptr_bin_sync2[11]_net_1\, C
         => \wptr[11]_net_1\, D => GND_net_1, FCI => 
        \wdiff_bus_cry_10\, S => \wdiff_bus[11]\, Y => OPEN, FCO
         => OPEN);
    
    \rptr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[7]_net_1\, S
         => \rptr_s[8]\, Y => OPEN, FCO => \rptr_cry[8]_net_1\);
    
    \rptr[7]\ : SLE
      port map(D => \rptr_s[7]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1006_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[7]_net_1\);
    
    rdiff_bus_cry_4 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[4]_net_1\, B => 
        \rptr[4]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_3\, S => \rdiff_bus[4]\, Y => OPEN, FCO
         => \rdiff_bus_cry_4\);
    
    \rptr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[9]_net_1\, S
         => \rptr_s[10]\, Y => OPEN, FCO => \rptr_cry[10]_net_1\);
    
    \rptr_bin_sync2[0]\ : SLE
      port map(D => \rptr_bin_sync[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[0]_net_1\);
    
    \L1.empty_r_3_0_a2_7\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \rdiff_bus[5]\, B => \rdiff_bus[6]\, C => 
        \rdiff_bus[7]\, D => \rdiff_bus[8]\, Y => 
        empty_r_3_0_a2_7);
    
    \wptr[11]\ : SLE
      port map(D => \wptr_s[11]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \wptr[11]_net_1\);
    
    rdiff_bus_cry_1 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[1]_net_1\, B => 
        \rptr[1]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_0\, S => \rdiff_bus[1]\, Y => OPEN, FCO
         => \rdiff_bus_cry_1\);
    
    \memraddr_r[1]\ : SLE
      port map(D => \memraddr_r_s[1]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1006_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[1]\);
    
    \L1.empty_r_3_0_a2_9\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \rdiff_bus[1]\, B => \rdiff_bus[2]\, C => 
        empty_r_3_0_a2_7, D => empty_r_3_0_a2_1, Y => 
        empty_r_3_0_a2_9);
    
    \rptr_bin_sync2[2]\ : SLE
      port map(D => \rptr_bin_sync[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[2]_net_1\);
    
    rdiff_bus_cry_6 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[6]_net_1\, B => 
        \rptr[6]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_5\, S => \rdiff_bus[6]\, Y => OPEN, FCO
         => \rdiff_bus_cry_6\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \memwaddr_r_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[3]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[2]_net_1\, S => \memwaddr_r_s[3]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[3]_net_1\);
    
    \rptr_gray[1]\ : SLE
      port map(D => \rptr_gray_1[1]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[1]_net_1\);
    
    \memwaddr_r[7]\ : SLE
      port map(D => \memwaddr_r_s[7]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_249, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[7]\);
    
    \memraddr_r_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[2]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[1]_net_1\, S => \memraddr_r_s[2]\, Y => 
        OPEN, FCO => \memraddr_r_cry[2]_net_1\);
    
    \wptr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[3]_net_1\, S
         => \wptr_s[4]\, Y => OPEN, FCO => \wptr_cry[4]_net_1\);
    
    \memraddr_r_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[8]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[7]_net_1\, S => \memraddr_r_s[8]\, Y => 
        OPEN, FCO => \memraddr_r_cry[8]_net_1\);
    
    \wptr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[9]_net_1\, S
         => \wptr_s[10]\, Y => OPEN, FCO => \wptr_cry[10]_net_1\);
    
    wdiff_bus_cry_5 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[5]_net_1\, B => 
        \rptr_bin_sync2[5]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_4\, S => \wdiff_bus[5]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_5\);
    
    \memwaddr_r[4]\ : SLE
      port map(D => \memwaddr_r_s[4]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_249, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[4]\);
    
    \wptr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[1]_net_1\, S
         => \wptr_s[2]\, Y => OPEN, FCO => \wptr_cry[2]_net_1\);
    
    wdiff_bus_cry_0 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[0]_net_1\, B => 
        \rptr_bin_sync2[0]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => VCC_net_1, S => OPEN, Y => wdiff_bus_cry_0_Y_3, 
        FCO => \wdiff_bus_cry_0\);
    
    \wptr[1]\ : SLE
      port map(D => \wptr_s[1]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[1]_net_1\);
    
    \rptr_bin_sync2[4]\ : SLE
      port map(D => \rptr_bin_sync[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[4]_net_1\);
    
    \wptr_bin_sync2[6]\ : SLE
      port map(D => \wptr_bin_sync[6]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[6]_net_1\);
    
    \memwaddr_r_cry_cy[0]\ : ARI1
      generic map(INIT => x"45500")

      port map(A => VCC_net_1, B => \iRX_FIFO_Full_0\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => memwaddr_r_cry_cy);
    
    \rptr[3]\ : SLE
      port map(D => \rptr_s[3]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1006_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[3]_net_1\);
    
    \wptr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[2]_net_1\, S
         => \wptr_s[3]\, Y => OPEN, FCO => \wptr_cry[3]_net_1\);
    
    \memwaddr_r_cry[0]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[0]\, C => 
        GND_net_1, D => GND_net_1, FCI => memwaddr_r_cry_cy, S
         => \memwaddr_r_s[0]\, Y => OPEN, FCO => 
        \memwaddr_r_cry[0]_net_1\);
    
    \rptr[6]\ : SLE
      port map(D => \rptr_s[6]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1006_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[6]_net_1\);
    
    rdiff_bus_cry_8 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[8]_net_1\, B => 
        \rptr[8]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_7\, S => \rdiff_bus[8]\, Y => OPEN, FCO
         => \rdiff_bus_cry_8\);
    
    \wptr_gray[10]\ : SLE
      port map(D => \wptr_gray_1[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[10]_net_1\);
    
    rdiff_bus_cry_7 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[7]_net_1\, B => 
        \rptr[7]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_6\, S => \rdiff_bus[7]\, Y => OPEN, FCO
         => \rdiff_bus_cry_7\);
    
    \wptr_bin_sync2[7]\ : SLE
      port map(D => \wptr_bin_sync[7]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[7]_net_1\);
    
    \rptr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[8]_net_1\, S
         => \rptr_s[9]\, Y => OPEN, FCO => \rptr_cry[9]_net_1\);
    
    \rptr_gray[5]\ : SLE
      port map(D => \rptr_gray_1[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[5]_net_1\);
    
    \wptr_gray_1[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[2]_net_1\, B => \wptr[3]_net_1\, Y => 
        \wptr_gray_1[2]_net_1\);
    
    \wptr[5]\ : SLE
      port map(D => \wptr_s[5]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[5]_net_1\);
    
    rdiff_bus_cry_5 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[5]_net_1\, B => 
        \rptr[5]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_4\, S => \rdiff_bus[5]\, Y => OPEN, FCO
         => \rdiff_bus_cry_5\);
    
    \wptr_bin_sync2[8]\ : SLE
      port map(D => \wptr_bin_sync[8]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[8]_net_1\);
    
    \wptr[7]\ : SLE
      port map(D => \wptr_s[7]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[7]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \wptr_gray[1]\ : SLE
      port map(D => \wptr_gray_1[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[1]_net_1\);
    
    \rptr_gray_1[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[9]_net_1\, B => \rptr[10]_net_1\, Y => 
        \rptr_gray_1[9]_net_1\);
    
    \rptr_bin_sync2[5]\ : SLE
      port map(D => \rptr_bin_sync[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[5]_net_1\);
    
    \rptr_bin_sync2[1]\ : SLE
      port map(D => \rptr_bin_sync[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[1]_net_1\);
    
    \memwaddr_r[10]\ : SLE
      port map(D => \memwaddr_r_s[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_249, ALn => irx_fifo_rst_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \fifo_MEMWADDR[10]\);
    
    wdiff_bus_cry_7 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[7]_net_1\, B => 
        \rptr_bin_sync2[7]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_6\, S => \wdiff_bus[7]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_7\);
    
    \wptr_bin_sync2[0]\ : SLE
      port map(D => \wptr_bin_sync[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rdiff_bus);
    
    \L1.un2_re_p_i_i_a3\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_133, B => \iRX_FIFO_Empty_0\, Y => 
        un2_re_p_i_i_a3_2);
    
    \L1.empty_r_3_0_a2_1\ : CFG2
      generic map(INIT => x"1")

      port map(A => \rdiff_bus[4]\, B => \rdiff_bus[3]\, Y => 
        empty_r_3_0_a2_1);
    
    \L1.un1_we_p_0_a2_0_a2\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_249, B => \iRX_FIFO_Full_0\, Y => un1_we_p);
    
    rdiff_bus_s_11 : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \rptr[11]_net_1\, C => 
        \wptr_bin_sync2[11]_net_1\, D => GND_net_1, FCI => 
        \rdiff_bus_cry_10\, S => \rdiff_bus[11]\, Y => OPEN, FCO
         => OPEN);
    
    \memwaddr_r_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[8]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[7]_net_1\, S => \memwaddr_r_s[8]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[8]_net_1\);
    
    \wptr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => wptr_s_376_FCO, S => 
        \wptr_s[1]\, Y => OPEN, FCO => \wptr_cry[1]_net_1\);
    
    \memraddr_r[8]\ : SLE
      port map(D => \memraddr_r_s[8]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1006_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[8]\);
    
    \rptr[9]\ : SLE
      port map(D => \rptr_s[9]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1006_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[9]_net_1\);
    
    \wptr_gray_1[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[6]_net_1\, B => \wptr[7]_net_1\, Y => 
        \wptr_gray_1[6]_net_1\);
    
    \wptr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[6]_net_1\, S
         => \wptr_s[7]\, Y => OPEN, FCO => \wptr_cry[7]_net_1\);
    
    \wptr_bin_sync2[2]\ : SLE
      port map(D => \wptr_bin_sync[2]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[2]_net_1\);
    
    \rptr_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \rptr[0]_net_1\, Y => \rptr_s[0]\);
    
    \rptr[4]\ : SLE
      port map(D => \rptr_s[4]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1006_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[4]_net_1\);
    
    \memwaddr_r_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[4]_net_1\, S => \memwaddr_r_s[5]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[5]_net_1\);
    
    \memraddr_r_s[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[9]_net_1\, S => \memraddr_r_s[10]_net_1\, 
        Y => OPEN, FCO => OPEN);
    
    \wptr_gray[6]\ : SLE
      port map(D => \wptr_gray_1[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[6]_net_1\);
    
    \wptr_gray_1[3]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[3]_net_1\, B => \wptr[4]_net_1\, Y => 
        \wptr_gray_1[3]_net_1\);
    
    \wptr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[4]_net_1\, S
         => \wptr_s[5]\, Y => OPEN, FCO => \wptr_cry[5]_net_1\);
    
    \memraddr_r_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[4]_net_1\, S => \memraddr_r_s[5]\, Y => 
        OPEN, FCO => \memraddr_r_cry[5]_net_1\);
    
    \memraddr_r_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[1]\, C => 
        GND_net_1, D => GND_net_1, FCI => memraddr_r_s_375_FCO, S
         => \memraddr_r_s[1]\, Y => OPEN, FCO => 
        \memraddr_r_cry[1]_net_1\);
    
    \rptr_gray[4]\ : SLE
      port map(D => \rptr_gray_1[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[4]_net_1\);
    
    \wptr_bin_sync2[4]\ : SLE
      port map(D => \wptr_bin_sync[4]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[4]_net_1\);
    
    \wptr[3]\ : SLE
      port map(D => \wptr_s[3]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[3]_net_1\);
    
    \memwaddr_r[6]\ : SLE
      port map(D => \memwaddr_r_s[6]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_249, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[6]\);
    
    rptr_s_374 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => rptr_s_374_FCO);
    
    \wptr_s[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[10]_net_1\, S
         => \wptr_s[11]_net_1\, Y => OPEN, FCO => OPEN);
    
    \wptr[6]\ : SLE
      port map(D => \wptr_s[6]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[6]_net_1\);
    
    \memwaddr_r[9]\ : SLE
      port map(D => \memwaddr_r_s[9]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_249, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[9]\);
    
    \memraddr_r_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[3]_net_1\, S => \memraddr_r_s[4]\, Y => 
        OPEN, FCO => \memraddr_r_cry[4]_net_1\);
    
    empty_r_RNI4GH71 : CFG3
      generic map(INIT => x"A6")

      port map(A => REN_d1, B => N_133, C => \iRX_FIFO_Empty_0\, 
        Y => N_154_i_i);
    
    \memraddr_r[10]\ : SLE
      port map(D => \memraddr_r_s[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1006_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[10]\);
    
    \memwaddr_r[3]\ : SLE
      port map(D => \memwaddr_r_s[3]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_249, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[3]\);
    
    full_r : SLE
      port map(D => fulli, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \iRX_FIFO_Full_0\);
    
    \rptr_bin_sync2[3]\ : SLE
      port map(D => \rptr_bin_sync[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[3]_net_1\);
    
    \wptr_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \wptr[0]_net_1\, Y => \wptr_s[0]\);
    
    \rptr[2]\ : SLE
      port map(D => \rptr_s[2]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1006_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[2]_net_1\);
    
    \memraddr_r[3]\ : SLE
      port map(D => \memraddr_r_s[3]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1006_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[3]\);
    
    \rptr_bin_sync2[9]\ : SLE
      port map(D => \rptr_bin_sync[9]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[9]_net_1\);
    
    \rptr[11]\ : SLE
      port map(D => \rptr_s[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1006_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rptr[11]_net_1\);
    
    memraddr_r_s_375 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[0]\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => memraddr_r_s_375_FCO);
    
    \wptr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[5]_net_1\, S
         => \wptr_s[6]\, Y => OPEN, FCO => \wptr_cry[6]_net_1\);
    
    \rptr_bin_sync2[11]\ : SLE
      port map(D => \rptr_bin_sync[11]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[11]_net_1\);
    
    \wptr_bin_sync2[5]\ : SLE
      port map(D => \wptr_bin_sync[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[5]_net_1\);
    
    \wptr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[7]_net_1\, S
         => \wptr_s[8]\, Y => OPEN, FCO => \wptr_cry[8]_net_1\);
    
    \wptr_bin_sync2[1]\ : SLE
      port map(D => \wptr_bin_sync[1]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[1]_net_1\);
    
    Wr_corefifo_grayToBinConv : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_6
      port map(wptr_bin_sync(11) => \wptr_bin_sync[11]\, 
        wptr_bin_sync(10) => \wptr_bin_sync[10]\, 
        wptr_bin_sync(9) => \wptr_bin_sync[9]\, wptr_bin_sync(8)
         => \wptr_bin_sync[8]\, wptr_bin_sync(7) => 
        \wptr_bin_sync[7]\, wptr_bin_sync(6) => 
        \wptr_bin_sync[6]\, wptr_bin_sync(5) => 
        \wptr_bin_sync[5]\, wptr_bin_sync(4) => 
        \wptr_bin_sync[4]\, wptr_bin_sync(3) => 
        \wptr_bin_sync[3]\, wptr_bin_sync(2) => 
        \wptr_bin_sync[2]\, wptr_bin_sync(1) => 
        \wptr_bin_sync[1]\, wptr_bin_sync(0) => 
        \wptr_bin_sync[0]\, wptr_gray_sync(10) => 
        \wptr_gray_sync[10]\, wptr_gray_sync(9) => 
        \wptr_gray_sync[9]\, wptr_gray_sync(8) => 
        \wptr_gray_sync[8]\, wptr_gray_sync(7) => 
        \wptr_gray_sync[7]\, wptr_gray_sync(6) => 
        \wptr_gray_sync[6]\, wptr_gray_sync(5) => 
        \wptr_gray_sync[5]\, wptr_gray_sync(4) => 
        \wptr_gray_sync[4]\, wptr_gray_sync(3) => 
        \wptr_gray_sync[3]\, wptr_gray_sync(2) => 
        \wptr_gray_sync[2]\, wptr_gray_sync(1) => 
        \wptr_gray_sync[1]\, wptr_gray_sync(0) => 
        \wptr_gray_sync[0]\);
    
    \wptr_gray_1[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[4]_net_1\, B => \wptr[5]_net_1\, Y => 
        \wptr_gray_1[4]_net_1\);
    
    overflow_r : SLE
      port map(D => un1_we_p, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        iRX_FIFO_OVERFLOW_0);
    
    fulli_0 : CFG4
      generic map(INIT => x"EAAA")

      port map(A => \wdiff_bus[11]\, B => \fulli_0_a2_7\, C => 
        N_249, D => \fulli_0_a2_8\, Y => fulli);
    
    \memraddr_r_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \fifo_MEMRADDR[0]\, Y => \memraddr_r_s[0]\);
    
    \rptr_gray[11]\ : SLE
      port map(D => \rptr[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[11]_net_1\);
    
    \wptr_bin_sync2[10]\ : SLE
      port map(D => \wptr_bin_sync[10]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[10]_net_1\);
    
    \rptr[10]\ : SLE
      port map(D => \rptr_s[10]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1006_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rptr[10]_net_1\);
    
    \wptr[9]\ : SLE
      port map(D => \wptr_s[9]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[9]_net_1\);
    
    Wr_corefifo_doubleSync : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_3
      port map(wptr_gray(11) => \wptr_gray[11]_net_1\, 
        wptr_gray(10) => \wptr_gray[10]_net_1\, wptr_gray(9) => 
        \wptr_gray[9]_net_1\, wptr_gray(8) => 
        \wptr_gray[8]_net_1\, wptr_gray(7) => 
        \wptr_gray[7]_net_1\, wptr_gray(6) => 
        \wptr_gray[6]_net_1\, wptr_gray(5) => 
        \wptr_gray[5]_net_1\, wptr_gray(4) => 
        \wptr_gray[4]_net_1\, wptr_gray(3) => 
        \wptr_gray[3]_net_1\, wptr_gray(2) => 
        \wptr_gray[2]_net_1\, wptr_gray(1) => 
        \wptr_gray[1]_net_1\, wptr_gray(0) => 
        \wptr_gray[0]_net_1\, wptr_gray_sync(10) => 
        \wptr_gray_sync[10]\, wptr_gray_sync(9) => 
        \wptr_gray_sync[9]\, wptr_gray_sync(8) => 
        \wptr_gray_sync[8]\, wptr_gray_sync(7) => 
        \wptr_gray_sync[7]\, wptr_gray_sync(6) => 
        \wptr_gray_sync[6]\, wptr_gray_sync(5) => 
        \wptr_gray_sync[5]\, wptr_gray_sync(4) => 
        \wptr_gray_sync[4]\, wptr_gray_sync(3) => 
        \wptr_gray_sync[3]\, wptr_gray_sync(2) => 
        \wptr_gray_sync[2]\, wptr_gray_sync(1) => 
        \wptr_gray_sync[1]\, wptr_gray_sync(0) => 
        \wptr_gray_sync[0]\, wptr_bin_sync_0 => 
        \wptr_bin_sync[11]\, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, irx_fifo_rst_i => 
        irx_fifo_rst_i);
    
    \rptr_gray[0]\ : SLE
      port map(D => \rptr_gray_1[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[0]_net_1\);
    
    empty_r : SLE
      port map(D => empty_r_3, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \iRX_FIFO_Empty_0\);
    
    \rptr_gray_1[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[7]_net_1\, B => \rptr[8]_net_1\, Y => 
        \rptr_gray_1[7]_net_1\);
    
    \wptr[4]\ : SLE
      port map(D => \wptr_s[4]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[4]_net_1\);
    
    \memwaddr_r[8]\ : SLE
      port map(D => \memwaddr_r_s[8]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_249, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[8]\);
    
    \memwaddr_r[2]\ : SLE
      port map(D => \memwaddr_r_s[2]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_249, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[2]\);
    
    \L1.empty_r_3_0_a2_5\ : CFG3
      generic map(INIT => x"0E")

      port map(A => N_133, B => rdiff_bus_cry_0_Y_3, C => 
        \rdiff_bus[11]\, Y => empty_r_3_0_a2_5);
    
    \wptr_bin_sync2[11]\ : SLE
      port map(D => \wptr_bin_sync[11]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[11]_net_1\);
    
    \wptr_gray_1[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[1]_net_1\, B => \wptr[2]_net_1\, Y => 
        \wptr_gray_1[1]_net_1\);
    
    underflow_r : SLE
      port map(D => un2_re_p_i_i_a3_2, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => iRX_FIFO_UNDERRUN_0);
    
    \memwaddr_r_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[6]_net_1\, S => \memwaddr_r_s[7]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[7]_net_1\);
    
    \wptr_gray[5]\ : SLE
      port map(D => \wptr_gray_1[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[5]_net_1\);
    
    \memraddr_r[7]\ : SLE
      port map(D => \memraddr_r_s[7]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1006_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[7]\);
    
    memwe_0_a2_0_a2 : CFG4
      generic map(INIT => x"2000")

      port map(A => ReadFIFO_Write_Ptr(1), B => \iRX_FIFO_Full_0\, 
        C => N_1466, D => ReadFIFO_Write_Ptr(0), Y => 
        \fifo_MEMWE\);
    
    \rptr_bin_sync2[10]\ : SLE
      port map(D => \rptr_bin_sync[10]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[10]_net_1\);
    
    wdiff_bus_cry_10 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[10]_net_1\, B => 
        \rptr_bin_sync2[10]_net_1\, C => GND_net_1, D => 
        GND_net_1, FCI => \wdiff_bus_cry_9\, S => \wdiff_bus[10]\, 
        Y => OPEN, FCO => \wdiff_bus_cry_10\);
    
    \memwaddr_r_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[9]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[8]_net_1\, S => \memwaddr_r_s[9]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[9]_net_1\);
    
    \wptr_gray[8]\ : SLE
      port map(D => \wptr_gray_1[8]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[8]_net_1\);
    
    \wptr_gray[7]\ : SLE
      port map(D => \wptr_gray_1[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[7]_net_1\);
    
    \wptr_gray_1[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[5]_net_1\, B => \wptr[6]_net_1\, Y => 
        \wptr_gray_1[5]_net_1\);
    
    \memwaddr_r[5]\ : SLE
      port map(D => \memwaddr_r_s[5]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_249, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[5]\);
    
    \L1.empty_r_3_0_a2\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \rdiff_bus[9]\, B => \rdiff_bus[10]\, C => 
        empty_r_3_0_a2_5, D => empty_r_3_0_a2_9, Y => empty_r_3);
    
    \rptr[8]\ : SLE
      port map(D => \rptr_s[8]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1006_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[8]_net_1\);
    
    Rd_corefifo_doubleSync : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_2
      port map(rptr_gray(11) => \rptr_gray[11]_net_1\, 
        rptr_gray(10) => \rptr_gray[10]_net_1\, rptr_gray(9) => 
        \rptr_gray[9]_net_1\, rptr_gray(8) => 
        \rptr_gray[8]_net_1\, rptr_gray(7) => 
        \rptr_gray[7]_net_1\, rptr_gray(6) => 
        \rptr_gray[6]_net_1\, rptr_gray(5) => 
        \rptr_gray[5]_net_1\, rptr_gray(4) => 
        \rptr_gray[4]_net_1\, rptr_gray(3) => 
        \rptr_gray[3]_net_1\, rptr_gray(2) => 
        \rptr_gray[2]_net_1\, rptr_gray(1) => 
        \rptr_gray[1]_net_1\, rptr_gray(0) => 
        \rptr_gray[0]_net_1\, rptr_gray_sync(10) => 
        \rptr_gray_sync[10]\, rptr_gray_sync(9) => 
        \rptr_gray_sync[9]\, rptr_gray_sync(8) => 
        \rptr_gray_sync[8]\, rptr_gray_sync(7) => 
        \rptr_gray_sync[7]\, rptr_gray_sync(6) => 
        \rptr_gray_sync[6]\, rptr_gray_sync(5) => 
        \rptr_gray_sync[5]\, rptr_gray_sync(4) => 
        \rptr_gray_sync[4]\, rptr_gray_sync(3) => 
        \rptr_gray_sync[3]\, rptr_gray_sync(2) => 
        \rptr_gray_sync[2]\, rptr_gray_sync(1) => 
        \rptr_gray_sync[1]\, rptr_gray_sync(0) => 
        \rptr_gray_sync[0]\, rptr_bin_sync_0 => 
        \rptr_bin_sync[11]\, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, irx_fifo_rst_i => irx_fifo_rst_i);
    
    \rptr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[3]_net_1\, S
         => \rptr_s[4]\, Y => OPEN, FCO => \rptr_cry[4]_net_1\);
    
    wdiff_bus_cry_2 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[2]_net_1\, B => 
        \rptr_bin_sync2[2]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_1\, S => \wdiff_bus[2]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_2\);
    
    \rptr_gray[2]\ : SLE
      port map(D => \rptr_gray_1[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[2]_net_1\);
    
    \wptr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[8]_net_1\, S
         => \wptr_s[9]\, Y => OPEN, FCO => \wptr_cry[9]_net_1\);
    
    \wptr_bin_sync2[3]\ : SLE
      port map(D => \wptr_bin_sync[3]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[3]_net_1\);
    
    \wptr[2]\ : SLE
      port map(D => \wptr_s[2]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[2]_net_1\);
    
    \rptr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[1]_net_1\, S
         => \rptr_s[2]\, Y => OPEN, FCO => \rptr_cry[2]_net_1\);
    
    rdiff_bus_cry_9 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[9]_net_1\, B => 
        \rptr[9]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_8\, S => \rdiff_bus[9]\, Y => OPEN, FCO
         => \rdiff_bus_cry_9\);
    
    \memwaddr_r[0]\ : SLE
      port map(D => \memwaddr_r_s[0]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_249, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[0]\);
    
    fulli_0_a2_7 : CFG4
      generic map(INIT => x"8000")

      port map(A => \wdiff_bus[6]\, B => \wdiff_bus[7]\, C => 
        \wdiff_bus[8]\, D => \wdiff_bus[9]\, Y => \fulli_0_a2_7\);
    
    \wptr_gray[2]\ : SLE
      port map(D => \wptr_gray_1[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[2]_net_1\);
    
    wdiff_bus_cry_4 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[4]_net_1\, B => 
        \rptr_bin_sync2[4]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_3\, S => \wdiff_bus[4]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_4\);
    
    \memwaddr_r_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[2]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[1]_net_1\, S => \memwaddr_r_s[2]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[2]_net_1\);
    
    \wptr_gray[11]\ : SLE
      port map(D => \wptr[11]_net_1\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr_gray[11]_net_1\);
    
    \wptr_bin_sync2[9]\ : SLE
      port map(D => \wptr_bin_sync[9]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[9]_net_1\);
    
    \rptr_gray_1[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[6]_net_1\, B => \rptr[7]_net_1\, Y => 
        \rptr_gray_1[6]_net_1\);
    
    \wptr_gray_1[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[11]_net_1\, B => \wptr[10]_net_1\, Y
         => \wptr_gray_1[10]_net_1\);
    
    wdiff_bus_cry_6 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[6]_net_1\, B => 
        \rptr_bin_sync2[6]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_5\, S => \wdiff_bus[6]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_6\);
    
    \rptr_s[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[10]_net_1\, S
         => \rptr_s[11]_net_1\, Y => OPEN, FCO => OPEN);
    
    \rptr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[2]_net_1\, S
         => \rptr_s[3]\, Y => OPEN, FCO => \rptr_cry[3]_net_1\);
    
    \memraddr_r[4]\ : SLE
      port map(D => \memraddr_r_s[4]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1006_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[4]\);
    
    wptr_s_376 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => wptr_s_376_FCO);
    
    \memraddr_r_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[6]_net_1\, S => \memraddr_r_s[7]\, Y => 
        OPEN, FCO => \memraddr_r_cry[7]_net_1\);
    
    fulli_0_a2_8 : CFG4
      generic map(INIT => x"4000")

      port map(A => wdiff_bus_cry_0_Y_3, B => \wdiff_bus[1]\, C
         => \wdiff_bus[10]\, D => \fulli_0_a2_6\, Y => 
        \fulli_0_a2_8\);
    
    empty_r_RNI3NBU : CFG2
      generic map(INIT => x"2")

      port map(A => N_133, B => \iRX_FIFO_Empty_0\, Y => 
        \N_1006_i\);
    
    \memraddr_r_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[9]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[8]_net_1\, S => \memraddr_r_s[9]\, Y => 
        OPEN, FCO => \memraddr_r_cry[9]_net_1\);
    
    \memraddr_r[5]\ : SLE
      port map(D => \memraddr_r_s[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1006_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[5]\);
    
    \rptr_gray[6]\ : SLE
      port map(D => \rptr_gray_1[6]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[6]_net_1\);
    
    \memraddr_r[9]\ : SLE
      port map(D => \memraddr_r_s[9]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1006_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[9]\);
    
    \rptr[0]\ : SLE
      port map(D => \rptr_s[0]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1006_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[0]_net_1\);
    
    \wptr[10]\ : SLE
      port map(D => \wptr_s[10]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[10]_net_1\);
    
    \memwaddr_r_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[3]_net_1\, S => \memwaddr_r_s[4]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[4]_net_1\);
    
    \memraddr_r_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[3]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[2]_net_1\, S => \memraddr_r_s[3]\, Y => 
        OPEN, FCO => \memraddr_r_cry[3]_net_1\);
    
    wdiff_bus_cry_1 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[1]_net_1\, B => 
        \rptr_bin_sync2[1]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_0\, S => \wdiff_bus[1]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_1\);
    
    rdiff_bus_cry_2 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[2]_net_1\, B => 
        \rptr[2]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_1\, S => \rdiff_bus[2]\, Y => OPEN, FCO
         => \rdiff_bus_cry_2\);
    
    \wptr_gray[9]\ : SLE
      port map(D => \wptr_gray_1[9]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[9]_net_1\);
    
    \rptr_gray_1[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[4]_net_1\, B => \rptr[5]_net_1\, Y => 
        \rptr_gray_1[4]_net_1\);
    
    \wptr_gray_1[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[8]_net_1\, B => \wptr[9]_net_1\, Y => 
        \wptr_gray_1[8]_net_1\);
    
    Rd_corefifo_grayToBinConv : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_5
      port map(rptr_bin_sync(11) => \rptr_bin_sync[11]\, 
        rptr_bin_sync(10) => \rptr_bin_sync[10]\, 
        rptr_bin_sync(9) => \rptr_bin_sync[9]\, rptr_bin_sync(8)
         => \rptr_bin_sync[8]\, rptr_bin_sync(7) => 
        \rptr_bin_sync[7]\, rptr_bin_sync(6) => 
        \rptr_bin_sync[6]\, rptr_bin_sync(5) => 
        \rptr_bin_sync[5]\, rptr_bin_sync(4) => 
        \rptr_bin_sync[4]\, rptr_bin_sync(3) => 
        \rptr_bin_sync[3]\, rptr_bin_sync(2) => 
        \rptr_bin_sync[2]\, rptr_bin_sync(1) => 
        \rptr_bin_sync[1]\, rptr_bin_sync(0) => 
        \rptr_bin_sync[0]\, rptr_gray_sync(10) => 
        \rptr_gray_sync[10]\, rptr_gray_sync(9) => 
        \rptr_gray_sync[9]\, rptr_gray_sync(8) => 
        \rptr_gray_sync[8]\, rptr_gray_sync(7) => 
        \rptr_gray_sync[7]\, rptr_gray_sync(6) => 
        \rptr_gray_sync[6]\, rptr_gray_sync(5) => 
        \rptr_gray_sync[5]\, rptr_gray_sync(4) => 
        \rptr_gray_sync[4]\, rptr_gray_sync(3) => 
        \rptr_gray_sync[3]\, rptr_gray_sync(2) => 
        \rptr_gray_sync[2]\, rptr_gray_sync(1) => 
        \rptr_gray_sync[1]\, rptr_gray_sync(0) => 
        \rptr_gray_sync[0]\);
    
    \rptr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => rptr_s_374_FCO, S => 
        \rptr_s[1]\, Y => OPEN, FCO => \rptr_cry[1]_net_1\);
    
    rdiff_bus_cry_3 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[3]_net_1\, B => 
        \rptr[3]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_2\, S => \rdiff_bus[3]\, Y => OPEN, FCO
         => \rdiff_bus_cry_3\);
    
    rdiff_bus_cry_10 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[10]_net_1\, B => 
        \rptr[10]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_9\, S => \rdiff_bus[10]\, Y => OPEN, FCO
         => \rdiff_bus_cry_10\);
    
    \memraddr_r_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[5]_net_1\, S => \memraddr_r_s[6]\, Y => 
        OPEN, FCO => \memraddr_r_cry[6]_net_1\);
    
    \memraddr_r[6]\ : SLE
      port map(D => \memraddr_r_s[6]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1006_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[6]\);
    
    \rptr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[6]_net_1\, S
         => \rptr_s[7]\, Y => OPEN, FCO => \rptr_cry[7]_net_1\);
    
    rdiff_bus_cry_0 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => rdiff_bus, B => \rptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => rdiff_bus_cry_0_Y_3, FCO => \rdiff_bus_cry_0\);
    
    \memraddr_r[2]\ : SLE
      port map(D => \memraddr_r_s[2]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1006_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[2]\);
    
    \wptr[8]\ : SLE
      port map(D => \wptr_s[8]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[8]_net_1\);
    
    wdiff_bus_cry_3 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[3]_net_1\, B => 
        \rptr_bin_sync2[3]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_2\, S => \wdiff_bus[3]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_3\);
    
    \rptr_gray[7]\ : SLE
      port map(D => \rptr_gray_1[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[7]_net_1\);
    
    \wptr_gray[0]\ : SLE
      port map(D => \wptr_gray_1[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[0]_net_1\);
    
    \rptr_gray_1[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[0]_net_1\, B => \rptr[1]_net_1\, Y => 
        \rptr_gray_1[0]_net_1\);
    
    \rptr_gray_1[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[8]_net_1\, B => \rptr[9]_net_1\, Y => 
        \rptr_gray_1[8]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_2 is

    port( RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          ReadFIFO_Write_Ptr        : in    std_logic_vector(1 downto 0);
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          RX_FIFO_DOUT_3_0          : out   std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          N_1466                    : in    std_logic;
          N_674                     : out   std_logic;
          N_676                     : out   std_logic;
          N_715                     : out   std_logic;
          N_677                     : out   std_logic;
          N_675                     : out   std_logic;
          N_673                     : out   std_logic;
          N_672                     : out   std_logic;
          N_671                     : out   std_logic;
          N_133                     : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          irx_fifo_rst_i            : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_2;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_2 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_2
    port( RDATA_int                 : out   std_logic_vector(8 downto 0);
          fifo_MEMRADDR             : in    std_logic_vector(10 downto 0) := (others => 'U');
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          fifo_MEMWADDR             : in    std_logic_vector(10 downto 0) := (others => 'U');
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          N_1006_i                  : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          fifo_MEMWE                : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_2
    port( ReadFIFO_Write_Ptr        : in    std_logic_vector(1 downto 0) := (others => 'U');
          fifo_MEMWADDR             : out   std_logic_vector(10 downto 0);
          fifo_MEMRADDR             : out   std_logic_vector(10 downto 0);
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          N_154_i_i                 : out   std_logic;
          N_89_i                    : out   std_logic;
          REN_d1                    : in    std_logic := 'U';
          N_133                     : in    std_logic := 'U';
          N_1466                    : in    std_logic := 'U';
          N_1006_i                  : out   std_logic;
          fifo_MEMWE                : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          irx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \RDATA_r[4]_net_1\, VCC_net_1, \RDATA_int[4]\, N_89_i, 
        GND_net_1, \RDATA_r[5]_net_1\, \RDATA_int[5]\, 
        \RDATA_r[6]_net_1\, \RDATA_int[6]\, \RDATA_r[7]_net_1\, 
        \RDATA_int[7]\, \RDATA_r[8]_net_1\, \RDATA_int[8]\, 
        \re_set\, \REN_d1\, N_154_i_i, \RDATA_r[0]_net_1\, 
        \RDATA_int[0]\, \RDATA_r[1]_net_1\, \RDATA_int[1]\, 
        \RDATA_r[2]_net_1\, \RDATA_int[2]\, \RDATA_r[3]_net_1\, 
        \RDATA_int[3]\, N_1006_i, \RE_d1\, \re_pulse_d1\, 
        \re_pulse\, \iRX_FIFO_Empty_0\, \fifo_MEMWADDR[0]\, 
        \fifo_MEMWADDR[1]\, \fifo_MEMWADDR[2]\, 
        \fifo_MEMWADDR[3]\, \fifo_MEMWADDR[4]\, 
        \fifo_MEMWADDR[5]\, \fifo_MEMWADDR[6]\, 
        \fifo_MEMWADDR[7]\, \fifo_MEMWADDR[8]\, 
        \fifo_MEMWADDR[9]\, \fifo_MEMWADDR[10]\, 
        \fifo_MEMRADDR[0]\, \fifo_MEMRADDR[1]\, 
        \fifo_MEMRADDR[2]\, \fifo_MEMRADDR[3]\, 
        \fifo_MEMRADDR[4]\, \fifo_MEMRADDR[5]\, 
        \fifo_MEMRADDR[6]\, \fifo_MEMRADDR[7]\, 
        \fifo_MEMRADDR[8]\, \fifo_MEMRADDR[9]\, 
        \fifo_MEMRADDR[10]\, fifo_MEMWE : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_2
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_2(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_2
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_2(DEF_ARCH);
begin 

    iRX_FIFO_Empty_0 <= \iRX_FIFO_Empty_0\;

    re_pulse : CFG4
      generic map(INIT => x"FAF2")

      port map(A => \REN_d1\, B => N_133, C => \re_set\, D => 
        \iRX_FIFO_Empty_0\, Y => \re_pulse\);
    
    \RDATA_r[3]\ : SLE
      port map(D => \RDATA_int[3]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[3]_net_1\);
    
    \Q_i_m2[2]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[2]_net_1\, C => 
        \RDATA_int[2]\, D => \RE_d1\, Y => N_672);
    
    re_pulse_d1 : SLE
      port map(D => \re_pulse\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \re_pulse_d1\);
    
    \RDATA_r[5]\ : SLE
      port map(D => \RDATA_int[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[5]_net_1\);
    
    \Q_i_m2[0]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[0]_net_1\, C => 
        \RDATA_int[0]\, D => \RE_d1\, Y => N_671);
    
    \Q_i_m2[3]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[3]_net_1\, C => 
        \RDATA_int[3]\, D => \RE_d1\, Y => N_673);
    
    \RDATA_r[8]\ : SLE
      port map(D => \RDATA_int[8]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[8]_net_1\);
    
    \Q_i_m2[7]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[7]_net_1\, C => 
        \RDATA_int[7]\, D => \RE_d1\, Y => N_677);
    
    \Q_i_m2[6]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[6]_net_1\, C => 
        \RDATA_int[6]\, D => \RE_d1\, Y => N_676);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \RW1.UI_ram_wrapper_1\ : FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_2
      port map(RDATA_int(8) => \RDATA_int[8]\, RDATA_int(7) => 
        \RDATA_int[7]\, RDATA_int(6) => \RDATA_int[6]\, 
        RDATA_int(5) => \RDATA_int[5]\, RDATA_int(4) => 
        \RDATA_int[4]\, RDATA_int(3) => \RDATA_int[3]\, 
        RDATA_int(2) => \RDATA_int[2]\, RDATA_int(1) => 
        \RDATA_int[1]\, RDATA_int(0) => \RDATA_int[0]\, 
        fifo_MEMRADDR(10) => \fifo_MEMRADDR[10]\, 
        fifo_MEMRADDR(9) => \fifo_MEMRADDR[9]\, fifo_MEMRADDR(8)
         => \fifo_MEMRADDR[8]\, fifo_MEMRADDR(7) => 
        \fifo_MEMRADDR[7]\, fifo_MEMRADDR(6) => 
        \fifo_MEMRADDR[6]\, fifo_MEMRADDR(5) => 
        \fifo_MEMRADDR[5]\, fifo_MEMRADDR(4) => 
        \fifo_MEMRADDR[4]\, fifo_MEMRADDR(3) => 
        \fifo_MEMRADDR[3]\, fifo_MEMRADDR(2) => 
        \fifo_MEMRADDR[2]\, fifo_MEMRADDR(1) => 
        \fifo_MEMRADDR[1]\, fifo_MEMRADDR(0) => 
        \fifo_MEMRADDR[0]\, RX_FIFO_DIN_pipe(8) => 
        RX_FIFO_DIN_pipe(8), RX_FIFO_DIN_pipe(7) => 
        RX_FIFO_DIN_pipe(7), RX_FIFO_DIN_pipe(6) => 
        RX_FIFO_DIN_pipe(6), RX_FIFO_DIN_pipe(5) => 
        RX_FIFO_DIN_pipe(5), RX_FIFO_DIN_pipe(4) => 
        RX_FIFO_DIN_pipe(4), RX_FIFO_DIN_pipe(3) => 
        RX_FIFO_DIN_pipe(3), RX_FIFO_DIN_pipe(2) => 
        RX_FIFO_DIN_pipe(2), RX_FIFO_DIN_pipe(1) => 
        RX_FIFO_DIN_pipe(1), RX_FIFO_DIN_pipe(0) => 
        RX_FIFO_DIN_pipe(0), fifo_MEMWADDR(10) => 
        \fifo_MEMWADDR[10]\, fifo_MEMWADDR(9) => 
        \fifo_MEMWADDR[9]\, fifo_MEMWADDR(8) => 
        \fifo_MEMWADDR[8]\, fifo_MEMWADDR(7) => 
        \fifo_MEMWADDR[7]\, fifo_MEMWADDR(6) => 
        \fifo_MEMWADDR[6]\, fifo_MEMWADDR(5) => 
        \fifo_MEMWADDR[5]\, fifo_MEMWADDR(4) => 
        \fifo_MEMWADDR[4]\, fifo_MEMWADDR(3) => 
        \fifo_MEMWADDR[3]\, fifo_MEMWADDR(2) => 
        \fifo_MEMWADDR[2]\, fifo_MEMWADDR(1) => 
        \fifo_MEMWADDR[1]\, fifo_MEMWADDR(0) => 
        \fifo_MEMWADDR[0]\, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, N_1006_i => N_1006_i, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, fifo_MEMWE
         => fifo_MEMWE);
    
    \RDATA_r[0]\ : SLE
      port map(D => \RDATA_int[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[0]_net_1\);
    
    \Q_i_m2[5]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[5]_net_1\, C => 
        \RDATA_int[5]\, D => \RE_d1\, Y => N_675);
    
    \RDATA_r[2]\ : SLE
      port map(D => \RDATA_int[2]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[2]_net_1\);
    
    \RDATA_r[6]\ : SLE
      port map(D => \RDATA_int[6]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[6]_net_1\);
    
    \L31.U_corefifo_async\ : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_2
      port map(ReadFIFO_Write_Ptr(1) => ReadFIFO_Write_Ptr(1), 
        ReadFIFO_Write_Ptr(0) => ReadFIFO_Write_Ptr(0), 
        fifo_MEMWADDR(10) => \fifo_MEMWADDR[10]\, 
        fifo_MEMWADDR(9) => \fifo_MEMWADDR[9]\, fifo_MEMWADDR(8)
         => \fifo_MEMWADDR[8]\, fifo_MEMWADDR(7) => 
        \fifo_MEMWADDR[7]\, fifo_MEMWADDR(6) => 
        \fifo_MEMWADDR[6]\, fifo_MEMWADDR(5) => 
        \fifo_MEMWADDR[5]\, fifo_MEMWADDR(4) => 
        \fifo_MEMWADDR[4]\, fifo_MEMWADDR(3) => 
        \fifo_MEMWADDR[3]\, fifo_MEMWADDR(2) => 
        \fifo_MEMWADDR[2]\, fifo_MEMWADDR(1) => 
        \fifo_MEMWADDR[1]\, fifo_MEMWADDR(0) => 
        \fifo_MEMWADDR[0]\, fifo_MEMRADDR(10) => 
        \fifo_MEMRADDR[10]\, fifo_MEMRADDR(9) => 
        \fifo_MEMRADDR[9]\, fifo_MEMRADDR(8) => 
        \fifo_MEMRADDR[8]\, fifo_MEMRADDR(7) => 
        \fifo_MEMRADDR[7]\, fifo_MEMRADDR(6) => 
        \fifo_MEMRADDR[6]\, fifo_MEMRADDR(5) => 
        \fifo_MEMRADDR[5]\, fifo_MEMRADDR(4) => 
        \fifo_MEMRADDR[4]\, fifo_MEMRADDR(3) => 
        \fifo_MEMRADDR[3]\, fifo_MEMRADDR(2) => 
        \fifo_MEMRADDR[2]\, fifo_MEMRADDR(1) => 
        \fifo_MEMRADDR[1]\, fifo_MEMRADDR(0) => 
        \fifo_MEMRADDR[0]\, iRX_FIFO_Empty_0 => 
        \iRX_FIFO_Empty_0\, iRX_FIFO_UNDERRUN_0 => 
        iRX_FIFO_UNDERRUN_0, iRX_FIFO_Full_0 => iRX_FIFO_Full_0, 
        iRX_FIFO_OVERFLOW_0 => iRX_FIFO_OVERFLOW_0, N_154_i_i => 
        N_154_i_i, N_89_i => N_89_i, REN_d1 => \REN_d1\, N_133
         => N_133, N_1466 => N_1466, N_1006_i => N_1006_i, 
        fifo_MEMWE => fifo_MEMWE, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, irx_fifo_rst_i => irx_fifo_rst_i);
    
    re_set : SLE
      port map(D => \REN_d1\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => N_154_i_i, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \re_set\);
    
    \Q_i_m2[8]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[8]_net_1\, C => 
        \RDATA_int[8]\, D => \RE_d1\, Y => N_715);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    RE_d1 : SLE
      port map(D => N_133, CLK => m2s010_som_sb_0_CCC_71MHz, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \RE_d1\);
    
    \RDATA_r[7]\ : SLE
      port map(D => \RDATA_int[7]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[7]_net_1\);
    
    \RDATA_r[4]\ : SLE
      port map(D => \RDATA_int[4]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[4]_net_1\);
    
    \Q[1]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[1]_net_1\, C => 
        \RDATA_int[1]\, D => \RE_d1\, Y => RX_FIFO_DOUT_3_0);
    
    REN_d1 : SLE
      port map(D => N_1006_i, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \REN_d1\);
    
    \Q_i_m2[4]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[4]_net_1\, C => 
        \RDATA_int[4]\, D => \RE_d1\, Y => N_674);
    
    \RDATA_r[1]\ : SLE
      port map(D => \RDATA_int[1]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[1]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_2 is

    port( ReadFIFO_Write_Ptr        : in    std_logic_vector(1 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          RX_FIFO_DOUT_3_0          : out   std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          irx_fifo_rst_i            : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          N_133                     : in    std_logic;
          N_671                     : out   std_logic;
          N_672                     : out   std_logic;
          N_673                     : out   std_logic;
          N_675                     : out   std_logic;
          N_677                     : out   std_logic;
          N_715                     : out   std_logic;
          N_676                     : out   std_logic;
          N_674                     : out   std_logic;
          N_1466                    : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic
        );

end FIFO_8Kx9_2;

architecture DEF_ARCH of FIFO_8Kx9_2 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_2
    port( RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          ReadFIFO_Write_Ptr        : in    std_logic_vector(1 downto 0) := (others => 'U');
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          RX_FIFO_DOUT_3_0          : out   std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          N_1466                    : in    std_logic := 'U';
          N_674                     : out   std_logic;
          N_676                     : out   std_logic;
          N_715                     : out   std_logic;
          N_677                     : out   std_logic;
          N_675                     : out   std_logic;
          N_673                     : out   std_logic;
          N_672                     : out   std_logic;
          N_671                     : out   std_logic;
          N_133                     : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          irx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_2
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_2(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    FIFO_8Kx9_0 : FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_2
      port map(RX_FIFO_DIN_pipe(8) => RX_FIFO_DIN_pipe(8), 
        RX_FIFO_DIN_pipe(7) => RX_FIFO_DIN_pipe(7), 
        RX_FIFO_DIN_pipe(6) => RX_FIFO_DIN_pipe(6), 
        RX_FIFO_DIN_pipe(5) => RX_FIFO_DIN_pipe(5), 
        RX_FIFO_DIN_pipe(4) => RX_FIFO_DIN_pipe(4), 
        RX_FIFO_DIN_pipe(3) => RX_FIFO_DIN_pipe(3), 
        RX_FIFO_DIN_pipe(2) => RX_FIFO_DIN_pipe(2), 
        RX_FIFO_DIN_pipe(1) => RX_FIFO_DIN_pipe(1), 
        RX_FIFO_DIN_pipe(0) => RX_FIFO_DIN_pipe(0), 
        ReadFIFO_Write_Ptr(1) => ReadFIFO_Write_Ptr(1), 
        ReadFIFO_Write_Ptr(0) => ReadFIFO_Write_Ptr(0), 
        iRX_FIFO_OVERFLOW_0 => iRX_FIFO_OVERFLOW_0, 
        iRX_FIFO_Full_0 => iRX_FIFO_Full_0, iRX_FIFO_UNDERRUN_0
         => iRX_FIFO_UNDERRUN_0, iRX_FIFO_Empty_0 => 
        iRX_FIFO_Empty_0, RX_FIFO_DOUT_3_0 => RX_FIFO_DOUT_3_0, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, N_1466 => 
        N_1466, N_674 => N_674, N_676 => N_676, N_715 => N_715, 
        N_677 => N_677, N_675 => N_675, N_673 => N_673, N_672 => 
        N_672, N_671 => N_671, N_133 => N_133, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz, 
        irx_fifo_rst_i => irx_fifo_rst_i);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top is

    port( fifo_MEMWADDR             : in    std_logic_vector(10 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          fifo_MEMRADDR             : in    std_logic_vector(10 downto 0);
          RDATA_int                 : out   std_logic_vector(8 downto 0);
          fifo_MEMWE                : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          N_1007_i                  : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component RAM1K18
    generic (MEMORYFILE:string := "");

    port( A_DOUT        : out   std_logic_vector(17 downto 0);
          B_DOUT        : out   std_logic_vector(17 downto 0);
          BUSY          : out   std_logic;
          A_CLK         : in    std_logic := 'U';
          A_DOUT_CLK    : in    std_logic := 'U';
          A_ARST_N      : in    std_logic := 'U';
          A_DOUT_EN     : in    std_logic := 'U';
          A_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_DOUT_ARST_N : in    std_logic := 'U';
          A_DOUT_SRST_N : in    std_logic := 'U';
          A_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          A_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          A_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          B_CLK         : in    std_logic := 'U';
          B_DOUT_CLK    : in    std_logic := 'U';
          B_ARST_N      : in    std_logic := 'U';
          B_DOUT_EN     : in    std_logic := 'U';
          B_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_DOUT_ARST_N : in    std_logic := 'U';
          B_DOUT_SRST_N : in    std_logic := 'U';
          B_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          B_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          B_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          A_EN          : in    std_logic := 'U';
          A_DOUT_LAT    : in    std_logic := 'U';
          A_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_WMODE       : in    std_logic := 'U';
          B_EN          : in    std_logic := 'U';
          B_DOUT_LAT    : in    std_logic := 'U';
          B_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_WMODE       : in    std_logic := 'U';
          SII_LOCK      : in    std_logic := 'U'
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;
    signal nc24, nc1, nc8, nc13, nc16, nc19, nc25, nc20, nc27, 
        nc9, nc22, nc14, nc5, nc21, nc15, nc3, nc10, nc7, nc17, 
        nc4, nc12, nc2, nc23, nc18, nc26, nc6, nc11 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C0 : RAM1K18
      port map(A_DOUT(17) => nc24, A_DOUT(16) => nc1, A_DOUT(15)
         => nc8, A_DOUT(14) => nc13, A_DOUT(13) => nc16, 
        A_DOUT(12) => nc19, A_DOUT(11) => nc25, A_DOUT(10) => 
        nc20, A_DOUT(9) => nc27, A_DOUT(8) => RDATA_int(8), 
        A_DOUT(7) => RDATA_int(7), A_DOUT(6) => RDATA_int(6), 
        A_DOUT(5) => RDATA_int(5), A_DOUT(4) => RDATA_int(4), 
        A_DOUT(3) => RDATA_int(3), A_DOUT(2) => RDATA_int(2), 
        A_DOUT(1) => RDATA_int(1), A_DOUT(0) => RDATA_int(0), 
        B_DOUT(17) => nc9, B_DOUT(16) => nc22, B_DOUT(15) => nc14, 
        B_DOUT(14) => nc5, B_DOUT(13) => nc21, B_DOUT(12) => nc15, 
        B_DOUT(11) => nc3, B_DOUT(10) => nc10, B_DOUT(9) => nc7, 
        B_DOUT(8) => nc17, B_DOUT(7) => nc4, B_DOUT(6) => nc12, 
        B_DOUT(5) => nc2, B_DOUT(4) => nc23, B_DOUT(3) => nc18, 
        B_DOUT(2) => nc26, B_DOUT(1) => nc6, B_DOUT(0) => nc11, 
        BUSY => OPEN, A_CLK => m2s010_som_sb_0_CCC_71MHz, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => VCC_net_1, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => N_1007_i, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => GND_net_1, A_DIN(15) => GND_net_1, 
        A_DIN(14) => GND_net_1, A_DIN(13) => GND_net_1, A_DIN(12)
         => GND_net_1, A_DIN(11) => GND_net_1, A_DIN(10) => 
        GND_net_1, A_DIN(9) => GND_net_1, A_DIN(8) => GND_net_1, 
        A_DIN(7) => GND_net_1, A_DIN(6) => GND_net_1, A_DIN(5)
         => GND_net_1, A_DIN(4) => GND_net_1, A_DIN(3) => 
        GND_net_1, A_DIN(2) => GND_net_1, A_DIN(1) => GND_net_1, 
        A_DIN(0) => GND_net_1, A_ADDR(13) => fifo_MEMRADDR(10), 
        A_ADDR(12) => fifo_MEMRADDR(9), A_ADDR(11) => 
        fifo_MEMRADDR(8), A_ADDR(10) => fifo_MEMRADDR(7), 
        A_ADDR(9) => fifo_MEMRADDR(6), A_ADDR(8) => 
        fifo_MEMRADDR(5), A_ADDR(7) => fifo_MEMRADDR(4), 
        A_ADDR(6) => fifo_MEMRADDR(3), A_ADDR(5) => 
        fifo_MEMRADDR(2), A_ADDR(4) => fifo_MEMRADDR(1), 
        A_ADDR(3) => fifo_MEMRADDR(0), A_ADDR(2) => GND_net_1, 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => RX_FIFO_DIN_pipe(8), B_DIN(7) => RX_FIFO_DIN_pipe(7), 
        B_DIN(6) => RX_FIFO_DIN_pipe(6), B_DIN(5) => 
        RX_FIFO_DIN_pipe(5), B_DIN(4) => RX_FIFO_DIN_pipe(4), 
        B_DIN(3) => RX_FIFO_DIN_pipe(3), B_DIN(2) => 
        RX_FIFO_DIN_pipe(2), B_DIN(1) => RX_FIFO_DIN_pipe(1), 
        B_DIN(0) => RX_FIFO_DIN_pipe(0), B_ADDR(13) => 
        fifo_MEMWADDR(10), B_ADDR(12) => fifo_MEMWADDR(9), 
        B_ADDR(11) => fifo_MEMWADDR(8), B_ADDR(10) => 
        fifo_MEMWADDR(7), B_ADDR(9) => fifo_MEMWADDR(6), 
        B_ADDR(8) => fifo_MEMWADDR(5), B_ADDR(7) => 
        fifo_MEMWADDR(4), B_ADDR(6) => fifo_MEMWADDR(3), 
        B_ADDR(5) => fifo_MEMWADDR(2), B_ADDR(4) => 
        fifo_MEMWADDR(1), B_ADDR(3) => fifo_MEMWADDR(0), 
        B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, B_ADDR(0)
         => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0) => 
        VCC_net_1, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper is

    port( RDATA_int                 : out   std_logic_vector(8 downto 0);
          fifo_MEMRADDR             : in    std_logic_vector(10 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          fifo_MEMWADDR             : in    std_logic_vector(10 downto 0);
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          N_1007_i                  : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          fifo_MEMWE                : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top
    port( fifo_MEMWADDR             : in    std_logic_vector(10 downto 0) := (others => 'U');
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          fifo_MEMRADDR             : in    std_logic_vector(10 downto 0) := (others => 'U');
          RDATA_int                 : out   std_logic_vector(8 downto 0);
          fifo_MEMWE                : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          N_1007_i                  : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    L1_asyncnonpipe : FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top
      port map(fifo_MEMWADDR(10) => fifo_MEMWADDR(10), 
        fifo_MEMWADDR(9) => fifo_MEMWADDR(9), fifo_MEMWADDR(8)
         => fifo_MEMWADDR(8), fifo_MEMWADDR(7) => 
        fifo_MEMWADDR(7), fifo_MEMWADDR(6) => fifo_MEMWADDR(6), 
        fifo_MEMWADDR(5) => fifo_MEMWADDR(5), fifo_MEMWADDR(4)
         => fifo_MEMWADDR(4), fifo_MEMWADDR(3) => 
        fifo_MEMWADDR(3), fifo_MEMWADDR(2) => fifo_MEMWADDR(2), 
        fifo_MEMWADDR(1) => fifo_MEMWADDR(1), fifo_MEMWADDR(0)
         => fifo_MEMWADDR(0), RX_FIFO_DIN_pipe(8) => 
        RX_FIFO_DIN_pipe(8), RX_FIFO_DIN_pipe(7) => 
        RX_FIFO_DIN_pipe(7), RX_FIFO_DIN_pipe(6) => 
        RX_FIFO_DIN_pipe(6), RX_FIFO_DIN_pipe(5) => 
        RX_FIFO_DIN_pipe(5), RX_FIFO_DIN_pipe(4) => 
        RX_FIFO_DIN_pipe(4), RX_FIFO_DIN_pipe(3) => 
        RX_FIFO_DIN_pipe(3), RX_FIFO_DIN_pipe(2) => 
        RX_FIFO_DIN_pipe(2), RX_FIFO_DIN_pipe(1) => 
        RX_FIFO_DIN_pipe(1), RX_FIFO_DIN_pipe(0) => 
        RX_FIFO_DIN_pipe(0), fifo_MEMRADDR(10) => 
        fifo_MEMRADDR(10), fifo_MEMRADDR(9) => fifo_MEMRADDR(9), 
        fifo_MEMRADDR(8) => fifo_MEMRADDR(8), fifo_MEMRADDR(7)
         => fifo_MEMRADDR(7), fifo_MEMRADDR(6) => 
        fifo_MEMRADDR(6), fifo_MEMRADDR(5) => fifo_MEMRADDR(5), 
        fifo_MEMRADDR(4) => fifo_MEMRADDR(4), fifo_MEMRADDR(3)
         => fifo_MEMRADDR(3), fifo_MEMRADDR(2) => 
        fifo_MEMRADDR(2), fifo_MEMRADDR(1) => fifo_MEMRADDR(1), 
        fifo_MEMRADDR(0) => fifo_MEMRADDR(0), RDATA_int(8) => 
        RDATA_int(8), RDATA_int(7) => RDATA_int(7), RDATA_int(6)
         => RDATA_int(6), RDATA_int(5) => RDATA_int(5), 
        RDATA_int(4) => RDATA_int(4), RDATA_int(3) => 
        RDATA_int(3), RDATA_int(2) => RDATA_int(2), RDATA_int(1)
         => RDATA_int(1), RDATA_int(0) => RDATA_int(0), 
        fifo_MEMWE => fifo_MEMWE, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, N_1007_i => N_1007_i, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_0 is

    port( wptr_bin_sync  : inout std_logic_vector(11 downto 0) := (others => 'Z');
          wptr_gray_sync : in    std_logic_vector(10 downto 0)
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_0;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    \bin_out_xhdl1_0_a2[1]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(3), B => wptr_gray_sync(1), C
         => wptr_bin_sync(4), D => wptr_gray_sync(2), Y => 
        wptr_bin_sync(1));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \bin_out_xhdl1_0_a2[5]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(7), B => wptr_gray_sync(6), C
         => wptr_gray_sync(5), D => wptr_bin_sync(8), Y => 
        wptr_bin_sync(5));
    
    \bin_out_xhdl1_0_a2[2]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(4), B => wptr_gray_sync(3), C
         => wptr_gray_sync(2), D => wptr_bin_sync(5), Y => 
        wptr_bin_sync(2));
    
    \bin_out_xhdl1_0_a2[0]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(2), B => wptr_bin_sync(3), C
         => wptr_gray_sync(0), D => wptr_gray_sync(1), Y => 
        wptr_bin_sync(0));
    
    \bin_out_xhdl1_i_o2[9]\ : CFG3
      generic map(INIT => x"96")

      port map(A => wptr_gray_sync(10), B => wptr_gray_sync(9), C
         => wptr_bin_sync(11), Y => wptr_bin_sync(9));
    
    \bin_out_xhdl1_i_o2[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => wptr_bin_sync(11), B => wptr_gray_sync(10), Y
         => wptr_bin_sync(10));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \bin_out_xhdl1_0_a2[6]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(8), B => wptr_gray_sync(7), C
         => wptr_gray_sync(6), D => wptr_bin_sync(9), Y => 
        wptr_bin_sync(6));
    
    \bin_out_xhdl1_0_a2[4]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(6), B => wptr_gray_sync(5), C
         => wptr_gray_sync(4), D => wptr_bin_sync(7), Y => 
        wptr_bin_sync(4));
    
    \bin_out_xhdl1_0_a2[8]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(10), B => wptr_gray_sync(9), C
         => wptr_gray_sync(8), D => wptr_bin_sync(11), Y => 
        wptr_bin_sync(8));
    
    \bin_out_xhdl1_0_a2[7]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(9), B => wptr_gray_sync(8), C
         => wptr_gray_sync(7), D => wptr_bin_sync(10), Y => 
        wptr_bin_sync(7));
    
    \bin_out_xhdl1_0_a2[3]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(5), B => wptr_gray_sync(4), C
         => wptr_gray_sync(3), D => wptr_bin_sync(6), Y => 
        wptr_bin_sync(3));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync is

    port( wptr_gray                 : in    std_logic_vector(11 downto 0);
          wptr_gray_sync            : out   std_logic_vector(10 downto 0);
          wptr_bin_sync_0           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          irx_fifo_rst_i            : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \sync_int[10]_net_1\, VCC_net_1, GND_net_1, 
        \sync_int[11]_net_1\, \sync_int[0]_net_1\, 
        \sync_int[1]_net_1\, \sync_int[2]_net_1\, 
        \sync_int[3]_net_1\, \sync_int[4]_net_1\, 
        \sync_int[5]_net_1\, \sync_int[6]_net_1\, 
        \sync_int[7]_net_1\, \sync_int[8]_net_1\, 
        \sync_int[9]_net_1\ : std_logic;

begin 


    \sync_int[9]\ : SLE
      port map(D => wptr_gray(9), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[9]_net_1\);
    
    \sync_int[4]\ : SLE
      port map(D => wptr_gray(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[4]_net_1\);
    
    \sync_out_xhdl1[10]\ : SLE
      port map(D => \sync_int[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(10));
    
    \sync_int[1]\ : SLE
      port map(D => wptr_gray(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[1]_net_1\);
    
    \sync_int[11]\ : SLE
      port map(D => wptr_gray(11), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[11]_net_1\);
    
    \sync_out_xhdl1[6]\ : SLE
      port map(D => \sync_int[6]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(6));
    
    \sync_out_xhdl1[3]\ : SLE
      port map(D => \sync_int[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(3));
    
    \sync_int[6]\ : SLE
      port map(D => wptr_gray(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[6]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \sync_out_xhdl1[11]\ : SLE
      port map(D => \sync_int[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_bin_sync_0);
    
    \sync_int[3]\ : SLE
      port map(D => wptr_gray(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[3]_net_1\);
    
    \sync_out_xhdl1[4]\ : SLE
      port map(D => \sync_int[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(4));
    
    \sync_int[0]\ : SLE
      port map(D => wptr_gray(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[0]_net_1\);
    
    \sync_out_xhdl1[1]\ : SLE
      port map(D => \sync_int[1]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(1));
    
    \sync_int[5]\ : SLE
      port map(D => wptr_gray(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[5]_net_1\);
    
    \sync_int[2]\ : SLE
      port map(D => wptr_gray(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[2]_net_1\);
    
    \sync_out_xhdl1[9]\ : SLE
      port map(D => \sync_int[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(9));
    
    \sync_out_xhdl1[2]\ : SLE
      port map(D => \sync_int[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(2));
    
    \sync_int[8]\ : SLE
      port map(D => wptr_gray(8), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[8]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sync_out_xhdl1[7]\ : SLE
      port map(D => \sync_int[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(7));
    
    \sync_out_xhdl1[5]\ : SLE
      port map(D => \sync_int[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(5));
    
    \sync_out_xhdl1[0]\ : SLE
      port map(D => \sync_int[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(0));
    
    \sync_out_xhdl1[8]\ : SLE
      port map(D => \sync_int[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(8));
    
    \sync_int[7]\ : SLE
      port map(D => wptr_gray(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[7]_net_1\);
    
    \sync_int[10]\ : SLE
      port map(D => wptr_gray(10), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0 is

    port( rptr_gray           : in    std_logic_vector(11 downto 0);
          rptr_gray_sync      : out   std_logic_vector(10 downto 0);
          rptr_bin_sync_0     : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          irx_fifo_rst_i      : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \sync_int[4]_net_1\, GND_net_1, 
        \sync_int[5]_net_1\, \sync_int[6]_net_1\, 
        \sync_int[7]_net_1\, \sync_int[8]_net_1\, 
        \sync_int[9]_net_1\, \sync_int[10]_net_1\, 
        \sync_int[11]_net_1\, \sync_int[1]_net_1\, 
        \sync_int[2]_net_1\, \sync_int[3]_net_1\, 
        \sync_int[0]_net_1\ : std_logic;

begin 


    \sync_int[9]\ : SLE
      port map(D => rptr_gray(9), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[9]_net_1\);
    
    \sync_int[4]\ : SLE
      port map(D => rptr_gray(4), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[4]_net_1\);
    
    \sync_out_xhdl1[10]\ : SLE
      port map(D => \sync_int[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(10));
    
    \sync_int[1]\ : SLE
      port map(D => rptr_gray(1), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[1]_net_1\);
    
    \sync_int[11]\ : SLE
      port map(D => rptr_gray(11), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[11]_net_1\);
    
    \sync_out_xhdl1[6]\ : SLE
      port map(D => \sync_int[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(6));
    
    \sync_out_xhdl1[3]\ : SLE
      port map(D => \sync_int[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(3));
    
    \sync_int[6]\ : SLE
      port map(D => rptr_gray(6), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[6]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \sync_out_xhdl1[11]\ : SLE
      port map(D => \sync_int[11]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_bin_sync_0);
    
    \sync_int[3]\ : SLE
      port map(D => rptr_gray(3), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[3]_net_1\);
    
    \sync_out_xhdl1[4]\ : SLE
      port map(D => \sync_int[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(4));
    
    \sync_int[0]\ : SLE
      port map(D => rptr_gray(0), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[0]_net_1\);
    
    \sync_out_xhdl1[1]\ : SLE
      port map(D => \sync_int[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(1));
    
    \sync_int[5]\ : SLE
      port map(D => rptr_gray(5), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[5]_net_1\);
    
    \sync_int[2]\ : SLE
      port map(D => rptr_gray(2), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[2]_net_1\);
    
    \sync_out_xhdl1[9]\ : SLE
      port map(D => \sync_int[9]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(9));
    
    \sync_out_xhdl1[2]\ : SLE
      port map(D => \sync_int[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(2));
    
    \sync_int[8]\ : SLE
      port map(D => rptr_gray(8), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[8]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sync_out_xhdl1[7]\ : SLE
      port map(D => \sync_int[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(7));
    
    \sync_out_xhdl1[5]\ : SLE
      port map(D => \sync_int[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(5));
    
    \sync_out_xhdl1[0]\ : SLE
      port map(D => \sync_int[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(0));
    
    \sync_out_xhdl1[8]\ : SLE
      port map(D => \sync_int[8]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(8));
    
    \sync_int[7]\ : SLE
      port map(D => rptr_gray(7), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[7]_net_1\);
    
    \sync_int[10]\ : SLE
      port map(D => rptr_gray(10), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3 is

    port( rptr_bin_sync  : inout std_logic_vector(11 downto 0) := (others => 'Z');
          rptr_gray_sync : in    std_logic_vector(10 downto 0)
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3 is 

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    \bin_out_xhdl1_0_a2[1]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(1), B => rptr_gray_sync(2), C
         => rptr_bin_sync(3), Y => rptr_bin_sync(1));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \bin_out_xhdl1_0_a2[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(6), B => rptr_gray_sync(5), Y
         => rptr_bin_sync(5));
    
    \bin_out_xhdl1_0_a2[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(3), B => rptr_gray_sync(2), Y
         => rptr_bin_sync(2));
    
    \bin_out_xhdl1_0_a2[0]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(1), B => rptr_gray_sync(0), C
         => rptr_bin_sync(3), D => rptr_gray_sync(2), Y => 
        rptr_bin_sync(0));
    
    \bin_out_xhdl1_i_o2[9]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(9), B => rptr_gray_sync(10), C
         => rptr_bin_sync(11), Y => rptr_bin_sync(9));
    
    \bin_out_xhdl1_i_o2[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(11), B => rptr_gray_sync(10), Y
         => rptr_bin_sync(10));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \bin_out_xhdl1_0_a2[6]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(6), B => rptr_gray_sync(7), C
         => rptr_gray_sync(8), D => rptr_bin_sync(9), Y => 
        rptr_bin_sync(6));
    
    \bin_out_xhdl1_0_a2[4]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(4), B => rptr_gray_sync(5), C
         => rptr_bin_sync(6), Y => rptr_bin_sync(4));
    
    \bin_out_xhdl1_0_a2[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(9), B => rptr_gray_sync(8), Y
         => rptr_bin_sync(8));
    
    \bin_out_xhdl1_0_a2[7]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(8), B => rptr_bin_sync(9), C
         => rptr_gray_sync(7), Y => rptr_bin_sync(7));
    
    \bin_out_xhdl1_0_a2[3]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(5), B => rptr_bin_sync(6), C
         => rptr_gray_sync(3), D => rptr_gray_sync(4), Y => 
        rptr_bin_sync(3));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3 is

    port( ReadFIFO_Write_Ptr        : in    std_logic_vector(1 downto 0);
          fifo_MEMWADDR             : out   std_logic_vector(10 downto 0);
          fifo_MEMRADDR             : out   std_logic_vector(10 downto 0);
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          N_153_i_i                 : out   std_logic;
          N_89_i                    : out   std_logic;
          REN_d1                    : in    std_logic;
          N_1004                    : in    std_logic;
          tx_col_detect_en          : in    std_logic;
          RX_InProcess_d1           : in    std_logic;
          sampler_clk1x_en          : in    std_logic;
          iRX_FIFO_wr_en            : in    std_logic;
          N_1466                    : out   std_logic;
          N_1007_i                  : out   std_logic;
          fifo_MEMWE                : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          irx_fifo_rst_i            : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3 is 

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_0
    port( wptr_bin_sync  : inout   std_logic_vector(11 downto 0);
          wptr_gray_sync : in    std_logic_vector(10 downto 0) := (others => 'U')
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync
    port( wptr_gray                 : in    std_logic_vector(11 downto 0) := (others => 'U');
          wptr_gray_sync            : out   std_logic_vector(10 downto 0);
          wptr_bin_sync_0           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          irx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0
    port( rptr_gray           : in    std_logic_vector(11 downto 0) := (others => 'U');
          rptr_gray_sync      : out   std_logic_vector(10 downto 0);
          rptr_bin_sync_0     : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          irx_fifo_rst_i      : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3
    port( rptr_bin_sync  : inout   std_logic_vector(11 downto 0);
          rptr_gray_sync : in    std_logic_vector(10 downto 0) := (others => 'U')
        );
  end component;

    signal \rptr[0]_net_1\, \rptr_s[0]\, \fifo_MEMRADDR[0]\, 
        \memraddr_r_s[0]\, \wptr[0]_net_1\, \wptr_s[0]\, 
        \wptr_gray[10]_net_1\, VCC_net_1, \wptr_gray_1[10]_net_1\, 
        GND_net_1, \wptr_gray[11]_net_1\, \wptr[11]_net_1\, 
        \rptr_gray[0]_net_1\, \rptr_gray_1[0]_net_1\, 
        \rptr_gray[1]_net_1\, \rptr_gray_1[1]_net_1\, 
        \rptr_gray[2]_net_1\, \rptr_gray_1[2]_net_1\, 
        \rptr_gray[3]_net_1\, \rptr_gray_1[3]_net_1\, 
        \rptr_gray[4]_net_1\, \rptr_gray_1[4]_net_1\, 
        \rptr_gray[5]_net_1\, \rptr_gray_1[5]_net_1\, 
        \rptr_gray[6]_net_1\, \rptr_gray_1[6]_net_1\, 
        \rptr_gray[7]_net_1\, \rptr_gray_1[7]_net_1\, 
        \rptr_gray[8]_net_1\, \rptr_gray_1[8]_net_1\, 
        \rptr_gray[9]_net_1\, \rptr_gray_1[9]_net_1\, 
        \rptr_gray[10]_net_1\, \rptr_gray_1[10]_net_1\, 
        \rptr_gray[11]_net_1\, \rptr[11]_net_1\, 
        \wptr_bin_sync2[7]_net_1\, \wptr_bin_sync[7]\, 
        \wptr_bin_sync2[8]_net_1\, \wptr_bin_sync[8]\, 
        \wptr_bin_sync2[9]_net_1\, \wptr_bin_sync[9]\, 
        \wptr_bin_sync2[10]_net_1\, \wptr_bin_sync[10]\, 
        \wptr_bin_sync2[11]_net_1\, \wptr_bin_sync[11]\, 
        \wptr_gray[0]_net_1\, \wptr_gray_1[0]_net_1\, 
        \wptr_gray[1]_net_1\, \wptr_gray_1[1]_net_1\, 
        \wptr_gray[2]_net_1\, \wptr_gray_1[2]_net_1\, 
        \wptr_gray[3]_net_1\, \wptr_gray_1[3]_net_1\, 
        \wptr_gray[4]_net_1\, \wptr_gray_1[4]_net_1\, 
        \wptr_gray[5]_net_1\, \wptr_gray_1[5]_net_1\, 
        \wptr_gray[6]_net_1\, \wptr_gray_1[6]_net_1\, 
        \wptr_gray[7]_net_1\, \wptr_gray_1[7]_net_1\, 
        \wptr_gray[8]_net_1\, \wptr_gray_1[8]_net_1\, 
        \wptr_gray[9]_net_1\, \wptr_gray_1[9]_net_1\, rdiff_bus, 
        \wptr_bin_sync[0]\, \wptr_bin_sync2[1]_net_1\, 
        \wptr_bin_sync[1]\, \wptr_bin_sync2[2]_net_1\, 
        \wptr_bin_sync[2]\, \wptr_bin_sync2[3]_net_1\, 
        \wptr_bin_sync[3]\, \wptr_bin_sync2[4]_net_1\, 
        \wptr_bin_sync[4]\, \wptr_bin_sync2[5]_net_1\, 
        \wptr_bin_sync[5]\, \wptr_bin_sync2[6]_net_1\, 
        \wptr_bin_sync[6]\, \rptr_bin_sync2[7]_net_1\, 
        \rptr_bin_sync[7]\, \rptr_bin_sync2[8]_net_1\, 
        \rptr_bin_sync[8]\, \rptr_bin_sync2[9]_net_1\, 
        \rptr_bin_sync[9]\, \rptr_bin_sync2[10]_net_1\, 
        \rptr_bin_sync[10]\, \rptr_bin_sync2[11]_net_1\, 
        \rptr_bin_sync[11]\, un1_we_p, \rptr_bin_sync2[0]_net_1\, 
        \rptr_bin_sync[0]\, \rptr_bin_sync2[1]_net_1\, 
        \rptr_bin_sync[1]\, \rptr_bin_sync2[2]_net_1\, 
        \rptr_bin_sync[2]\, \rptr_bin_sync2[3]_net_1\, 
        \rptr_bin_sync[3]\, \rptr_bin_sync2[4]_net_1\, 
        \rptr_bin_sync[4]\, \rptr_bin_sync2[5]_net_1\, 
        \rptr_bin_sync[5]\, \rptr_bin_sync2[6]_net_1\, 
        \rptr_bin_sync[6]\, \iRX_FIFO_Full_0\, fulli, 
        un2_re_p_i_i_a3, \iRX_FIFO_Empty_0\, empty_r_3, 
        \fifo_MEMWE\, \wptr[1]_net_1\, \wptr_s[1]\, 
        \wptr[2]_net_1\, \wptr_s[2]\, \wptr[3]_net_1\, 
        \wptr_s[3]\, \wptr[4]_net_1\, \wptr_s[4]\, 
        \wptr[5]_net_1\, \wptr_s[5]\, \wptr[6]_net_1\, 
        \wptr_s[6]\, \wptr[7]_net_1\, \wptr_s[7]\, 
        \wptr[8]_net_1\, \wptr_s[8]\, \wptr[9]_net_1\, 
        \wptr_s[9]\, \wptr[10]_net_1\, \wptr_s[10]\, 
        \wptr_s[11]_net_1\, \N_1007_i\, \fifo_MEMRADDR[1]\, 
        \memraddr_r_s[1]\, \fifo_MEMRADDR[2]\, \memraddr_r_s[2]\, 
        \fifo_MEMRADDR[3]\, \memraddr_r_s[3]\, \fifo_MEMRADDR[4]\, 
        \memraddr_r_s[4]\, \fifo_MEMRADDR[5]\, \memraddr_r_s[5]\, 
        \fifo_MEMRADDR[6]\, \memraddr_r_s[6]\, \fifo_MEMRADDR[7]\, 
        \memraddr_r_s[7]\, \fifo_MEMRADDR[8]\, \memraddr_r_s[8]\, 
        \fifo_MEMRADDR[9]\, \memraddr_r_s[9]\, 
        \fifo_MEMRADDR[10]\, \memraddr_r_s[10]_net_1\, 
        \fifo_MEMWADDR[0]\, \memwaddr_r_s[0]\, N_248, 
        \fifo_MEMWADDR[1]\, \memwaddr_r_s[1]\, \fifo_MEMWADDR[2]\, 
        \memwaddr_r_s[2]\, \fifo_MEMWADDR[3]\, \memwaddr_r_s[3]\, 
        \fifo_MEMWADDR[4]\, \memwaddr_r_s[4]\, \fifo_MEMWADDR[5]\, 
        \memwaddr_r_s[5]\, \fifo_MEMWADDR[6]\, \memwaddr_r_s[6]\, 
        \fifo_MEMWADDR[7]\, \memwaddr_r_s[7]\, \fifo_MEMWADDR[8]\, 
        \memwaddr_r_s[8]\, \fifo_MEMWADDR[9]\, \memwaddr_r_s[9]\, 
        \fifo_MEMWADDR[10]\, \memwaddr_r_s[10]_net_1\, 
        \rptr[1]_net_1\, \rptr_s[1]\, \rptr[2]_net_1\, 
        \rptr_s[2]\, \rptr[3]_net_1\, \rptr_s[3]\, 
        \rptr[4]_net_1\, \rptr_s[4]\, \rptr[5]_net_1\, 
        \rptr_s[5]\, \rptr[6]_net_1\, \rptr_s[6]\, 
        \rptr[7]_net_1\, \rptr_s[7]\, \rptr[8]_net_1\, 
        \rptr_s[8]\, \rptr[9]_net_1\, \rptr_s[9]\, 
        \rptr[10]_net_1\, \rptr_s[10]\, \rptr_s[11]_net_1\, 
        memwaddr_r_cry_cy, \memwaddr_r_cry[0]_net_1\, 
        \memwaddr_r_cry[1]_net_1\, \memwaddr_r_cry[2]_net_1\, 
        \memwaddr_r_cry[3]_net_1\, \memwaddr_r_cry[4]_net_1\, 
        \memwaddr_r_cry[5]_net_1\, \memwaddr_r_cry[6]_net_1\, 
        \memwaddr_r_cry[7]_net_1\, \memwaddr_r_cry[8]_net_1\, 
        \memwaddr_r_cry[9]_net_1\, \rdiff_bus_cry_0\, 
        rdiff_bus_cry_0_Y_0, \rdiff_bus_cry_1\, \rdiff_bus[1]\, 
        \rdiff_bus_cry_2\, \rdiff_bus[2]\, \rdiff_bus_cry_3\, 
        \rdiff_bus[3]\, \rdiff_bus_cry_4\, \rdiff_bus[4]\, 
        \rdiff_bus_cry_5\, \rdiff_bus[5]\, \rdiff_bus_cry_6\, 
        \rdiff_bus[6]\, \rdiff_bus_cry_7\, \rdiff_bus[7]\, 
        \rdiff_bus_cry_8\, \rdiff_bus[8]\, \rdiff_bus_cry_9\, 
        \rdiff_bus[9]\, \rdiff_bus[11]\, \rdiff_bus_cry_10\, 
        \rdiff_bus[10]\, \wdiff_bus_cry_0\, wdiff_bus_cry_0_Y_0, 
        \wdiff_bus_cry_1\, \wdiff_bus[1]\, \wdiff_bus_cry_2\, 
        \wdiff_bus[2]\, \wdiff_bus_cry_3\, \wdiff_bus[3]\, 
        \wdiff_bus_cry_4\, \wdiff_bus[4]\, \wdiff_bus_cry_5\, 
        \wdiff_bus[5]\, \wdiff_bus_cry_6\, \wdiff_bus[6]\, 
        \wdiff_bus_cry_7\, \wdiff_bus[7]\, \wdiff_bus_cry_8\, 
        \wdiff_bus[8]\, \wdiff_bus_cry_9\, \wdiff_bus[9]\, 
        \wdiff_bus[11]\, \wdiff_bus_cry_10\, \wdiff_bus[10]\, 
        rptr_s_383_FCO, \rptr_cry[1]_net_1\, \rptr_cry[2]_net_1\, 
        \rptr_cry[3]_net_1\, \rptr_cry[4]_net_1\, 
        \rptr_cry[5]_net_1\, \rptr_cry[6]_net_1\, 
        \rptr_cry[7]_net_1\, \rptr_cry[8]_net_1\, 
        \rptr_cry[9]_net_1\, \rptr_cry[10]_net_1\, 
        memraddr_r_s_384_FCO, \memraddr_r_cry[1]_net_1\, 
        \memraddr_r_cry[2]_net_1\, \memraddr_r_cry[3]_net_1\, 
        \memraddr_r_cry[4]_net_1\, \memraddr_r_cry[5]_net_1\, 
        \memraddr_r_cry[6]_net_1\, \memraddr_r_cry[7]_net_1\, 
        \memraddr_r_cry[8]_net_1\, \memraddr_r_cry[9]_net_1\, 
        wptr_s_385_FCO, \wptr_cry[1]_net_1\, \wptr_cry[2]_net_1\, 
        \wptr_cry[3]_net_1\, \wptr_cry[4]_net_1\, 
        \wptr_cry[5]_net_1\, \wptr_cry[6]_net_1\, 
        \wptr_cry[7]_net_1\, \wptr_cry[8]_net_1\, 
        \wptr_cry[9]_net_1\, \wptr_cry[10]_net_1\, \N_1466\, 
        empty_r_3_0_a2_1, \fulli_0_a2_7\, \fulli_0_a2_6\, 
        empty_r_3_0_a2_7, empty_r_3_0_a2_9, \fulli_0_a2_8\, 
        empty_r_3_0_a2_5, \wptr_gray_sync[0]\, 
        \wptr_gray_sync[1]\, \wptr_gray_sync[2]\, 
        \wptr_gray_sync[3]\, \wptr_gray_sync[4]\, 
        \wptr_gray_sync[5]\, \wptr_gray_sync[6]\, 
        \wptr_gray_sync[7]\, \wptr_gray_sync[8]\, 
        \wptr_gray_sync[9]\, \wptr_gray_sync[10]\, 
        \rptr_gray_sync[0]\, \rptr_gray_sync[1]\, 
        \rptr_gray_sync[2]\, \rptr_gray_sync[3]\, 
        \rptr_gray_sync[4]\, \rptr_gray_sync[5]\, 
        \rptr_gray_sync[6]\, \rptr_gray_sync[7]\, 
        \rptr_gray_sync[8]\, \rptr_gray_sync[9]\, 
        \rptr_gray_sync[10]\ : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_0
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_0(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3(DEF_ARCH);
begin 

    fifo_MEMWADDR(10) <= \fifo_MEMWADDR[10]\;
    fifo_MEMWADDR(9) <= \fifo_MEMWADDR[9]\;
    fifo_MEMWADDR(8) <= \fifo_MEMWADDR[8]\;
    fifo_MEMWADDR(7) <= \fifo_MEMWADDR[7]\;
    fifo_MEMWADDR(6) <= \fifo_MEMWADDR[6]\;
    fifo_MEMWADDR(5) <= \fifo_MEMWADDR[5]\;
    fifo_MEMWADDR(4) <= \fifo_MEMWADDR[4]\;
    fifo_MEMWADDR(3) <= \fifo_MEMWADDR[3]\;
    fifo_MEMWADDR(2) <= \fifo_MEMWADDR[2]\;
    fifo_MEMWADDR(1) <= \fifo_MEMWADDR[1]\;
    fifo_MEMWADDR(0) <= \fifo_MEMWADDR[0]\;
    fifo_MEMRADDR(10) <= \fifo_MEMRADDR[10]\;
    fifo_MEMRADDR(9) <= \fifo_MEMRADDR[9]\;
    fifo_MEMRADDR(8) <= \fifo_MEMRADDR[8]\;
    fifo_MEMRADDR(7) <= \fifo_MEMRADDR[7]\;
    fifo_MEMRADDR(6) <= \fifo_MEMRADDR[6]\;
    fifo_MEMRADDR(5) <= \fifo_MEMRADDR[5]\;
    fifo_MEMRADDR(4) <= \fifo_MEMRADDR[4]\;
    fifo_MEMRADDR(3) <= \fifo_MEMRADDR[3]\;
    fifo_MEMRADDR(2) <= \fifo_MEMRADDR[2]\;
    fifo_MEMRADDR(1) <= \fifo_MEMRADDR[1]\;
    fifo_MEMRADDR(0) <= \fifo_MEMRADDR[0]\;
    iRX_FIFO_Empty_0 <= \iRX_FIFO_Empty_0\;
    iRX_FIFO_Full_0 <= \iRX_FIFO_Full_0\;
    N_1466 <= \N_1466\;
    N_1007_i <= \N_1007_i\;
    fifo_MEMWE <= \fifo_MEMWE\;

    \rptr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[4]_net_1\, S
         => \rptr_s[5]\, Y => OPEN, FCO => \rptr_cry[5]_net_1\);
    
    empty_r_RNIUREJ1 : CFG3
      generic map(INIT => x"A6")

      port map(A => REN_d1, B => N_1004, C => \iRX_FIFO_Empty_0\, 
        Y => N_153_i_i);
    
    wdiff_bus_cry_8 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[8]_net_1\, B => 
        \rptr_bin_sync2[8]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_7\, S => \wdiff_bus[8]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_8\);
    
    \wptr_gray[4]\ : SLE
      port map(D => \wptr_gray_1[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[4]_net_1\);
    
    \rptr_gray_1[3]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[3]_net_1\, B => \rptr[4]_net_1\, Y => 
        \rptr_gray_1[3]_net_1\);
    
    \rptr_bin_sync2[6]\ : SLE
      port map(D => \rptr_bin_sync[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[6]_net_1\);
    
    fulli_0_a2_0_0_a2 : CFG3
      generic map(INIT => x"04")

      port map(A => ReadFIFO_Write_Ptr(0), B => \N_1466\, C => 
        ReadFIFO_Write_Ptr(1), Y => N_248);
    
    \rptr[1]\ : SLE
      port map(D => \rptr_s[1]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1007_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[1]_net_1\);
    
    \wptr_gray_1[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[9]_net_1\, B => \wptr[10]_net_1\, Y => 
        \wptr_gray_1[9]_net_1\);
    
    \rptr_gray_1[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[5]_net_1\, B => \rptr[6]_net_1\, Y => 
        \rptr_gray_1[5]_net_1\);
    
    \rptr_gray[9]\ : SLE
      port map(D => \rptr_gray_1[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[9]_net_1\);
    
    \rptr_gray[8]\ : SLE
      port map(D => \rptr_gray_1[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[8]_net_1\);
    
    \rptr_gray_1[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[2]_net_1\, B => \rptr[3]_net_1\, Y => 
        \rptr_gray_1[2]_net_1\);
    
    \rptr_bin_sync2[7]\ : SLE
      port map(D => \rptr_bin_sync[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[7]_net_1\);
    
    \memwaddr_r[1]\ : SLE
      port map(D => \memwaddr_r_s[1]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_248, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[1]\);
    
    empty_r_RNI0SB51 : CFG2
      generic map(INIT => x"2")

      port map(A => N_1004, B => \iRX_FIFO_Empty_0\, Y => 
        \N_1007_i\);
    
    \memwaddr_r_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[5]_net_1\, S => \memwaddr_r_s[6]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[6]_net_1\);
    
    \memwaddr_r_s[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[9]_net_1\, S => \memwaddr_r_s[10]_net_1\, 
        Y => OPEN, FCO => OPEN);
    
    \wptr_gray_1[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[7]_net_1\, B => \wptr[8]_net_1\, Y => 
        \wptr_gray_1[7]_net_1\);
    
    \memraddr_r[0]\ : SLE
      port map(D => \memraddr_r_s[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1007_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[0]\);
    
    \wptr[0]\ : SLE
      port map(D => \wptr_s[0]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[0]_net_1\);
    
    \rptr_bin_sync2[8]\ : SLE
      port map(D => \rptr_bin_sync[8]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[8]_net_1\);
    
    \rptr_gray_1[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[1]_net_1\, B => \rptr[2]_net_1\, Y => 
        \rptr_gray_1[1]_net_1\);
    
    \rptr_gray[10]\ : SLE
      port map(D => \rptr_gray_1[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[10]_net_1\);
    
    \wptr_gray_1[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[0]_net_1\, B => \wptr[1]_net_1\, Y => 
        \wptr_gray_1[0]_net_1\);
    
    wdiff_bus_cry_9 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[9]_net_1\, B => 
        \rptr_bin_sync2[9]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_8\, S => \wdiff_bus[9]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_9\);
    
    \rptr[5]\ : SLE
      port map(D => \rptr_s[5]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1007_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[5]_net_1\);
    
    \rptr_gray[3]\ : SLE
      port map(D => \rptr_gray_1[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[3]_net_1\);
    
    \rptr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[5]_net_1\, S
         => \rptr_s[6]\, Y => OPEN, FCO => \rptr_cry[6]_net_1\);
    
    \memwaddr_r_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[1]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[0]_net_1\, S => \memwaddr_r_s[1]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[1]_net_1\);
    
    fulli_0_a2_6 : CFG4
      generic map(INIT => x"8000")

      port map(A => \wdiff_bus[2]\, B => \wdiff_bus[3]\, C => 
        \wdiff_bus[5]\, D => \wdiff_bus[4]\, Y => \fulli_0_a2_6\);
    
    \wptr_gray[3]\ : SLE
      port map(D => \wptr_gray_1[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[3]_net_1\);
    
    \rptr_gray_1[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[11]_net_1\, B => \rptr[10]_net_1\, Y
         => \rptr_gray_1[10]_net_1\);
    
    wdiff_bus_s_11 : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \rptr_bin_sync2[11]_net_1\, C
         => \wptr[11]_net_1\, D => GND_net_1, FCI => 
        \wdiff_bus_cry_10\, S => \wdiff_bus[11]\, Y => OPEN, FCO
         => OPEN);
    
    \rptr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[7]_net_1\, S
         => \rptr_s[8]\, Y => OPEN, FCO => \rptr_cry[8]_net_1\);
    
    \rptr[7]\ : SLE
      port map(D => \rptr_s[7]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1007_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[7]_net_1\);
    
    rdiff_bus_cry_4 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[4]_net_1\, B => 
        \rptr[4]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_3\, S => \rdiff_bus[4]\, Y => OPEN, FCO
         => \rdiff_bus_cry_4\);
    
    \rptr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[9]_net_1\, S
         => \rptr_s[10]\, Y => OPEN, FCO => \rptr_cry[10]_net_1\);
    
    \rptr_bin_sync2[0]\ : SLE
      port map(D => \rptr_bin_sync[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[0]_net_1\);
    
    \L1.empty_r_3_0_a2_7\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \rdiff_bus[5]\, B => \rdiff_bus[6]\, C => 
        \rdiff_bus[7]\, D => \rdiff_bus[8]\, Y => 
        empty_r_3_0_a2_7);
    
    \wptr[11]\ : SLE
      port map(D => \wptr_s[11]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \wptr[11]_net_1\);
    
    rdiff_bus_cry_1 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[1]_net_1\, B => 
        \rptr[1]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_0\, S => \rdiff_bus[1]\, Y => OPEN, FCO
         => \rdiff_bus_cry_1\);
    
    rptr_s_383 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => rptr_s_383_FCO);
    
    \memraddr_r[1]\ : SLE
      port map(D => \memraddr_r_s[1]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1007_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[1]\);
    
    \L1.empty_r_3_0_a2_9\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \rdiff_bus[1]\, B => \rdiff_bus[2]\, C => 
        empty_r_3_0_a2_7, D => empty_r_3_0_a2_1, Y => 
        empty_r_3_0_a2_9);
    
    \rptr_bin_sync2[2]\ : SLE
      port map(D => \rptr_bin_sync[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[2]_net_1\);
    
    rdiff_bus_cry_6 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[6]_net_1\, B => 
        \rptr[6]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_5\, S => \rdiff_bus[6]\, Y => OPEN, FCO
         => \rdiff_bus_cry_6\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \memwaddr_r_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[3]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[2]_net_1\, S => \memwaddr_r_s[3]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[3]_net_1\);
    
    \rptr_gray[1]\ : SLE
      port map(D => \rptr_gray_1[1]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[1]_net_1\);
    
    \memwaddr_r[7]\ : SLE
      port map(D => \memwaddr_r_s[7]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_248, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[7]\);
    
    \memraddr_r_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[2]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[1]_net_1\, S => \memraddr_r_s[2]\, Y => 
        OPEN, FCO => \memraddr_r_cry[2]_net_1\);
    
    \wptr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[3]_net_1\, S
         => \wptr_s[4]\, Y => OPEN, FCO => \wptr_cry[4]_net_1\);
    
    \memraddr_r_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[8]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[7]_net_1\, S => \memraddr_r_s[8]\, Y => 
        OPEN, FCO => \memraddr_r_cry[8]_net_1\);
    
    \wptr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[9]_net_1\, S
         => \wptr_s[10]\, Y => OPEN, FCO => \wptr_cry[10]_net_1\);
    
    wdiff_bus_cry_5 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[5]_net_1\, B => 
        \rptr_bin_sync2[5]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_4\, S => \wdiff_bus[5]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_5\);
    
    \memwaddr_r[4]\ : SLE
      port map(D => \memwaddr_r_s[4]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_248, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[4]\);
    
    \wptr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[1]_net_1\, S
         => \wptr_s[2]\, Y => OPEN, FCO => \wptr_cry[2]_net_1\);
    
    wdiff_bus_cry_0 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[0]_net_1\, B => 
        \rptr_bin_sync2[0]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => VCC_net_1, S => OPEN, Y => wdiff_bus_cry_0_Y_0, 
        FCO => \wdiff_bus_cry_0\);
    
    \wptr[1]\ : SLE
      port map(D => \wptr_s[1]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[1]_net_1\);
    
    \rptr_bin_sync2[4]\ : SLE
      port map(D => \rptr_bin_sync[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[4]_net_1\);
    
    \wptr_bin_sync2[6]\ : SLE
      port map(D => \wptr_bin_sync[6]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[6]_net_1\);
    
    \memwaddr_r_cry_cy[0]\ : ARI1
      generic map(INIT => x"45500")

      port map(A => VCC_net_1, B => \iRX_FIFO_Full_0\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => memwaddr_r_cry_cy);
    
    \rptr[3]\ : SLE
      port map(D => \rptr_s[3]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1007_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[3]_net_1\);
    
    \wptr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[2]_net_1\, S
         => \wptr_s[3]\, Y => OPEN, FCO => \wptr_cry[3]_net_1\);
    
    \memwaddr_r_cry[0]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[0]\, C => 
        GND_net_1, D => GND_net_1, FCI => memwaddr_r_cry_cy, S
         => \memwaddr_r_s[0]\, Y => OPEN, FCO => 
        \memwaddr_r_cry[0]_net_1\);
    
    \rptr[6]\ : SLE
      port map(D => \rptr_s[6]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1007_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[6]_net_1\);
    
    rdiff_bus_cry_8 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[8]_net_1\, B => 
        \rptr[8]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_7\, S => \rdiff_bus[8]\, Y => OPEN, FCO
         => \rdiff_bus_cry_8\);
    
    \wptr_gray[10]\ : SLE
      port map(D => \wptr_gray_1[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[10]_net_1\);
    
    rdiff_bus_cry_7 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[7]_net_1\, B => 
        \rptr[7]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_6\, S => \rdiff_bus[7]\, Y => OPEN, FCO
         => \rdiff_bus_cry_7\);
    
    \wptr_bin_sync2[7]\ : SLE
      port map(D => \wptr_bin_sync[7]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[7]_net_1\);
    
    \rptr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[8]_net_1\, S
         => \rptr_s[9]\, Y => OPEN, FCO => \rptr_cry[9]_net_1\);
    
    \rptr_gray[5]\ : SLE
      port map(D => \rptr_gray_1[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[5]_net_1\);
    
    \wptr_gray_1[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[2]_net_1\, B => \wptr[3]_net_1\, Y => 
        \wptr_gray_1[2]_net_1\);
    
    \wptr[5]\ : SLE
      port map(D => \wptr_s[5]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[5]_net_1\);
    
    rdiff_bus_cry_5 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[5]_net_1\, B => 
        \rptr[5]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_4\, S => \rdiff_bus[5]\, Y => OPEN, FCO
         => \rdiff_bus_cry_5\);
    
    \wptr_bin_sync2[8]\ : SLE
      port map(D => \wptr_bin_sync[8]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[8]_net_1\);
    
    \wptr[7]\ : SLE
      port map(D => \wptr_s[7]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[7]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \wptr_gray[1]\ : SLE
      port map(D => \wptr_gray_1[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[1]_net_1\);
    
    \rptr_gray_1[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[9]_net_1\, B => \rptr[10]_net_1\, Y => 
        \rptr_gray_1[9]_net_1\);
    
    \rptr_bin_sync2[5]\ : SLE
      port map(D => \rptr_bin_sync[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[5]_net_1\);
    
    \rptr_bin_sync2[1]\ : SLE
      port map(D => \rptr_bin_sync[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[1]_net_1\);
    
    \memwaddr_r[10]\ : SLE
      port map(D => \memwaddr_r_s[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_248, ALn => irx_fifo_rst_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \fifo_MEMWADDR[10]\);
    
    wdiff_bus_cry_7 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[7]_net_1\, B => 
        \rptr_bin_sync2[7]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_6\, S => \wdiff_bus[7]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_7\);
    
    \wptr_bin_sync2[0]\ : SLE
      port map(D => \wptr_bin_sync[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rdiff_bus);
    
    \L1.un2_re_p_i_i_a3\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_1004, B => \iRX_FIFO_Empty_0\, Y => 
        un2_re_p_i_i_a3);
    
    \L1.empty_r_3_0_a2_1\ : CFG2
      generic map(INIT => x"1")

      port map(A => \rdiff_bus[4]\, B => \rdiff_bus[3]\, Y => 
        empty_r_3_0_a2_1);
    
    \L1.un1_we_p_0_a2_0_a2\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_248, B => \iRX_FIFO_Full_0\, Y => un1_we_p);
    
    rdiff_bus_s_11 : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \rptr[11]_net_1\, C => 
        \wptr_bin_sync2[11]_net_1\, D => GND_net_1, FCI => 
        \rdiff_bus_cry_10\, S => \rdiff_bus[11]\, Y => OPEN, FCO
         => OPEN);
    
    \memwaddr_r_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[8]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[7]_net_1\, S => \memwaddr_r_s[8]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[8]_net_1\);
    
    \wptr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => wptr_s_385_FCO, S => 
        \wptr_s[1]\, Y => OPEN, FCO => \wptr_cry[1]_net_1\);
    
    \memraddr_r[8]\ : SLE
      port map(D => \memraddr_r_s[8]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1007_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[8]\);
    
    \rptr[9]\ : SLE
      port map(D => \rptr_s[9]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1007_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[9]_net_1\);
    
    \wptr_gray_1[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[6]_net_1\, B => \wptr[7]_net_1\, Y => 
        \wptr_gray_1[6]_net_1\);
    
    \wptr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[6]_net_1\, S
         => \wptr_s[7]\, Y => OPEN, FCO => \wptr_cry[7]_net_1\);
    
    \wptr_bin_sync2[2]\ : SLE
      port map(D => \wptr_bin_sync[2]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[2]_net_1\);
    
    \rptr_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \rptr[0]_net_1\, Y => \rptr_s[0]\);
    
    \rptr[4]\ : SLE
      port map(D => \rptr_s[4]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1007_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[4]_net_1\);
    
    \memwaddr_r_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[4]_net_1\, S => \memwaddr_r_s[5]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[5]_net_1\);
    
    \memraddr_r_s[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[9]_net_1\, S => \memraddr_r_s[10]_net_1\, 
        Y => OPEN, FCO => OPEN);
    
    \wptr_gray[6]\ : SLE
      port map(D => \wptr_gray_1[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[6]_net_1\);
    
    \wptr_gray_1[3]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[3]_net_1\, B => \wptr[4]_net_1\, Y => 
        \wptr_gray_1[3]_net_1\);
    
    \wptr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[4]_net_1\, S
         => \wptr_s[5]\, Y => OPEN, FCO => \wptr_cry[5]_net_1\);
    
    \memraddr_r_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[4]_net_1\, S => \memraddr_r_s[5]\, Y => 
        OPEN, FCO => \memraddr_r_cry[5]_net_1\);
    
    \memraddr_r_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[1]\, C => 
        GND_net_1, D => GND_net_1, FCI => memraddr_r_s_384_FCO, S
         => \memraddr_r_s[1]\, Y => OPEN, FCO => 
        \memraddr_r_cry[1]_net_1\);
    
    \rptr_gray[4]\ : SLE
      port map(D => \rptr_gray_1[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[4]_net_1\);
    
    \wptr_bin_sync2[4]\ : SLE
      port map(D => \wptr_bin_sync[4]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[4]_net_1\);
    
    \wptr[3]\ : SLE
      port map(D => \wptr_s[3]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[3]_net_1\);
    
    \memwaddr_r[6]\ : SLE
      port map(D => \memwaddr_r_s[6]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_248, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[6]\);
    
    \wptr_s[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[10]_net_1\, S
         => \wptr_s[11]_net_1\, Y => OPEN, FCO => OPEN);
    
    \wptr[6]\ : SLE
      port map(D => \wptr_s[6]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[6]_net_1\);
    
    \memwaddr_r[9]\ : SLE
      port map(D => \memwaddr_r_s[9]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_248, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[9]\);
    
    \memraddr_r_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[3]_net_1\, S => \memraddr_r_s[4]\, Y => 
        OPEN, FCO => \memraddr_r_cry[4]_net_1\);
    
    \memraddr_r[10]\ : SLE
      port map(D => \memraddr_r_s[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1007_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[10]\);
    
    \memwaddr_r[3]\ : SLE
      port map(D => \memwaddr_r_s[3]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_248, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[3]\);
    
    full_r : SLE
      port map(D => fulli, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \iRX_FIFO_Full_0\);
    
    \rptr_bin_sync2[3]\ : SLE
      port map(D => \rptr_bin_sync[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[3]_net_1\);
    
    \wptr_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \wptr[0]_net_1\, Y => \wptr_s[0]\);
    
    \rptr[2]\ : SLE
      port map(D => \rptr_s[2]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1007_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[2]_net_1\);
    
    \memraddr_r[3]\ : SLE
      port map(D => \memraddr_r_s[3]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1007_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[3]\);
    
    \rptr_bin_sync2[9]\ : SLE
      port map(D => \rptr_bin_sync[9]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[9]_net_1\);
    
    \rptr[11]\ : SLE
      port map(D => \rptr_s[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1007_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rptr[11]_net_1\);
    
    \wptr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[5]_net_1\, S
         => \wptr_s[6]\, Y => OPEN, FCO => \wptr_cry[6]_net_1\);
    
    \rptr_bin_sync2[11]\ : SLE
      port map(D => \rptr_bin_sync[11]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[11]_net_1\);
    
    \wptr_bin_sync2[5]\ : SLE
      port map(D => \wptr_bin_sync[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[5]_net_1\);
    
    \wptr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[7]_net_1\, S
         => \wptr_s[8]\, Y => OPEN, FCO => \wptr_cry[8]_net_1\);
    
    \wptr_bin_sync2[1]\ : SLE
      port map(D => \wptr_bin_sync[1]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[1]_net_1\);
    
    Wr_corefifo_grayToBinConv : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_0
      port map(wptr_bin_sync(11) => \wptr_bin_sync[11]\, 
        wptr_bin_sync(10) => \wptr_bin_sync[10]\, 
        wptr_bin_sync(9) => \wptr_bin_sync[9]\, wptr_bin_sync(8)
         => \wptr_bin_sync[8]\, wptr_bin_sync(7) => 
        \wptr_bin_sync[7]\, wptr_bin_sync(6) => 
        \wptr_bin_sync[6]\, wptr_bin_sync(5) => 
        \wptr_bin_sync[5]\, wptr_bin_sync(4) => 
        \wptr_bin_sync[4]\, wptr_bin_sync(3) => 
        \wptr_bin_sync[3]\, wptr_bin_sync(2) => 
        \wptr_bin_sync[2]\, wptr_bin_sync(1) => 
        \wptr_bin_sync[1]\, wptr_bin_sync(0) => 
        \wptr_bin_sync[0]\, wptr_gray_sync(10) => 
        \wptr_gray_sync[10]\, wptr_gray_sync(9) => 
        \wptr_gray_sync[9]\, wptr_gray_sync(8) => 
        \wptr_gray_sync[8]\, wptr_gray_sync(7) => 
        \wptr_gray_sync[7]\, wptr_gray_sync(6) => 
        \wptr_gray_sync[6]\, wptr_gray_sync(5) => 
        \wptr_gray_sync[5]\, wptr_gray_sync(4) => 
        \wptr_gray_sync[4]\, wptr_gray_sync(3) => 
        \wptr_gray_sync[3]\, wptr_gray_sync(2) => 
        \wptr_gray_sync[2]\, wptr_gray_sync(1) => 
        \wptr_gray_sync[1]\, wptr_gray_sync(0) => 
        \wptr_gray_sync[0]\);
    
    \wptr_gray_1[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[4]_net_1\, B => \wptr[5]_net_1\, Y => 
        \wptr_gray_1[4]_net_1\);
    
    overflow_r : SLE
      port map(D => un1_we_p, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        iRX_FIFO_OVERFLOW_0);
    
    fulli_0 : CFG4
      generic map(INIT => x"EAAA")

      port map(A => \wdiff_bus[11]\, B => \fulli_0_a2_7\, C => 
        N_248, D => \fulli_0_a2_8\, Y => fulli);
    
    \memraddr_r_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \fifo_MEMRADDR[0]\, Y => \memraddr_r_s[0]\);
    
    \rptr_gray[11]\ : SLE
      port map(D => \rptr[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[11]_net_1\);
    
    \wptr_bin_sync2[10]\ : SLE
      port map(D => \wptr_bin_sync[10]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[10]_net_1\);
    
    \rptr[10]\ : SLE
      port map(D => \rptr_s[10]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1007_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rptr[10]_net_1\);
    
    \wptr[9]\ : SLE
      port map(D => \wptr_s[9]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[9]_net_1\);
    
    Wr_corefifo_doubleSync : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync
      port map(wptr_gray(11) => \wptr_gray[11]_net_1\, 
        wptr_gray(10) => \wptr_gray[10]_net_1\, wptr_gray(9) => 
        \wptr_gray[9]_net_1\, wptr_gray(8) => 
        \wptr_gray[8]_net_1\, wptr_gray(7) => 
        \wptr_gray[7]_net_1\, wptr_gray(6) => 
        \wptr_gray[6]_net_1\, wptr_gray(5) => 
        \wptr_gray[5]_net_1\, wptr_gray(4) => 
        \wptr_gray[4]_net_1\, wptr_gray(3) => 
        \wptr_gray[3]_net_1\, wptr_gray(2) => 
        \wptr_gray[2]_net_1\, wptr_gray(1) => 
        \wptr_gray[1]_net_1\, wptr_gray(0) => 
        \wptr_gray[0]_net_1\, wptr_gray_sync(10) => 
        \wptr_gray_sync[10]\, wptr_gray_sync(9) => 
        \wptr_gray_sync[9]\, wptr_gray_sync(8) => 
        \wptr_gray_sync[8]\, wptr_gray_sync(7) => 
        \wptr_gray_sync[7]\, wptr_gray_sync(6) => 
        \wptr_gray_sync[6]\, wptr_gray_sync(5) => 
        \wptr_gray_sync[5]\, wptr_gray_sync(4) => 
        \wptr_gray_sync[4]\, wptr_gray_sync(3) => 
        \wptr_gray_sync[3]\, wptr_gray_sync(2) => 
        \wptr_gray_sync[2]\, wptr_gray_sync(1) => 
        \wptr_gray_sync[1]\, wptr_gray_sync(0) => 
        \wptr_gray_sync[0]\, wptr_bin_sync_0 => 
        \wptr_bin_sync[11]\, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, irx_fifo_rst_i => 
        irx_fifo_rst_i);
    
    \rptr_gray[0]\ : SLE
      port map(D => \rptr_gray_1[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[0]_net_1\);
    
    empty_r : SLE
      port map(D => empty_r_3, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \iRX_FIFO_Empty_0\);
    
    \rptr_gray_1[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[7]_net_1\, B => \rptr[8]_net_1\, Y => 
        \rptr_gray_1[7]_net_1\);
    
    fulli_0_a2_0_0_a2_1 : CFG4
      generic map(INIT => x"0080")

      port map(A => iRX_FIFO_wr_en, B => sampler_clk1x_en, C => 
        RX_InProcess_d1, D => tx_col_detect_en, Y => \N_1466\);
    
    \wptr[4]\ : SLE
      port map(D => \wptr_s[4]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[4]_net_1\);
    
    \memwaddr_r[8]\ : SLE
      port map(D => \memwaddr_r_s[8]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_248, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[8]\);
    
    \memwaddr_r[2]\ : SLE
      port map(D => \memwaddr_r_s[2]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_248, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[2]\);
    
    \L1.empty_r_3_0_a2_5\ : CFG3
      generic map(INIT => x"0E")

      port map(A => N_1004, B => rdiff_bus_cry_0_Y_0, C => 
        \rdiff_bus[11]\, Y => empty_r_3_0_a2_5);
    
    \wptr_bin_sync2[11]\ : SLE
      port map(D => \wptr_bin_sync[11]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[11]_net_1\);
    
    \wptr_gray_1[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[1]_net_1\, B => \wptr[2]_net_1\, Y => 
        \wptr_gray_1[1]_net_1\);
    
    underflow_r : SLE
      port map(D => un2_re_p_i_i_a3, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => iRX_FIFO_UNDERRUN_0);
    
    \memwaddr_r_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[6]_net_1\, S => \memwaddr_r_s[7]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[7]_net_1\);
    
    \wptr_gray[5]\ : SLE
      port map(D => \wptr_gray_1[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[5]_net_1\);
    
    \memraddr_r[7]\ : SLE
      port map(D => \memraddr_r_s[7]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1007_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[7]\);
    
    memwe_0_a2_0_a2 : CFG4
      generic map(INIT => x"0010")

      port map(A => ReadFIFO_Write_Ptr(1), B => \iRX_FIFO_Full_0\, 
        C => \N_1466\, D => ReadFIFO_Write_Ptr(0), Y => 
        \fifo_MEMWE\);
    
    \rptr_bin_sync2[10]\ : SLE
      port map(D => \rptr_bin_sync[10]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[10]_net_1\);
    
    wdiff_bus_cry_10 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[10]_net_1\, B => 
        \rptr_bin_sync2[10]_net_1\, C => GND_net_1, D => 
        GND_net_1, FCI => \wdiff_bus_cry_9\, S => \wdiff_bus[10]\, 
        Y => OPEN, FCO => \wdiff_bus_cry_10\);
    
    \memwaddr_r_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[9]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[8]_net_1\, S => \memwaddr_r_s[9]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[9]_net_1\);
    
    \wptr_gray[8]\ : SLE
      port map(D => \wptr_gray_1[8]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[8]_net_1\);
    
    \wptr_gray[7]\ : SLE
      port map(D => \wptr_gray_1[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[7]_net_1\);
    
    \wptr_gray_1[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[5]_net_1\, B => \wptr[6]_net_1\, Y => 
        \wptr_gray_1[5]_net_1\);
    
    \memwaddr_r[5]\ : SLE
      port map(D => \memwaddr_r_s[5]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_248, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[5]\);
    
    \L1.empty_r_3_0_a2\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \rdiff_bus[9]\, B => \rdiff_bus[10]\, C => 
        empty_r_3_0_a2_5, D => empty_r_3_0_a2_9, Y => empty_r_3);
    
    \rptr[8]\ : SLE
      port map(D => \rptr_s[8]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1007_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[8]_net_1\);
    
    Rd_corefifo_doubleSync : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0
      port map(rptr_gray(11) => \rptr_gray[11]_net_1\, 
        rptr_gray(10) => \rptr_gray[10]_net_1\, rptr_gray(9) => 
        \rptr_gray[9]_net_1\, rptr_gray(8) => 
        \rptr_gray[8]_net_1\, rptr_gray(7) => 
        \rptr_gray[7]_net_1\, rptr_gray(6) => 
        \rptr_gray[6]_net_1\, rptr_gray(5) => 
        \rptr_gray[5]_net_1\, rptr_gray(4) => 
        \rptr_gray[4]_net_1\, rptr_gray(3) => 
        \rptr_gray[3]_net_1\, rptr_gray(2) => 
        \rptr_gray[2]_net_1\, rptr_gray(1) => 
        \rptr_gray[1]_net_1\, rptr_gray(0) => 
        \rptr_gray[0]_net_1\, rptr_gray_sync(10) => 
        \rptr_gray_sync[10]\, rptr_gray_sync(9) => 
        \rptr_gray_sync[9]\, rptr_gray_sync(8) => 
        \rptr_gray_sync[8]\, rptr_gray_sync(7) => 
        \rptr_gray_sync[7]\, rptr_gray_sync(6) => 
        \rptr_gray_sync[6]\, rptr_gray_sync(5) => 
        \rptr_gray_sync[5]\, rptr_gray_sync(4) => 
        \rptr_gray_sync[4]\, rptr_gray_sync(3) => 
        \rptr_gray_sync[3]\, rptr_gray_sync(2) => 
        \rptr_gray_sync[2]\, rptr_gray_sync(1) => 
        \rptr_gray_sync[1]\, rptr_gray_sync(0) => 
        \rptr_gray_sync[0]\, rptr_bin_sync_0 => 
        \rptr_bin_sync[11]\, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, irx_fifo_rst_i => irx_fifo_rst_i);
    
    \rptr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[3]_net_1\, S
         => \rptr_s[4]\, Y => OPEN, FCO => \rptr_cry[4]_net_1\);
    
    wdiff_bus_cry_2 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[2]_net_1\, B => 
        \rptr_bin_sync2[2]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_1\, S => \wdiff_bus[2]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_2\);
    
    \rptr_gray[2]\ : SLE
      port map(D => \rptr_gray_1[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[2]_net_1\);
    
    \wptr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[8]_net_1\, S
         => \wptr_s[9]\, Y => OPEN, FCO => \wptr_cry[9]_net_1\);
    
    \wptr_bin_sync2[3]\ : SLE
      port map(D => \wptr_bin_sync[3]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[3]_net_1\);
    
    \wptr[2]\ : SLE
      port map(D => \wptr_s[2]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[2]_net_1\);
    
    \rptr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[1]_net_1\, S
         => \rptr_s[2]\, Y => OPEN, FCO => \rptr_cry[2]_net_1\);
    
    rdiff_bus_cry_9 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[9]_net_1\, B => 
        \rptr[9]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_8\, S => \rdiff_bus[9]\, Y => OPEN, FCO
         => \rdiff_bus_cry_9\);
    
    \memwaddr_r[0]\ : SLE
      port map(D => \memwaddr_r_s[0]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_248, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMWADDR[0]\);
    
    fulli_0_a2_7 : CFG4
      generic map(INIT => x"8000")

      port map(A => \wdiff_bus[6]\, B => \wdiff_bus[7]\, C => 
        \wdiff_bus[8]\, D => \wdiff_bus[9]\, Y => \fulli_0_a2_7\);
    
    \wptr_gray[2]\ : SLE
      port map(D => \wptr_gray_1[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[2]_net_1\);
    
    wdiff_bus_cry_4 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[4]_net_1\, B => 
        \rptr_bin_sync2[4]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_3\, S => \wdiff_bus[4]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_4\);
    
    \memwaddr_r_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[2]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[1]_net_1\, S => \memwaddr_r_s[2]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[2]_net_1\);
    
    \wptr_gray[11]\ : SLE
      port map(D => \wptr[11]_net_1\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr_gray[11]_net_1\);
    
    \wptr_bin_sync2[9]\ : SLE
      port map(D => \wptr_bin_sync[9]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[9]_net_1\);
    
    \rptr_gray_1[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[6]_net_1\, B => \rptr[7]_net_1\, Y => 
        \rptr_gray_1[6]_net_1\);
    
    \wptr_gray_1[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[11]_net_1\, B => \wptr[10]_net_1\, Y
         => \wptr_gray_1[10]_net_1\);
    
    wdiff_bus_cry_6 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[6]_net_1\, B => 
        \rptr_bin_sync2[6]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_5\, S => \wdiff_bus[6]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_6\);
    
    \rptr_s[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[10]_net_1\, S
         => \rptr_s[11]_net_1\, Y => OPEN, FCO => OPEN);
    
    \rptr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[2]_net_1\, S
         => \rptr_s[3]\, Y => OPEN, FCO => \rptr_cry[3]_net_1\);
    
    \memraddr_r[4]\ : SLE
      port map(D => \memraddr_r_s[4]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1007_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[4]\);
    
    \memraddr_r_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[6]_net_1\, S => \memraddr_r_s[7]\, Y => 
        OPEN, FCO => \memraddr_r_cry[7]_net_1\);
    
    fulli_0_a2_8 : CFG4
      generic map(INIT => x"4000")

      port map(A => wdiff_bus_cry_0_Y_0, B => \wdiff_bus[1]\, C
         => \wdiff_bus[10]\, D => \fulli_0_a2_6\, Y => 
        \fulli_0_a2_8\);
    
    memraddr_r_s_384 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[0]\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => memraddr_r_s_384_FCO);
    
    \memraddr_r_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[9]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[8]_net_1\, S => \memraddr_r_s[9]\, Y => 
        OPEN, FCO => \memraddr_r_cry[9]_net_1\);
    
    \memraddr_r[5]\ : SLE
      port map(D => \memraddr_r_s[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1007_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[5]\);
    
    \rptr_gray[6]\ : SLE
      port map(D => \rptr_gray_1[6]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[6]_net_1\);
    
    \memraddr_r[9]\ : SLE
      port map(D => \memraddr_r_s[9]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1007_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[9]\);
    
    \rptr[0]\ : SLE
      port map(D => \rptr_s[0]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \N_1007_i\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr[0]_net_1\);
    
    wptr_s_385 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => wptr_s_385_FCO);
    
    \wptr[10]\ : SLE
      port map(D => \wptr_s[10]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[10]_net_1\);
    
    \memwaddr_r_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[3]_net_1\, S => \memwaddr_r_s[4]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[4]_net_1\);
    
    \memraddr_r_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[3]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[2]_net_1\, S => \memraddr_r_s[3]\, Y => 
        OPEN, FCO => \memraddr_r_cry[3]_net_1\);
    
    wdiff_bus_cry_1 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[1]_net_1\, B => 
        \rptr_bin_sync2[1]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_0\, S => \wdiff_bus[1]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_1\);
    
    rdiff_bus_cry_2 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[2]_net_1\, B => 
        \rptr[2]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_1\, S => \rdiff_bus[2]\, Y => OPEN, FCO
         => \rdiff_bus_cry_2\);
    
    \wptr_gray[9]\ : SLE
      port map(D => \wptr_gray_1[9]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[9]_net_1\);
    
    \rptr_gray_1[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[4]_net_1\, B => \rptr[5]_net_1\, Y => 
        \rptr_gray_1[4]_net_1\);
    
    \wptr_gray_1[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[8]_net_1\, B => \wptr[9]_net_1\, Y => 
        \wptr_gray_1[8]_net_1\);
    
    Rd_corefifo_grayToBinConv : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3
      port map(rptr_bin_sync(11) => \rptr_bin_sync[11]\, 
        rptr_bin_sync(10) => \rptr_bin_sync[10]\, 
        rptr_bin_sync(9) => \rptr_bin_sync[9]\, rptr_bin_sync(8)
         => \rptr_bin_sync[8]\, rptr_bin_sync(7) => 
        \rptr_bin_sync[7]\, rptr_bin_sync(6) => 
        \rptr_bin_sync[6]\, rptr_bin_sync(5) => 
        \rptr_bin_sync[5]\, rptr_bin_sync(4) => 
        \rptr_bin_sync[4]\, rptr_bin_sync(3) => 
        \rptr_bin_sync[3]\, rptr_bin_sync(2) => 
        \rptr_bin_sync[2]\, rptr_bin_sync(1) => 
        \rptr_bin_sync[1]\, rptr_bin_sync(0) => 
        \rptr_bin_sync[0]\, rptr_gray_sync(10) => 
        \rptr_gray_sync[10]\, rptr_gray_sync(9) => 
        \rptr_gray_sync[9]\, rptr_gray_sync(8) => 
        \rptr_gray_sync[8]\, rptr_gray_sync(7) => 
        \rptr_gray_sync[7]\, rptr_gray_sync(6) => 
        \rptr_gray_sync[6]\, rptr_gray_sync(5) => 
        \rptr_gray_sync[5]\, rptr_gray_sync(4) => 
        \rptr_gray_sync[4]\, rptr_gray_sync(3) => 
        \rptr_gray_sync[3]\, rptr_gray_sync(2) => 
        \rptr_gray_sync[2]\, rptr_gray_sync(1) => 
        \rptr_gray_sync[1]\, rptr_gray_sync(0) => 
        \rptr_gray_sync[0]\);
    
    \rptr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => rptr_s_383_FCO, S => 
        \rptr_s[1]\, Y => OPEN, FCO => \rptr_cry[1]_net_1\);
    
    rdiff_bus_cry_3 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[3]_net_1\, B => 
        \rptr[3]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_2\, S => \rdiff_bus[3]\, Y => OPEN, FCO
         => \rdiff_bus_cry_3\);
    
    rdiff_bus_cry_10 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[10]_net_1\, B => 
        \rptr[10]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_9\, S => \rdiff_bus[10]\, Y => OPEN, FCO
         => \rdiff_bus_cry_10\);
    
    \memraddr_r_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[5]_net_1\, S => \memraddr_r_s[6]\, Y => 
        OPEN, FCO => \memraddr_r_cry[6]_net_1\);
    
    \memraddr_r[6]\ : SLE
      port map(D => \memraddr_r_s[6]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1007_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[6]\);
    
    \rptr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[6]_net_1\, S
         => \rptr_s[7]\, Y => OPEN, FCO => \rptr_cry[7]_net_1\);
    
    rdiff_bus_cry_0 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => rdiff_bus, B => \rptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => rdiff_bus_cry_0_Y_0, FCO => \rdiff_bus_cry_0\);
    
    \memraddr_r[2]\ : SLE
      port map(D => \memraddr_r_s[2]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \N_1007_i\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[2]\);
    
    \wptr[8]\ : SLE
      port map(D => \wptr_s[8]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[8]_net_1\);
    
    empty_r_RNIUREJ1_0 : CFG3
      generic map(INIT => x"A2")

      port map(A => REN_d1, B => N_1004, C => \iRX_FIFO_Empty_0\, 
        Y => N_89_i);
    
    wdiff_bus_cry_3 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[3]_net_1\, B => 
        \rptr_bin_sync2[3]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_2\, S => \wdiff_bus[3]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_3\);
    
    \rptr_gray[7]\ : SLE
      port map(D => \rptr_gray_1[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[7]_net_1\);
    
    \wptr_gray[0]\ : SLE
      port map(D => \wptr_gray_1[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[0]_net_1\);
    
    \rptr_gray_1[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[0]_net_1\, B => \rptr[1]_net_1\, Y => 
        \rptr_gray_1[0]_net_1\);
    
    \rptr_gray_1[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[8]_net_1\, B => \rptr[9]_net_1\, Y => 
        \rptr_gray_1[8]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO is

    port( RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          ReadFIFO_Write_Ptr        : in    std_logic_vector(1 downto 0);
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          RX_FIFO_DOUT_0_0          : out   std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          N_1466                    : out   std_logic;
          iRX_FIFO_wr_en            : in    std_logic;
          sampler_clk1x_en          : in    std_logic;
          RX_InProcess_d1           : in    std_logic;
          tx_col_detect_en          : in    std_logic;
          N_653                     : out   std_logic;
          N_655                     : out   std_logic;
          N_656                     : out   std_logic;
          N_718                     : out   std_logic;
          N_654                     : out   std_logic;
          N_652                     : out   std_logic;
          N_651                     : out   std_logic;
          N_650                     : out   std_logic;
          N_1004                    : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          irx_fifo_rst_i            : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper
    port( RDATA_int                 : out   std_logic_vector(8 downto 0);
          fifo_MEMRADDR             : in    std_logic_vector(10 downto 0) := (others => 'U');
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          fifo_MEMWADDR             : in    std_logic_vector(10 downto 0) := (others => 'U');
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          N_1007_i                  : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          fifo_MEMWE                : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3
    port( ReadFIFO_Write_Ptr        : in    std_logic_vector(1 downto 0) := (others => 'U');
          fifo_MEMWADDR             : out   std_logic_vector(10 downto 0);
          fifo_MEMRADDR             : out   std_logic_vector(10 downto 0);
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          N_153_i_i                 : out   std_logic;
          N_89_i                    : out   std_logic;
          REN_d1                    : in    std_logic := 'U';
          N_1004                    : in    std_logic := 'U';
          tx_col_detect_en          : in    std_logic := 'U';
          RX_InProcess_d1           : in    std_logic := 'U';
          sampler_clk1x_en          : in    std_logic := 'U';
          iRX_FIFO_wr_en            : in    std_logic := 'U';
          N_1466                    : out   std_logic;
          N_1007_i                  : out   std_logic;
          fifo_MEMWE                : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          irx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \RDATA_r[4]_net_1\, VCC_net_1, \RDATA_int[4]\, N_89_i, 
        GND_net_1, \RDATA_r[5]_net_1\, \RDATA_int[5]\, 
        \RDATA_r[6]_net_1\, \RDATA_int[6]\, \RDATA_r[7]_net_1\, 
        \RDATA_int[7]\, \RDATA_r[8]_net_1\, \RDATA_int[8]\, 
        \re_set\, \REN_d1\, N_153_i_i, \RDATA_r[0]_net_1\, 
        \RDATA_int[0]\, \RDATA_r[1]_net_1\, \RDATA_int[1]\, 
        \RDATA_r[2]_net_1\, \RDATA_int[2]\, \RDATA_r[3]_net_1\, 
        \RDATA_int[3]\, N_1007_i, \RE_d1\, \re_pulse_d1\, 
        \re_pulse\, \iRX_FIFO_Empty_0\, \fifo_MEMWADDR[0]\, 
        \fifo_MEMWADDR[1]\, \fifo_MEMWADDR[2]\, 
        \fifo_MEMWADDR[3]\, \fifo_MEMWADDR[4]\, 
        \fifo_MEMWADDR[5]\, \fifo_MEMWADDR[6]\, 
        \fifo_MEMWADDR[7]\, \fifo_MEMWADDR[8]\, 
        \fifo_MEMWADDR[9]\, \fifo_MEMWADDR[10]\, 
        \fifo_MEMRADDR[0]\, \fifo_MEMRADDR[1]\, 
        \fifo_MEMRADDR[2]\, \fifo_MEMRADDR[3]\, 
        \fifo_MEMRADDR[4]\, \fifo_MEMRADDR[5]\, 
        \fifo_MEMRADDR[6]\, \fifo_MEMRADDR[7]\, 
        \fifo_MEMRADDR[8]\, \fifo_MEMRADDR[9]\, 
        \fifo_MEMRADDR[10]\, fifo_MEMWE : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3(DEF_ARCH);
begin 

    iRX_FIFO_Empty_0 <= \iRX_FIFO_Empty_0\;

    re_pulse : CFG4
      generic map(INIT => x"FAF2")

      port map(A => \REN_d1\, B => N_1004, C => \re_set\, D => 
        \iRX_FIFO_Empty_0\, Y => \re_pulse\);
    
    \RDATA_r[3]\ : SLE
      port map(D => \RDATA_int[3]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[3]_net_1\);
    
    \Q_i_m2[2]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[2]_net_1\, C => 
        \RDATA_int[2]\, D => \RE_d1\, Y => N_651);
    
    re_pulse_d1 : SLE
      port map(D => \re_pulse\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \re_pulse_d1\);
    
    \RDATA_r[5]\ : SLE
      port map(D => \RDATA_int[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[5]_net_1\);
    
    \Q_i_m2[0]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[0]_net_1\, C => 
        \RDATA_int[0]\, D => \RE_d1\, Y => N_650);
    
    \Q_i_m2[3]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[3]_net_1\, C => 
        \RDATA_int[3]\, D => \RE_d1\, Y => N_652);
    
    \RDATA_r[8]\ : SLE
      port map(D => \RDATA_int[8]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[8]_net_1\);
    
    \Q_i_m2[7]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[7]_net_1\, C => 
        \RDATA_int[7]\, D => \RE_d1\, Y => N_656);
    
    \Q_i_m2[6]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[6]_net_1\, C => 
        \RDATA_int[6]\, D => \RE_d1\, Y => N_655);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \RW1.UI_ram_wrapper_1\ : FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper
      port map(RDATA_int(8) => \RDATA_int[8]\, RDATA_int(7) => 
        \RDATA_int[7]\, RDATA_int(6) => \RDATA_int[6]\, 
        RDATA_int(5) => \RDATA_int[5]\, RDATA_int(4) => 
        \RDATA_int[4]\, RDATA_int(3) => \RDATA_int[3]\, 
        RDATA_int(2) => \RDATA_int[2]\, RDATA_int(1) => 
        \RDATA_int[1]\, RDATA_int(0) => \RDATA_int[0]\, 
        fifo_MEMRADDR(10) => \fifo_MEMRADDR[10]\, 
        fifo_MEMRADDR(9) => \fifo_MEMRADDR[9]\, fifo_MEMRADDR(8)
         => \fifo_MEMRADDR[8]\, fifo_MEMRADDR(7) => 
        \fifo_MEMRADDR[7]\, fifo_MEMRADDR(6) => 
        \fifo_MEMRADDR[6]\, fifo_MEMRADDR(5) => 
        \fifo_MEMRADDR[5]\, fifo_MEMRADDR(4) => 
        \fifo_MEMRADDR[4]\, fifo_MEMRADDR(3) => 
        \fifo_MEMRADDR[3]\, fifo_MEMRADDR(2) => 
        \fifo_MEMRADDR[2]\, fifo_MEMRADDR(1) => 
        \fifo_MEMRADDR[1]\, fifo_MEMRADDR(0) => 
        \fifo_MEMRADDR[0]\, RX_FIFO_DIN_pipe(8) => 
        RX_FIFO_DIN_pipe(8), RX_FIFO_DIN_pipe(7) => 
        RX_FIFO_DIN_pipe(7), RX_FIFO_DIN_pipe(6) => 
        RX_FIFO_DIN_pipe(6), RX_FIFO_DIN_pipe(5) => 
        RX_FIFO_DIN_pipe(5), RX_FIFO_DIN_pipe(4) => 
        RX_FIFO_DIN_pipe(4), RX_FIFO_DIN_pipe(3) => 
        RX_FIFO_DIN_pipe(3), RX_FIFO_DIN_pipe(2) => 
        RX_FIFO_DIN_pipe(2), RX_FIFO_DIN_pipe(1) => 
        RX_FIFO_DIN_pipe(1), RX_FIFO_DIN_pipe(0) => 
        RX_FIFO_DIN_pipe(0), fifo_MEMWADDR(10) => 
        \fifo_MEMWADDR[10]\, fifo_MEMWADDR(9) => 
        \fifo_MEMWADDR[9]\, fifo_MEMWADDR(8) => 
        \fifo_MEMWADDR[8]\, fifo_MEMWADDR(7) => 
        \fifo_MEMWADDR[7]\, fifo_MEMWADDR(6) => 
        \fifo_MEMWADDR[6]\, fifo_MEMWADDR(5) => 
        \fifo_MEMWADDR[5]\, fifo_MEMWADDR(4) => 
        \fifo_MEMWADDR[4]\, fifo_MEMWADDR(3) => 
        \fifo_MEMWADDR[3]\, fifo_MEMWADDR(2) => 
        \fifo_MEMWADDR[2]\, fifo_MEMWADDR(1) => 
        \fifo_MEMWADDR[1]\, fifo_MEMWADDR(0) => 
        \fifo_MEMWADDR[0]\, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, N_1007_i => N_1007_i, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, fifo_MEMWE
         => fifo_MEMWE);
    
    \RDATA_r[0]\ : SLE
      port map(D => \RDATA_int[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[0]_net_1\);
    
    \Q_i_m2[5]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[5]_net_1\, C => 
        \RDATA_int[5]\, D => \RE_d1\, Y => N_654);
    
    \RDATA_r[2]\ : SLE
      port map(D => \RDATA_int[2]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[2]_net_1\);
    
    \RDATA_r[6]\ : SLE
      port map(D => \RDATA_int[6]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[6]_net_1\);
    
    \L31.U_corefifo_async\ : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3
      port map(ReadFIFO_Write_Ptr(1) => ReadFIFO_Write_Ptr(1), 
        ReadFIFO_Write_Ptr(0) => ReadFIFO_Write_Ptr(0), 
        fifo_MEMWADDR(10) => \fifo_MEMWADDR[10]\, 
        fifo_MEMWADDR(9) => \fifo_MEMWADDR[9]\, fifo_MEMWADDR(8)
         => \fifo_MEMWADDR[8]\, fifo_MEMWADDR(7) => 
        \fifo_MEMWADDR[7]\, fifo_MEMWADDR(6) => 
        \fifo_MEMWADDR[6]\, fifo_MEMWADDR(5) => 
        \fifo_MEMWADDR[5]\, fifo_MEMWADDR(4) => 
        \fifo_MEMWADDR[4]\, fifo_MEMWADDR(3) => 
        \fifo_MEMWADDR[3]\, fifo_MEMWADDR(2) => 
        \fifo_MEMWADDR[2]\, fifo_MEMWADDR(1) => 
        \fifo_MEMWADDR[1]\, fifo_MEMWADDR(0) => 
        \fifo_MEMWADDR[0]\, fifo_MEMRADDR(10) => 
        \fifo_MEMRADDR[10]\, fifo_MEMRADDR(9) => 
        \fifo_MEMRADDR[9]\, fifo_MEMRADDR(8) => 
        \fifo_MEMRADDR[8]\, fifo_MEMRADDR(7) => 
        \fifo_MEMRADDR[7]\, fifo_MEMRADDR(6) => 
        \fifo_MEMRADDR[6]\, fifo_MEMRADDR(5) => 
        \fifo_MEMRADDR[5]\, fifo_MEMRADDR(4) => 
        \fifo_MEMRADDR[4]\, fifo_MEMRADDR(3) => 
        \fifo_MEMRADDR[3]\, fifo_MEMRADDR(2) => 
        \fifo_MEMRADDR[2]\, fifo_MEMRADDR(1) => 
        \fifo_MEMRADDR[1]\, fifo_MEMRADDR(0) => 
        \fifo_MEMRADDR[0]\, iRX_FIFO_Empty_0 => 
        \iRX_FIFO_Empty_0\, iRX_FIFO_UNDERRUN_0 => 
        iRX_FIFO_UNDERRUN_0, iRX_FIFO_Full_0 => iRX_FIFO_Full_0, 
        iRX_FIFO_OVERFLOW_0 => iRX_FIFO_OVERFLOW_0, N_153_i_i => 
        N_153_i_i, N_89_i => N_89_i, REN_d1 => \REN_d1\, N_1004
         => N_1004, tx_col_detect_en => tx_col_detect_en, 
        RX_InProcess_d1 => RX_InProcess_d1, sampler_clk1x_en => 
        sampler_clk1x_en, iRX_FIFO_wr_en => iRX_FIFO_wr_en, 
        N_1466 => N_1466, N_1007_i => N_1007_i, fifo_MEMWE => 
        fifo_MEMWE, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, irx_fifo_rst_i => irx_fifo_rst_i);
    
    re_set : SLE
      port map(D => \REN_d1\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => N_153_i_i, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \re_set\);
    
    \Q_i_m2[8]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[8]_net_1\, C => 
        \RDATA_int[8]\, D => \RE_d1\, Y => N_718);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    RE_d1 : SLE
      port map(D => N_1004, CLK => m2s010_som_sb_0_CCC_71MHz, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \RE_d1\);
    
    \RDATA_r[7]\ : SLE
      port map(D => \RDATA_int[7]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[7]_net_1\);
    
    \RDATA_r[4]\ : SLE
      port map(D => \RDATA_int[4]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[4]_net_1\);
    
    \Q[1]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[1]_net_1\, C => 
        \RDATA_int[1]\, D => \RE_d1\, Y => RX_FIFO_DOUT_0_0);
    
    REN_d1 : SLE
      port map(D => N_1007_i, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \REN_d1\);
    
    \Q_i_m2[4]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[4]_net_1\, C => 
        \RDATA_int[4]\, D => \RE_d1\, Y => N_653);
    
    \RDATA_r[1]\ : SLE
      port map(D => \RDATA_int[1]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_89_i, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RDATA_r[1]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9 is

    port( ReadFIFO_Write_Ptr        : in    std_logic_vector(1 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          RX_FIFO_DOUT_0_0          : out   std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          irx_fifo_rst_i            : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          N_1004                    : in    std_logic;
          N_650                     : out   std_logic;
          N_651                     : out   std_logic;
          N_652                     : out   std_logic;
          N_654                     : out   std_logic;
          N_718                     : out   std_logic;
          N_656                     : out   std_logic;
          N_655                     : out   std_logic;
          N_653                     : out   std_logic;
          tx_col_detect_en          : in    std_logic;
          RX_InProcess_d1           : in    std_logic;
          sampler_clk1x_en          : in    std_logic;
          iRX_FIFO_wr_en            : in    std_logic;
          N_1466                    : out   std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic
        );

end FIFO_8Kx9;

architecture DEF_ARCH of FIFO_8Kx9 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO
    port( RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          ReadFIFO_Write_Ptr        : in    std_logic_vector(1 downto 0) := (others => 'U');
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          RX_FIFO_DOUT_0_0          : out   std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          N_1466                    : out   std_logic;
          iRX_FIFO_wr_en            : in    std_logic := 'U';
          sampler_clk1x_en          : in    std_logic := 'U';
          RX_InProcess_d1           : in    std_logic := 'U';
          tx_col_detect_en          : in    std_logic := 'U';
          N_653                     : out   std_logic;
          N_655                     : out   std_logic;
          N_656                     : out   std_logic;
          N_718                     : out   std_logic;
          N_654                     : out   std_logic;
          N_652                     : out   std_logic;
          N_651                     : out   std_logic;
          N_650                     : out   std_logic;
          N_1004                    : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          irx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    FIFO_8Kx9_0 : FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO
      port map(RX_FIFO_DIN_pipe(8) => RX_FIFO_DIN_pipe(8), 
        RX_FIFO_DIN_pipe(7) => RX_FIFO_DIN_pipe(7), 
        RX_FIFO_DIN_pipe(6) => RX_FIFO_DIN_pipe(6), 
        RX_FIFO_DIN_pipe(5) => RX_FIFO_DIN_pipe(5), 
        RX_FIFO_DIN_pipe(4) => RX_FIFO_DIN_pipe(4), 
        RX_FIFO_DIN_pipe(3) => RX_FIFO_DIN_pipe(3), 
        RX_FIFO_DIN_pipe(2) => RX_FIFO_DIN_pipe(2), 
        RX_FIFO_DIN_pipe(1) => RX_FIFO_DIN_pipe(1), 
        RX_FIFO_DIN_pipe(0) => RX_FIFO_DIN_pipe(0), 
        ReadFIFO_Write_Ptr(1) => ReadFIFO_Write_Ptr(1), 
        ReadFIFO_Write_Ptr(0) => ReadFIFO_Write_Ptr(0), 
        iRX_FIFO_OVERFLOW_0 => iRX_FIFO_OVERFLOW_0, 
        iRX_FIFO_Full_0 => iRX_FIFO_Full_0, iRX_FIFO_UNDERRUN_0
         => iRX_FIFO_UNDERRUN_0, iRX_FIFO_Empty_0 => 
        iRX_FIFO_Empty_0, RX_FIFO_DOUT_0_0 => RX_FIFO_DOUT_0_0, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, N_1466 => 
        N_1466, iRX_FIFO_wr_en => iRX_FIFO_wr_en, 
        sampler_clk1x_en => sampler_clk1x_en, RX_InProcess_d1 => 
        RX_InProcess_d1, tx_col_detect_en => tx_col_detect_en, 
        N_653 => N_653, N_655 => N_655, N_656 => N_656, N_718 => 
        N_718, N_654 => N_654, N_652 => N_652, N_651 => N_651, 
        N_650 => N_650, N_1004 => N_1004, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz, 
        irx_fifo_rst_i => irx_fifo_rst_i);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFOs is

    port( iRX_FIFO_Full                   : out   std_logic_vector(3 downto 0);
          RX_FIFO_DIN_pipe                : in    std_logic_vector(8 downto 0);
          CoreAPB3_0_APBmslave0_PWDATA    : in    std_logic_vector(7 downto 0);
          up_EOP_sync                     : in    std_logic_vector(2 downto 1);
          RX_FIFO_DOUT                    : out   std_logic_vector(7 downto 5);
          ReadFIFO_Read_Ptr               : out   std_logic_vector(1 downto 0);
          RX_FIFO_DOUT_3_0                : out   std_logic;
          RX_FIFO_DOUT_2_0                : out   std_logic;
          RX_FIFO_DOUT_1_0                : out   std_logic;
          RX_FIFO_DOUT_0_0                : out   std_logic;
          N_674                           : out   std_logic;
          N_673                           : out   std_logic;
          N_672                           : out   std_logic;
          N_667                           : out   std_logic;
          N_666                           : out   std_logic;
          N_665                           : out   std_logic;
          N_660                           : out   std_logic;
          N_659                           : out   std_logic;
          N_658                           : out   std_logic;
          iRX_FIFO_wr_en                  : in    std_logic;
          sampler_clk1x_en                : in    std_logic;
          RX_InProcess_d1                 : in    std_logic;
          tx_col_detect_en                : in    std_logic;
          N_653                           : out   std_logic;
          N_652                           : out   std_logic;
          N_651                           : out   std_logic;
          TX_FIFO_UNDERRUN                : out   std_logic;
          TX_FIFO_UNDERRUN_i              : out   std_logic;
          TX_FIFO_OVERFLOW                : out   std_logic;
          TX_FIFO_OVERFLOW_i              : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz       : in    std_logic;
          TX_FIFO_Full                    : out   std_logic;
          TX_FIFO_wr_en                   : in    std_logic;
          un1_tx_packet_length_0_sqmuxa_o : in    std_logic;
          TX_DataEn_1_o                   : in    std_logic;
          TX_PreAmble                     : in    std_logic;
          N_704                           : out   std_logic;
          N_705                           : out   std_logic;
          N_706                           : out   std_logic;
          N_707                           : out   std_logic;
          N_708                           : out   std_logic;
          N_709                           : out   std_logic;
          N_710                           : out   std_logic;
          N_711                           : out   std_logic;
          byte_clk_en                     : in    std_logic;
          TX_FIFO_Empty                   : out   std_logic;
          BIT_CLK                         : in    std_logic;
          RX_FIFO_RST                     : in    std_logic;
          RX_FIFO_rd_en                   : in    std_logic;
          TX_FIFO_RST                     : in    std_logic;
          un2_apb3_reset                  : in    std_logic;
          rx_packet_complt                : in    std_logic;
          N_678                           : out   std_logic;
          N_712                           : out   std_logic;
          N_693                           : out   std_logic;
          CommsFPGA_CCC_0_GL0             : in    std_logic;
          RX_FIFO_OVERFLOW_i              : out   std_logic;
          RX_FIFO_OVERFLOW                : out   std_logic;
          RX_FIFO_UNDERRUN_i              : out   std_logic;
          RX_FIFO_UNDERRUN                : out   std_logic
        );

end FIFOs;

architecture DEF_ARCH of FIFOs is 

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component FIFO_2Kx8
    port( CoreAPB3_0_APBmslave0_PWDATA    : in    std_logic_vector(7 downto 0) := (others => 'U');
          itx_fifo_rst_i                  : in    std_logic := 'U';
          BIT_CLK                         : in    std_logic := 'U';
          TX_FIFO_Empty                   : out   std_logic;
          byte_clk_en                     : in    std_logic := 'U';
          N_711                           : out   std_logic;
          N_710                           : out   std_logic;
          N_709                           : out   std_logic;
          N_708                           : out   std_logic;
          N_707                           : out   std_logic;
          N_706                           : out   std_logic;
          N_705                           : out   std_logic;
          N_704                           : out   std_logic;
          TX_PreAmble                     : in    std_logic := 'U';
          TX_DataEn_1_o                   : in    std_logic := 'U';
          un1_tx_packet_length_0_sqmuxa_o : in    std_logic := 'U';
          TX_FIFO_wr_en                   : in    std_logic := 'U';
          TX_FIFO_Full                    : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz       : in    std_logic := 'U';
          TX_FIFO_OVERFLOW_i              : out   std_logic;
          TX_FIFO_OVERFLOW                : out   std_logic;
          TX_FIFO_UNDERRUN_i              : out   std_logic;
          TX_FIFO_UNDERRUN                : out   std_logic
        );
  end component;

  component FIFO_8Kx9_0
    port( ReadFIFO_Write_Ptr        : in    std_logic_vector(1 downto 0) := (others => 'U');
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          RX_FIFO_DOUT_1_0          : out   std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          irx_fifo_rst_i            : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          N_1003                    : in    std_logic := 'U';
          N_657                     : out   std_logic;
          N_658                     : out   std_logic;
          N_659                     : out   std_logic;
          N_661                     : out   std_logic;
          N_717                     : out   std_logic;
          N_663                     : out   std_logic;
          N_662                     : out   std_logic;
          N_660                     : out   std_logic;
          N_1466                    : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9_1
    port( ReadFIFO_Write_Ptr        : in    std_logic_vector(1 downto 0) := (others => 'U');
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          RX_FIFO_DOUT_2_0          : out   std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          irx_fifo_rst_i            : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          N_134                     : in    std_logic := 'U';
          N_664                     : out   std_logic;
          N_665                     : out   std_logic;
          N_666                     : out   std_logic;
          N_668                     : out   std_logic;
          N_670                     : out   std_logic;
          N_716                     : out   std_logic;
          N_669                     : out   std_logic;
          N_667                     : out   std_logic;
          N_1466                    : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_2
    port( ReadFIFO_Write_Ptr        : in    std_logic_vector(1 downto 0) := (others => 'U');
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          RX_FIFO_DOUT_3_0          : out   std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          irx_fifo_rst_i            : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          N_133                     : in    std_logic := 'U';
          N_671                     : out   std_logic;
          N_672                     : out   std_logic;
          N_673                     : out   std_logic;
          N_675                     : out   std_logic;
          N_677                     : out   std_logic;
          N_715                     : out   std_logic;
          N_676                     : out   std_logic;
          N_674                     : out   std_logic;
          N_1466                    : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9
    port( ReadFIFO_Write_Ptr        : in    std_logic_vector(1 downto 0) := (others => 'U');
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          RX_FIFO_DOUT_0_0          : out   std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          irx_fifo_rst_i            : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          N_1004                    : in    std_logic := 'U';
          N_650                     : out   std_logic;
          N_651                     : out   std_logic;
          N_652                     : out   std_logic;
          N_654                     : out   std_logic;
          N_718                     : out   std_logic;
          N_656                     : out   std_logic;
          N_655                     : out   std_logic;
          N_653                     : out   std_logic;
          tx_col_detect_en          : in    std_logic := 'U';
          RX_InProcess_d1           : in    std_logic := 'U';
          sampler_clk1x_en          : in    std_logic := 'U';
          iRX_FIFO_wr_en            : in    std_logic := 'U';
          N_1466                    : out   std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U'
        );
  end component;

    signal itx_fifo_rst_i, \itx_fifo_rst\, irx_fifo_rst_i, 
        \irx_fifo_rst\, \RX_FIFO_UNDERRUN\, \RX_FIFO_OVERFLOW\, 
        \ReadFIFO_Read_Ptr[0]_net_1\, VCC_net_1, N_128_i, 
        GND_net_1, \ReadFIFO_Read_Ptr[1]_net_1\, 
        \ReadFIFO_Read_Ptr_2[1]\, \ReadFIFO_Write_Ptr[0]_net_1\, 
        N_601_i, \ReadFIFO_Write_Ptr[1]_net_1\, N_631_i_i, 
        \iRX_FIFO_UNDERRUN[2]\, \iRX_FIFO_UNDERRUN[3]\, 
        RX_FIFO_UNDERRUN_3_0_0_y0, RX_FIFO_UNDERRUN_3_0_0_co0, 
        \iRX_FIFO_UNDERRUN[0]\, \iRX_FIFO_UNDERRUN[1]\, 
        \iRX_FIFO_Empty[2]\, \iRX_FIFO_Empty[3]\, 
        RX_FIFO_Empty_3_i_m2_0_0_y0, RX_FIFO_Empty_3_i_m2_0_0_co0, 
        \iRX_FIFO_Empty[0]\, \iRX_FIFO_Empty[1]\, 
        \iRX_FIFO_OVERFLOW[2]\, \iRX_FIFO_OVERFLOW[3]\, 
        RX_FIFO_OVERFLOW_3_0_0_y0, RX_FIFO_OVERFLOW_3_0_0_co0, 
        \iRX_FIFO_OVERFLOW[0]\, \iRX_FIFO_OVERFLOW[1]\, N_670, 
        N_677, \RX_FIFO_DOUT_3_0_0_y0[7]\, 
        \RX_FIFO_DOUT_3_0_0_co0[7]\, N_656, N_663, N_716, N_715, 
        \RX_FIFO_DOUT_3_i_m2_i_m2_0_0_y0[8]\, 
        \RX_FIFO_DOUT_3_i_m2_i_m2_0_0_co0[8]\, N_718, N_717, 
        N_669, N_676, \RX_FIFO_DOUT_3_0_0_y0[6]\, 
        \RX_FIFO_DOUT_3_0_0_co0[6]\, N_655, N_662, N_664, N_671, 
        \RX_FIFO_DOUT_3_i_m2_0_0_y0[0]\, 
        \RX_FIFO_DOUT_3_i_m2_0_0_co0[0]\, N_650, N_657, N_668, 
        N_675, \RX_FIFO_DOUT_3_0_0_y0[5]\, 
        \RX_FIFO_DOUT_3_0_0_co0[5]\, N_654, N_661, N_134, N_133, 
        N_1004, N_1003, N_1466 : std_logic;

    for all : FIFO_2Kx8
	Use entity work.FIFO_2Kx8(DEF_ARCH);
    for all : FIFO_8Kx9_0
	Use entity work.FIFO_8Kx9_0(DEF_ARCH);
    for all : FIFO_8Kx9_1
	Use entity work.FIFO_8Kx9_1(DEF_ARCH);
    for all : FIFO_8Kx9_2
	Use entity work.FIFO_8Kx9_2(DEF_ARCH);
    for all : FIFO_8Kx9
	Use entity work.FIFO_8Kx9(DEF_ARCH);
begin 

    ReadFIFO_Read_Ptr(1) <= \ReadFIFO_Read_Ptr[1]_net_1\;
    ReadFIFO_Read_Ptr(0) <= \ReadFIFO_Read_Ptr[0]_net_1\;
    RX_FIFO_OVERFLOW <= \RX_FIFO_OVERFLOW\;
    RX_FIFO_UNDERRUN <= \RX_FIFO_UNDERRUN\;

    \RX_FIFO_DOUT_3_0_0_wmux_0[6]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \RX_FIFO_DOUT_3_0_0_y0[6]\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => N_669, D => N_676, FCI
         => \RX_FIFO_DOUT_3_0_0_co0[6]\, S => OPEN, Y => 
        RX_FIFO_DOUT(6), FCO => OPEN);
    
    irx_fifo_rst_RNIS228 : CLKINT
      port map(A => \irx_fifo_rst\, Y => irx_fifo_rst_i);
    
    \RX_FIFO_DOUT_3_0_0_wmux[6]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => \ReadFIFO_Read_Ptr[0]_net_1\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => N_655, D => N_662, FCI
         => VCC_net_1, S => OPEN, Y => \RX_FIFO_DOUT_3_0_0_y0[6]\, 
        FCO => \RX_FIFO_DOUT_3_0_0_co0[6]\);
    
    \ReadFIFO_Read_Ptr_RNO[1]\ : CFG4
      generic map(INIT => x"B4F0")

      port map(A => up_EOP_sync(1), B => up_EOP_sync(2), C => 
        \ReadFIFO_Read_Ptr[1]_net_1\, D => 
        \ReadFIFO_Read_Ptr[0]_net_1\, Y => 
        \ReadFIFO_Read_Ptr_2[1]\);
    
    RX_FIFO_UNDERRUN_3_0_0_wmux : ARI1
      generic map(INIT => x"0FA44")

      port map(A => \ReadFIFO_Read_Ptr[0]_net_1\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \iRX_FIFO_UNDERRUN[0]\, 
        D => \iRX_FIFO_UNDERRUN[1]\, FCI => VCC_net_1, S => OPEN, 
        Y => RX_FIFO_UNDERRUN_3_0_0_y0, FCO => 
        RX_FIFO_UNDERRUN_3_0_0_co0);
    
    \iRX_FIFO_rd_en_0_o2[0]\ : CFG3
      generic map(INIT => x"04")

      port map(A => \ReadFIFO_Read_Ptr[0]_net_1\, B => 
        RX_FIFO_rd_en, C => \ReadFIFO_Read_Ptr[1]_net_1\, Y => 
        N_1004);
    
    RX_FIFO_OVERFLOW_3_0_0_wmux : ARI1
      generic map(INIT => x"0FA44")

      port map(A => \ReadFIFO_Read_Ptr[0]_net_1\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \iRX_FIFO_OVERFLOW[0]\, 
        D => \iRX_FIFO_OVERFLOW[1]\, FCI => VCC_net_1, S => OPEN, 
        Y => RX_FIFO_OVERFLOW_3_0_0_y0, FCO => 
        RX_FIFO_OVERFLOW_3_0_0_co0);
    
    \RX_FIFO_DOUT_3_0_0_wmux[7]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => \ReadFIFO_Read_Ptr[0]_net_1\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => N_656, D => N_663, FCI
         => VCC_net_1, S => OPEN, Y => \RX_FIFO_DOUT_3_0_0_y0[7]\, 
        FCO => \RX_FIFO_DOUT_3_0_0_co0[7]\);
    
    \ReadFIFO_Read_Ptr_RNO[0]\ : CFG3
      generic map(INIT => x"D2")

      port map(A => up_EOP_sync(2), B => up_EOP_sync(1), C => 
        \ReadFIFO_Read_Ptr[0]_net_1\, Y => N_128_i);
    
    TRANSMIT_FIFO : FIFO_2Kx8
      port map(CoreAPB3_0_APBmslave0_PWDATA(7) => 
        CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), itx_fifo_rst_i => 
        itx_fifo_rst_i, BIT_CLK => BIT_CLK, TX_FIFO_Empty => 
        TX_FIFO_Empty, byte_clk_en => byte_clk_en, N_711 => N_711, 
        N_710 => N_710, N_709 => N_709, N_708 => N_708, N_707 => 
        N_707, N_706 => N_706, N_705 => N_705, N_704 => N_704, 
        TX_PreAmble => TX_PreAmble, TX_DataEn_1_o => 
        TX_DataEn_1_o, un1_tx_packet_length_0_sqmuxa_o => 
        un1_tx_packet_length_0_sqmuxa_o, TX_FIFO_wr_en => 
        TX_FIFO_wr_en, TX_FIFO_Full => TX_FIFO_Full, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz, 
        TX_FIFO_OVERFLOW_i => TX_FIFO_OVERFLOW_i, 
        TX_FIFO_OVERFLOW => TX_FIFO_OVERFLOW, TX_FIFO_UNDERRUN_i
         => TX_FIFO_UNDERRUN_i, TX_FIFO_UNDERRUN => 
        TX_FIFO_UNDERRUN);
    
    \iRX_FIFO_rd_en_0_o2[1]\ : CFG3
      generic map(INIT => x"08")

      port map(A => \ReadFIFO_Read_Ptr[0]_net_1\, B => 
        RX_FIFO_rd_en, C => \ReadFIFO_Read_Ptr[1]_net_1\, Y => 
        N_1003);
    
    RECEIVE_FIFO_1 : FIFO_8Kx9_0
      port map(ReadFIFO_Write_Ptr(1) => 
        \ReadFIFO_Write_Ptr[1]_net_1\, ReadFIFO_Write_Ptr(0) => 
        \ReadFIFO_Write_Ptr[0]_net_1\, RX_FIFO_DIN_pipe(8) => 
        RX_FIFO_DIN_pipe(8), RX_FIFO_DIN_pipe(7) => 
        RX_FIFO_DIN_pipe(7), RX_FIFO_DIN_pipe(6) => 
        RX_FIFO_DIN_pipe(6), RX_FIFO_DIN_pipe(5) => 
        RX_FIFO_DIN_pipe(5), RX_FIFO_DIN_pipe(4) => 
        RX_FIFO_DIN_pipe(4), RX_FIFO_DIN_pipe(3) => 
        RX_FIFO_DIN_pipe(3), RX_FIFO_DIN_pipe(2) => 
        RX_FIFO_DIN_pipe(2), RX_FIFO_DIN_pipe(1) => 
        RX_FIFO_DIN_pipe(1), RX_FIFO_DIN_pipe(0) => 
        RX_FIFO_DIN_pipe(0), RX_FIFO_DOUT_1_0 => RX_FIFO_DOUT_1_0, 
        iRX_FIFO_Empty_0 => \iRX_FIFO_Empty[1]\, 
        iRX_FIFO_UNDERRUN_0 => \iRX_FIFO_UNDERRUN[1]\, 
        iRX_FIFO_Full_0 => iRX_FIFO_Full(1), iRX_FIFO_OVERFLOW_0
         => \iRX_FIFO_OVERFLOW[1]\, irx_fifo_rst_i => 
        irx_fifo_rst_i, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, N_1003 => N_1003, N_657 => 
        N_657, N_658 => N_658, N_659 => N_659, N_661 => N_661, 
        N_717 => N_717, N_663 => N_663, N_662 => N_662, N_660 => 
        N_660, N_1466 => N_1466, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0);
    
    \RX_FIFO_DOUT_3_i_m2_0_0_wmux[0]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => \ReadFIFO_Read_Ptr[0]_net_1\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => N_650, D => N_657, FCI
         => VCC_net_1, S => OPEN, Y => 
        \RX_FIFO_DOUT_3_i_m2_0_0_y0[0]\, FCO => 
        \RX_FIFO_DOUT_3_i_m2_0_0_co0[0]\);
    
    \RX_FIFO_DOUT_3_0_0_wmux_0[5]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \RX_FIFO_DOUT_3_0_0_y0[5]\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => N_668, D => N_675, FCI
         => \RX_FIFO_DOUT_3_0_0_co0[5]\, S => OPEN, Y => 
        RX_FIFO_DOUT(5), FCO => OPEN);
    
    RECEIVE_FIFO_2 : FIFO_8Kx9_1
      port map(ReadFIFO_Write_Ptr(1) => 
        \ReadFIFO_Write_Ptr[1]_net_1\, ReadFIFO_Write_Ptr(0) => 
        \ReadFIFO_Write_Ptr[0]_net_1\, RX_FIFO_DIN_pipe(8) => 
        RX_FIFO_DIN_pipe(8), RX_FIFO_DIN_pipe(7) => 
        RX_FIFO_DIN_pipe(7), RX_FIFO_DIN_pipe(6) => 
        RX_FIFO_DIN_pipe(6), RX_FIFO_DIN_pipe(5) => 
        RX_FIFO_DIN_pipe(5), RX_FIFO_DIN_pipe(4) => 
        RX_FIFO_DIN_pipe(4), RX_FIFO_DIN_pipe(3) => 
        RX_FIFO_DIN_pipe(3), RX_FIFO_DIN_pipe(2) => 
        RX_FIFO_DIN_pipe(2), RX_FIFO_DIN_pipe(1) => 
        RX_FIFO_DIN_pipe(1), RX_FIFO_DIN_pipe(0) => 
        RX_FIFO_DIN_pipe(0), RX_FIFO_DOUT_2_0 => RX_FIFO_DOUT_2_0, 
        iRX_FIFO_Empty_0 => \iRX_FIFO_Empty[2]\, 
        iRX_FIFO_UNDERRUN_0 => \iRX_FIFO_UNDERRUN[2]\, 
        iRX_FIFO_Full_0 => iRX_FIFO_Full(2), iRX_FIFO_OVERFLOW_0
         => \iRX_FIFO_OVERFLOW[2]\, irx_fifo_rst_i => 
        irx_fifo_rst_i, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, N_134 => N_134, N_664 => N_664, 
        N_665 => N_665, N_666 => N_666, N_668 => N_668, N_670 => 
        N_670, N_716 => N_716, N_669 => N_669, N_667 => N_667, 
        N_1466 => N_1466, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    RX_FIFO_Empty_3_i_m2_0_0_wmux_0 : ARI1
      generic map(INIT => x"0F588")

      port map(A => RX_FIFO_Empty_3_i_m2_0_0_y0, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \iRX_FIFO_Empty[2]\, D
         => \iRX_FIFO_Empty[3]\, FCI => 
        RX_FIFO_Empty_3_i_m2_0_0_co0, S => OPEN, Y => N_693, FCO
         => OPEN);
    
    \ReadFIFO_Read_Ptr[0]\ : SLE
      port map(D => N_128_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ReadFIFO_Read_Ptr[0]_net_1\);
    
    itx_fifo_rst_RNIUMSA : CLKINT
      port map(A => \itx_fifo_rst\, Y => itx_fifo_rst_i);
    
    RX_FIFO_UNDERRUN_3_0_0_wmux_0_RNIS837 : CFG1
      generic map(INIT => "01")

      port map(A => \RX_FIFO_UNDERRUN\, Y => RX_FIFO_UNDERRUN_i);
    
    irx_fifo_rst : CFG2
      generic map(INIT => x"1")

      port map(A => un2_apb3_reset, B => RX_FIFO_RST, Y => 
        \irx_fifo_rst\);
    
    \RX_FIFO_DOUT_3_0_0_wmux_0[7]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \RX_FIFO_DOUT_3_0_0_y0[7]\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => N_670, D => N_677, FCI
         => \RX_FIFO_DOUT_3_0_0_co0[7]\, S => OPEN, Y => 
        RX_FIFO_DOUT(7), FCO => OPEN);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \ReadFIFO_Write_Ptr_RNO[1]\ : CFG3
      generic map(INIT => x"78")

      port map(A => \ReadFIFO_Write_Ptr[0]_net_1\, B => 
        rx_packet_complt, C => \ReadFIFO_Write_Ptr[1]_net_1\, Y
         => N_631_i_i);
    
    RX_FIFO_UNDERRUN_3_0_0_wmux_0 : ARI1
      generic map(INIT => x"0F588")

      port map(A => RX_FIFO_UNDERRUN_3_0_0_y0, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \iRX_FIFO_UNDERRUN[2]\, 
        D => \iRX_FIFO_UNDERRUN[3]\, FCI => 
        RX_FIFO_UNDERRUN_3_0_0_co0, S => OPEN, Y => 
        \RX_FIFO_UNDERRUN\, FCO => OPEN);
    
    \ReadFIFO_Write_Ptr[0]\ : SLE
      port map(D => N_601_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ReadFIFO_Write_Ptr[0]_net_1\);
    
    RECEIVE_FIFO_3 : FIFO_8Kx9_2
      port map(ReadFIFO_Write_Ptr(1) => 
        \ReadFIFO_Write_Ptr[1]_net_1\, ReadFIFO_Write_Ptr(0) => 
        \ReadFIFO_Write_Ptr[0]_net_1\, RX_FIFO_DIN_pipe(8) => 
        RX_FIFO_DIN_pipe(8), RX_FIFO_DIN_pipe(7) => 
        RX_FIFO_DIN_pipe(7), RX_FIFO_DIN_pipe(6) => 
        RX_FIFO_DIN_pipe(6), RX_FIFO_DIN_pipe(5) => 
        RX_FIFO_DIN_pipe(5), RX_FIFO_DIN_pipe(4) => 
        RX_FIFO_DIN_pipe(4), RX_FIFO_DIN_pipe(3) => 
        RX_FIFO_DIN_pipe(3), RX_FIFO_DIN_pipe(2) => 
        RX_FIFO_DIN_pipe(2), RX_FIFO_DIN_pipe(1) => 
        RX_FIFO_DIN_pipe(1), RX_FIFO_DIN_pipe(0) => 
        RX_FIFO_DIN_pipe(0), RX_FIFO_DOUT_3_0 => RX_FIFO_DOUT_3_0, 
        iRX_FIFO_Empty_0 => \iRX_FIFO_Empty[3]\, 
        iRX_FIFO_UNDERRUN_0 => \iRX_FIFO_UNDERRUN[3]\, 
        iRX_FIFO_Full_0 => iRX_FIFO_Full(3), iRX_FIFO_OVERFLOW_0
         => \iRX_FIFO_OVERFLOW[3]\, irx_fifo_rst_i => 
        irx_fifo_rst_i, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, N_133 => N_133, N_671 => N_671, 
        N_672 => N_672, N_673 => N_673, N_675 => N_675, N_677 => 
        N_677, N_715 => N_715, N_676 => N_676, N_674 => N_674, 
        N_1466 => N_1466, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0);
    
    \RX_FIFO_DOUT_3_i_m2_i_m2_0_0_wmux[8]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => \ReadFIFO_Read_Ptr[0]_net_1\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => N_718, D => N_717, FCI
         => VCC_net_1, S => OPEN, Y => 
        \RX_FIFO_DOUT_3_i_m2_i_m2_0_0_y0[8]\, FCO => 
        \RX_FIFO_DOUT_3_i_m2_i_m2_0_0_co0[8]\);
    
    RX_FIFO_Empty_3_i_m2_0_0_wmux : ARI1
      generic map(INIT => x"0FA44")

      port map(A => \ReadFIFO_Read_Ptr[0]_net_1\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \iRX_FIFO_Empty[0]\, D
         => \iRX_FIFO_Empty[1]\, FCI => VCC_net_1, S => OPEN, Y
         => RX_FIFO_Empty_3_i_m2_0_0_y0, FCO => 
        RX_FIFO_Empty_3_i_m2_0_0_co0);
    
    \ReadFIFO_Write_Ptr_RNO[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rx_packet_complt, B => 
        \ReadFIFO_Write_Ptr[0]_net_1\, Y => N_601_i);
    
    \RX_FIFO_DOUT_3_i_m2_i_m2_0_0_wmux_0[8]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \RX_FIFO_DOUT_3_i_m2_i_m2_0_0_y0[8]\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => N_716, D => N_715, FCI
         => \RX_FIFO_DOUT_3_i_m2_i_m2_0_0_co0[8]\, S => OPEN, Y
         => N_712, FCO => OPEN);
    
    itx_fifo_rst : CFG2
      generic map(INIT => x"1")

      port map(A => un2_apb3_reset, B => TX_FIFO_RST, Y => 
        \itx_fifo_rst\);
    
    RECEIVE_FIFO_0 : FIFO_8Kx9
      port map(ReadFIFO_Write_Ptr(1) => 
        \ReadFIFO_Write_Ptr[1]_net_1\, ReadFIFO_Write_Ptr(0) => 
        \ReadFIFO_Write_Ptr[0]_net_1\, RX_FIFO_DIN_pipe(8) => 
        RX_FIFO_DIN_pipe(8), RX_FIFO_DIN_pipe(7) => 
        RX_FIFO_DIN_pipe(7), RX_FIFO_DIN_pipe(6) => 
        RX_FIFO_DIN_pipe(6), RX_FIFO_DIN_pipe(5) => 
        RX_FIFO_DIN_pipe(5), RX_FIFO_DIN_pipe(4) => 
        RX_FIFO_DIN_pipe(4), RX_FIFO_DIN_pipe(3) => 
        RX_FIFO_DIN_pipe(3), RX_FIFO_DIN_pipe(2) => 
        RX_FIFO_DIN_pipe(2), RX_FIFO_DIN_pipe(1) => 
        RX_FIFO_DIN_pipe(1), RX_FIFO_DIN_pipe(0) => 
        RX_FIFO_DIN_pipe(0), RX_FIFO_DOUT_0_0 => RX_FIFO_DOUT_0_0, 
        iRX_FIFO_Empty_0 => \iRX_FIFO_Empty[0]\, 
        iRX_FIFO_UNDERRUN_0 => \iRX_FIFO_UNDERRUN[0]\, 
        iRX_FIFO_Full_0 => iRX_FIFO_Full(0), iRX_FIFO_OVERFLOW_0
         => \iRX_FIFO_OVERFLOW[0]\, irx_fifo_rst_i => 
        irx_fifo_rst_i, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, N_1004 => N_1004, N_650 => 
        N_650, N_651 => N_651, N_652 => N_652, N_654 => N_654, 
        N_718 => N_718, N_656 => N_656, N_655 => N_655, N_653 => 
        N_653, tx_col_detect_en => tx_col_detect_en, 
        RX_InProcess_d1 => RX_InProcess_d1, sampler_clk1x_en => 
        sampler_clk1x_en, iRX_FIFO_wr_en => iRX_FIFO_wr_en, 
        N_1466 => N_1466, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0);
    
    \ReadFIFO_Read_Ptr[1]\ : SLE
      port map(D => \ReadFIFO_Read_Ptr_2[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \ReadFIFO_Read_Ptr[1]_net_1\);
    
    \RX_FIFO_DOUT_3_i_m2_0_0_wmux_0[0]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \RX_FIFO_DOUT_3_i_m2_0_0_y0[0]\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => N_664, D => N_671, FCI
         => \RX_FIFO_DOUT_3_i_m2_0_0_co0[0]\, S => OPEN, Y => 
        N_678, FCO => OPEN);
    
    RX_FIFO_OVERFLOW_3_0_0_wmux_0 : ARI1
      generic map(INIT => x"0F588")

      port map(A => RX_FIFO_OVERFLOW_3_0_0_y0, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \iRX_FIFO_OVERFLOW[2]\, 
        D => \iRX_FIFO_OVERFLOW[3]\, FCI => 
        RX_FIFO_OVERFLOW_3_0_0_co0, S => OPEN, Y => 
        \RX_FIFO_OVERFLOW\, FCO => OPEN);
    
    RX_FIFO_OVERFLOW_3_0_0_wmux_0_RNITUE2 : CFG1
      generic map(INIT => "01")

      port map(A => \RX_FIFO_OVERFLOW\, Y => RX_FIFO_OVERFLOW_i);
    
    \RX_FIFO_DOUT_3_0_0_wmux[5]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => \ReadFIFO_Read_Ptr[0]_net_1\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => N_654, D => N_661, FCI
         => VCC_net_1, S => OPEN, Y => \RX_FIFO_DOUT_3_0_0_y0[5]\, 
        FCO => \RX_FIFO_DOUT_3_0_0_co0[5]\);
    
    \ReadFIFO_Write_Ptr[1]\ : SLE
      port map(D => N_631_i_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ReadFIFO_Write_Ptr[1]_net_1\);
    
    \iRX_FIFO_rd_en_0_o2[2]\ : CFG3
      generic map(INIT => x"40")

      port map(A => \ReadFIFO_Read_Ptr[0]_net_1\, B => 
        RX_FIFO_rd_en, C => \ReadFIFO_Read_Ptr[1]_net_1\, Y => 
        N_134);
    
    \iRX_FIFO_rd_en_0_o2[3]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \ReadFIFO_Read_Ptr[0]_net_1\, B => 
        RX_FIFO_rd_en, C => \ReadFIFO_Read_Ptr[1]_net_1\, Y => 
        N_133);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity Interrupts is

    port( CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 1);
          i_int_mask_reg               : in    std_logic_vector(7 downto 1);
          N_799                        : in    std_logic;
          N_789                        : in    std_logic;
          N_790                        : in    std_logic;
          N_791                        : in    std_logic;
          write_reg_en                 : in    std_logic;
          CommsFPGA_top_0_INT          : out   std_logic;
          RX_packet_depth_status       : in    std_logic;
          un2_apb3_reset               : in    std_logic;
          N_385                        : out   std_logic;
          N_384                        : out   std_logic;
          N_381                        : out   std_logic;
          TX_FIFO_UNDERRUN             : in    std_logic;
          un15_int_reg_clr             : out   std_logic;
          tx_FIFO_UNDERRUN_int         : out   std_logic;
          TX_FIFO_UNDERRUN_set         : in    std_logic;
          TX_FIFO_OVERFLOW             : in    std_logic;
          un19_int_reg_clr             : out   std_logic;
          tx_FIFO_OVERFLOW_int         : out   std_logic;
          TX_FIFO_OVERFLOW_set         : in    std_logic;
          RX_FIFO_UNDERRUN             : in    std_logic;
          un23_int_reg_clr             : out   std_logic;
          RX_FIFO_UNDERRUN_set         : in    std_logic;
          RX_FIFO_OVERFLOW             : in    std_logic;
          un27_int_reg_clr             : out   std_logic;
          rx_FIFO_OVERFLOW_int         : out   std_logic;
          RX_FIFO_OVERFLOW_set         : in    std_logic;
          rx_CRC_error                 : in    std_logic;
          un31_int_reg_clr             : out   std_logic;
          rx_CRC_error_int             : out   std_logic;
          rx_CRC_error_set             : in    std_logic;
          iup_EOP                      : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic;
          tx_packet_complt             : in    std_logic;
          CommsFPGA_CCC_0_GL0          : in    std_logic;
          BIT_CLK                      : in    std_logic;
          un2_apb3_reset_i             : in    std_logic;
          un2_apb3_reset_set           : out   std_logic
        );

end Interrupts;

architecture DEF_ARCH of Interrupts is 

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \block_int_until_rd\, block_int_until_rd_i, 
        \tx_packet_complt_toClk16x\, tx_packet_complt_toClk16x_i, 
        GND_net_1, VCC_net_1, \tx_packet_complt_d[7]_net_1\, 
        \tx_packet_complt_d[6]_net_1\, 
        \tx_packet_complt_d[0]_net_1\, 
        \tx_packet_complt_d[1]_net_1\, 
        \tx_packet_complt_d[2]_net_1\, 
        \tx_packet_complt_d[3]_net_1\, 
        \tx_packet_complt_d[4]_net_1\, 
        \tx_packet_complt_d[5]_net_1\, \up_EOP_del[0]_net_1\, 
        \up_EOP_del[1]_net_1\, \up_EOP_del[2]_net_1\, 
        \up_EOP_del[3]_net_1\, \up_EOP_del[4]_net_1\, 
        \up_EOP_del[5]_net_1\, un15_apb3_reset_i, 
        \block_int_until_rd_RNO\, N_61, \irx_packet_avail_int\, 
        rx_CRC_error_intrs, un2_apb3_reset_rs_3, 
        rx_CRC_error_int_net_1, \un31_int_reg_clr\, 
        rx_FIFO_OVERFLOW_intrs, un2_apb3_reset_rs_2, 
        rx_FIFO_OVERFLOW_int_net_1, \un27_int_reg_clr\, 
        rx_FIFO_UNDERRUN_intrs, un2_apb3_reset_rs_1, 
        \rx_FIFO_UNDERRUN_int\, \un23_int_reg_clr\, 
        tx_FIFO_OVERFLOW_intrs, un2_apb3_reset_rs_0, 
        tx_FIFO_OVERFLOW_int_net_1, \un19_int_reg_clr\, 
        tx_FIFO_UNDERRUN_intrs, un2_apb3_reset_rs, 
        tx_FIFO_UNDERRUN_int_net_1, \un15_int_reg_clr\, 
        \tx_packet_complt_toClk16x_set\, tx_packet_complt_intrs, 
        un6_apb3_reset_rs, \tx_packet_complt_int\, 
        un6_apb3_reset_i, un5_int_reg_clr, \N_381\, \N_384\, 
        \N_385\, \INT_2\, \INT_1\, \un1_int_reg_clr_2_i_0_0\, 
        \INT_3\, N_400 : std_logic;

begin 

    N_385 <= \N_385\;
    N_384 <= \N_384\;
    N_381 <= \N_381\;
    un15_int_reg_clr <= \un15_int_reg_clr\;
    tx_FIFO_UNDERRUN_int <= tx_FIFO_UNDERRUN_int_net_1;
    un19_int_reg_clr <= \un19_int_reg_clr\;
    tx_FIFO_OVERFLOW_int <= tx_FIFO_OVERFLOW_int_net_1;
    un23_int_reg_clr <= \un23_int_reg_clr\;
    un27_int_reg_clr <= \un27_int_reg_clr\;
    rx_FIFO_OVERFLOW_int <= rx_FIFO_OVERFLOW_int_net_1;
    un31_int_reg_clr <= \un31_int_reg_clr\;
    rx_CRC_error_int <= rx_CRC_error_int_net_1;

    irx_packet_avail_int_RNIF9DL : CFG2
      generic map(INIT => x"2")

      port map(A => \irx_packet_avail_int\, B => 
        i_int_mask_reg(6), Y => \N_384\);
    
    \TX_PACKET_COMPLETE_INTR.un2_apb3_reset_rs_3\ : SLE
      port map(D => VCC_net_1, CLK => rx_CRC_error, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        un2_apb3_reset_rs_3);
    
    \up_EOP_del[1]\ : SLE
      port map(D => \up_EOP_del[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \up_EOP_del[1]_net_1\);
    
    \TX_PACKET_COMPLETE_INTR.un2_apb3_reset_rs_1_RNIVKP21\ : CFG2
      generic map(INIT => x"2")

      port map(A => \rx_FIFO_UNDERRUN_int\, B => 
        i_int_mask_reg(3), Y => \N_381\);
    
    tx_packet_complt_toClk16x_set_RNO : CFG1
      generic map(INIT => "01")

      port map(A => \tx_packet_complt_toClk16x\, Y => 
        tx_packet_complt_toClk16x_i);
    
    \RX_PACKET_AVAILABLE_INTR.un15_apb3_reset\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \rx_FIFO_UNDERRUN_int\, B => 
        rx_FIFO_OVERFLOW_int_net_1, C => rx_CRC_error_int_net_1, 
        D => un2_apb3_reset, Y => un15_apb3_reset_i);
    
    tx_FIFO_UNDERRUN_int_RNI6GG01 : CFG3
      generic map(INIT => x"EC")

      port map(A => TX_FIFO_UNDERRUN_set, B => 
        tx_FIFO_UNDERRUN_intrs, C => un2_apb3_reset_rs, Y => 
        tx_FIFO_UNDERRUN_int_net_1);
    
    \RX_FIFO_OVERFLOW_INTR.un27_int_reg_clr\ : CFG4
      generic map(INIT => x"8000")

      port map(A => write_reg_en, B => 
        CoreAPB3_0_APBmslave0_PWDATA(2), C => N_790, D => N_799, 
        Y => \un27_int_reg_clr\);
    
    \up_EOP_del[0]\ : SLE
      port map(D => iup_EOP, CLK => m2s010_som_sb_0_CCC_71MHz, EN
         => VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \up_EOP_del[0]_net_1\);
    
    un1_int_reg_clr_2_i_0_0 : CFG4
      generic map(INIT => x"C0E2")

      port map(A => RX_packet_depth_status, B => 
        \block_int_until_rd\, C => \up_EOP_del[5]_net_1\, D => 
        \irx_packet_avail_int\, Y => \un1_int_reg_clr_2_i_0_0\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \up_EOP_del[5]\ : SLE
      port map(D => \up_EOP_del[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \up_EOP_del[5]_net_1\);
    
    irx_packet_avail_int : SLE
      port map(D => block_int_until_rd_i, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_61, ALn => 
        un15_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \irx_packet_avail_int\);
    
    \TX_FIFO_OVERFLOW_INTR.un19_int_reg_clr\ : CFG4
      generic map(INIT => x"8000")

      port map(A => write_reg_en, B => 
        CoreAPB3_0_APBmslave0_PWDATA(4), C => N_790, D => N_799, 
        Y => \un19_int_reg_clr\);
    
    \tx_packet_complt_d[0]\ : SLE
      port map(D => tx_packet_complt, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => un2_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_packet_complt_d[0]_net_1\);
    
    \RX_CRC_ERROR_INTR.un31_int_reg_clr\ : CFG4
      generic map(INIT => x"8000")

      port map(A => write_reg_en, B => 
        CoreAPB3_0_APBmslave0_PWDATA(1), C => N_790, D => N_799, 
        Y => \un31_int_reg_clr\);
    
    \TX_PACKET_COMPLETE_INTR.un5_int_reg_clr\ : CFG4
      generic map(INIT => x"8000")

      port map(A => write_reg_en, B => 
        CoreAPB3_0_APBmslave0_PWDATA(7), C => N_790, D => N_799, 
        Y => un5_int_reg_clr);
    
    \TX_PACKET_COMPLETE_INTR.un2_apb3_reset_rs_2_RNIL9OK\ : CFG3
      generic map(INIT => x"EC")

      port map(A => RX_FIFO_OVERFLOW_set, B => 
        rx_FIFO_OVERFLOW_intrs, C => un2_apb3_reset_rs_2, Y => 
        rx_FIFO_OVERFLOW_int_net_1);
    
    \tx_packet_complt_d[7]\ : SLE
      port map(D => \tx_packet_complt_d[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \tx_packet_complt_d[7]_net_1\);
    
    \TX_PACKET_COMPLETE_INTR.un2_apb3_reset_rs_2\ : SLE
      port map(D => VCC_net_1, CLK => RX_FIFO_OVERFLOW, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        un2_apb3_reset_rs_2);
    
    \tx_FIFO_OVERFLOW_int\ : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \un19_int_reg_clr\, ALn => un2_apb3_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => tx_FIFO_OVERFLOW_intrs);
    
    \rx_CRC_error_int\ : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \un31_int_reg_clr\, ALn => un2_apb3_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => rx_CRC_error_intrs);
    
    \TX_PACKET_COMPLETE_INTR.un2_apb3_reset_rs\ : SLE
      port map(D => VCC_net_1, CLK => TX_FIFO_UNDERRUN, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        un2_apb3_reset_rs);
    
    \tx_FIFO_UNDERRUN_int\ : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \un15_int_reg_clr\, ALn => un2_apb3_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => tx_FIFO_UNDERRUN_intrs);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \tx_packet_complt_d[5]\ : SLE
      port map(D => \tx_packet_complt_d[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \tx_packet_complt_d[5]_net_1\);
    
    \tx_packet_complt_d[4]\ : SLE
      port map(D => \tx_packet_complt_d[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \tx_packet_complt_d[4]_net_1\);
    
    \TX_PACKET_COMPLETE_INTR.un2_apb3_reset_rs_1_RNIIFJR\ : CFG3
      generic map(INIT => x"EC")

      port map(A => RX_FIFO_UNDERRUN_set, B => 
        rx_FIFO_UNDERRUN_intrs, C => un2_apb3_reset_rs_1, Y => 
        \rx_FIFO_UNDERRUN_int\);
    
    \tx_packet_complt_d[3]\ : SLE
      port map(D => \tx_packet_complt_d[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \tx_packet_complt_d[3]_net_1\);
    
    \TX_PACKET_COMPLETE_INTR.un2_apb3_reset_rs_3_RNIA45O\ : CFG3
      generic map(INIT => x"EC")

      port map(A => rx_CRC_error_set, B => rx_CRC_error_intrs, C
         => un2_apb3_reset_rs_3, Y => rx_CRC_error_int_net_1);
    
    INT_3 : CFG4
      generic map(INIT => x"FBFA")

      port map(A => \N_384\, B => i_int_mask_reg(5), C => \N_385\, 
        D => tx_FIFO_UNDERRUN_int_net_1, Y => \INT_3\);
    
    tx_packet_complt_int : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => un5_int_reg_clr, ALn => un6_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => tx_packet_complt_intrs);
    
    irx_packet_avail_int_RNO : CFG1
      generic map(INIT => "01")

      port map(A => \block_int_until_rd\, Y => 
        block_int_until_rd_i);
    
    \tx_packet_complt_d[6]\ : SLE
      port map(D => \tx_packet_complt_d[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \tx_packet_complt_d[6]_net_1\);
    
    block_int_until_rd : SLE
      port map(D => \block_int_until_rd_RNO\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_61, ALn => 
        un15_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \block_int_until_rd\);
    
    \TX_PACKET_COMPLETE_INTR.un2_apb3_reset_rs_0\ : SLE
      port map(D => VCC_net_1, CLK => TX_FIFO_OVERFLOW, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        un2_apb3_reset_rs_0);
    
    un1_int_reg_clr_2_i_0 : CFG4
      generic map(INIT => x"EAAA")

      port map(A => \un1_int_reg_clr_2_i_0_0\, B => 
        \block_int_until_rd\, C => N_400, D => 
        CoreAPB3_0_APBmslave0_PWDATA(6), Y => N_61);
    
    tx_packet_complt_toClk16x : CFG2
      generic map(INIT => x"2")

      port map(A => \tx_packet_complt_d[6]_net_1\, B => 
        \tx_packet_complt_d[7]_net_1\, Y => 
        \tx_packet_complt_toClk16x\);
    
    \TX_FIFO_UNDERRUN_INTR.un15_int_reg_clr\ : CFG4
      generic map(INIT => x"8000")

      port map(A => write_reg_en, B => 
        CoreAPB3_0_APBmslave0_PWDATA(5), C => N_790, D => N_799, 
        Y => \un15_int_reg_clr\);
    
    INT_1 : CFG4
      generic map(INIT => x"7350")

      port map(A => i_int_mask_reg(2), B => i_int_mask_reg(1), C
         => rx_FIFO_OVERFLOW_int_net_1, D => 
        rx_CRC_error_int_net_1, Y => \INT_1\);
    
    \RX_FIFO_UNDERRUN_INTR.un23_int_reg_clr\ : CFG4
      generic map(INIT => x"8000")

      port map(A => write_reg_en, B => 
        CoreAPB3_0_APBmslave0_PWDATA(3), C => N_790, D => N_799, 
        Y => \un23_int_reg_clr\);
    
    \rx_FIFO_OVERFLOW_int\ : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \un27_int_reg_clr\, ALn => un2_apb3_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => rx_FIFO_OVERFLOW_intrs);
    
    \TX_PACKET_COMPLETE_INTR.un2_apb3_reset_set\ : SLE
      port map(D => GND_net_1, CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => un2_apb3_reset_i, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        un2_apb3_reset_set);
    
    \up_EOP_del[4]\ : SLE
      port map(D => \up_EOP_del[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \up_EOP_del[4]_net_1\);
    
    \tx_packet_complt_d[1]\ : SLE
      port map(D => \tx_packet_complt_d[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \tx_packet_complt_d[1]_net_1\);
    
    INT_2 : CFG3
      generic map(INIT => x"BA")

      port map(A => \N_381\, B => i_int_mask_reg(4), C => 
        tx_FIFO_OVERFLOW_int_net_1, Y => \INT_2\);
    
    \tx_packet_complt_d[2]\ : SLE
      port map(D => \tx_packet_complt_d[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \tx_packet_complt_d[2]_net_1\);
    
    block_int_until_rd_RNO : CFG3
      generic map(INIT => x"B3")

      port map(A => N_400, B => \block_int_until_rd\, C => 
        CoreAPB3_0_APBmslave0_PWDATA(6), Y => 
        \block_int_until_rd_RNO\);
    
    tx_packet_complt_toClk16x_set_RNI9HQV : CFG2
      generic map(INIT => x"2")

      port map(A => \tx_packet_complt_int\, B => 
        i_int_mask_reg(7), Y => \N_385\);
    
    \TX_PACKET_COMPLETE_INTR.un6_apb3_reset\ : CFG2
      generic map(INIT => x"1")

      port map(A => un2_apb3_reset, B => 
        tx_FIFO_UNDERRUN_int_net_1, Y => un6_apb3_reset_i);
    
    \TX_PACKET_COMPLETE_INTR.un6_apb3_reset_rs\ : SLE
      port map(D => VCC_net_1, CLK => \tx_packet_complt_toClk16x\, 
        EN => VCC_net_1, ALn => un6_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        VCC_net_1, Q => un6_apb3_reset_rs);
    
    \TX_PACKET_COMPLETE_INTR.un2_apb3_reset_rs_1\ : SLE
      port map(D => VCC_net_1, CLK => RX_FIFO_UNDERRUN, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        un2_apb3_reset_rs_1);
    
    \TX_PACKET_COMPLETE_INTR.un2_apb3_reset_rs_0_RNINL6E\ : CFG3
      generic map(INIT => x"EC")

      port map(A => TX_FIFO_OVERFLOW_set, B => 
        tx_FIFO_OVERFLOW_intrs, C => un2_apb3_reset_rs_0, Y => 
        tx_FIFO_OVERFLOW_int_net_1);
    
    INT : CFG3
      generic map(INIT => x"FE")

      port map(A => \INT_1\, B => \INT_2\, C => \INT_3\, Y => 
        CommsFPGA_top_0_INT);
    
    \REGISTER_CLEAR_INST.un1_write_reg_en_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => write_reg_en, B => N_791, C => N_790, D => 
        N_789, Y => N_400);
    
    \up_EOP_del[3]\ : SLE
      port map(D => \up_EOP_del[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \up_EOP_del[3]_net_1\);
    
    \up_EOP_del[2]\ : SLE
      port map(D => \up_EOP_del[1]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \up_EOP_del[2]_net_1\);
    
    tx_packet_complt_toClk16x_set : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => un5_int_reg_clr, ALn => tx_packet_complt_toClk16x_i, 
        ADn => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \tx_packet_complt_toClk16x_set\);
    
    tx_packet_complt_toClk16x_set_RNIO7KO : CFG3
      generic map(INIT => x"EC")

      port map(A => \tx_packet_complt_toClk16x_set\, B => 
        tx_packet_complt_intrs, C => un6_apb3_reset_rs, Y => 
        \tx_packet_complt_int\);
    
    rx_FIFO_UNDERRUN_int : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \un23_int_reg_clr\, ALn => un2_apb3_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => rx_FIFO_UNDERRUN_intrs);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity uP_if is

    port( RX_FIFO_DIN                        : in    std_logic_vector(3 downto 2);
          rx_crc_data_calc                   : in    std_logic_vector(11 downto 10);
          CoreAPB3_0_APBmslave0_PADDR        : in    std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PRDATA_m     : out   std_logic_vector(7 downto 0);
          RX_FIFO_DOUT                       : in    std_logic_vector(7 downto 5);
          iRX_FIFO_Full                      : in    std_logic_vector(3 downto 0);
          ReadFIFO_Read_Ptr                  : in    std_logic_vector(1 downto 0);
          consumer_type4_reg                 : out   std_logic_vector(9 downto 0);
          consumer_type3_reg                 : out   std_logic_vector(9 downto 0);
          consumer_type2_reg                 : out   std_logic_vector(9 downto 0);
          consumer_type1_reg                 : out   std_logic_vector(9 downto 0);
          CoreAPB3_0_APBmslave0_PWDATA       : in    std_logic_vector(7 downto 0);
          up_EOP_sync                        : out   std_logic_vector(2 downto 1);
          lfsr_c_i_i_0                       : out   std_logic;
          RX_FIFO_DIN_pipe_0                 : in    std_logic;
          RX_FIFO_DOUT_1_0                   : in    std_logic;
          RX_FIFO_DOUT_0_0                   : in    std_logic;
          RX_FIFO_DOUT_3_0                   : in    std_logic;
          RX_FIFO_DOUT_2_0                   : in    std_logic;
          un2_apb3_reset_set                 : out   std_logic;
          un2_apb3_reset_i                   : in    std_logic;
          BIT_CLK                            : in    std_logic;
          tx_packet_complt                   : in    std_logic;
          rx_CRC_error_set                   : in    std_logic;
          un31_int_reg_clr                   : out   std_logic;
          rx_CRC_error                       : in    std_logic;
          RX_FIFO_OVERFLOW_set               : in    std_logic;
          un27_int_reg_clr                   : out   std_logic;
          RX_FIFO_OVERFLOW                   : in    std_logic;
          RX_FIFO_UNDERRUN_set               : in    std_logic;
          un23_int_reg_clr                   : out   std_logic;
          RX_FIFO_UNDERRUN                   : in    std_logic;
          TX_FIFO_OVERFLOW_set               : in    std_logic;
          un19_int_reg_clr                   : out   std_logic;
          TX_FIFO_OVERFLOW                   : in    std_logic;
          TX_FIFO_UNDERRUN_set               : in    std_logic;
          un15_int_reg_clr                   : out   std_logic;
          TX_FIFO_UNDERRUN                   : in    std_logic;
          un2_apb3_reset                     : in    std_logic;
          CommsFPGA_top_0_INT                : out   std_logic;
          TX_PreAmble                        : in    std_logic;
          N_712                              : in    std_logic;
          N_855_i                            : out   std_logic;
          CoreAPB3_0_APBmslave0_PWRITE       : in    std_logic;
          N_993_i                            : out   std_logic;
          sampler_clk1x_en                   : in    std_logic;
          SM_advance_i                       : in    std_logic;
          N_41_i                             : out   std_logic;
          rx_crc_HighByte_en                 : in    std_logic;
          N_535                              : in    std_logic;
          CoreAPB3_0_APBmslave0_PREADY_i_m_i : out   std_logic;
          CoreAPB3_0_APBmslave0_PENABLE      : in    std_logic;
          RX_FIFO_RST_1                      : out   std_logic;
          RX_EarlyTerm                       : in    std_logic;
          CoreAPB3_0_APBmslave0_PSELx        : in    std_logic;
          TX_FIFO_Empty                      : in    std_logic;
          TX_FIFO_Full                       : in    std_logic;
          N_693                              : in    std_logic;
          N_678                              : in    std_logic;
          N_658                              : in    std_logic;
          N_651                              : in    std_logic;
          N_672                              : in    std_logic;
          N_665                              : in    std_logic;
          N_659                              : in    std_logic;
          N_652                              : in    std_logic;
          N_673                              : in    std_logic;
          N_666                              : in    std_logic;
          N_660                              : in    std_logic;
          N_653                              : in    std_logic;
          N_674                              : in    std_logic;
          N_667                              : in    std_logic;
          rx_packet_complt                   : in    std_logic;
          RX_FIFO_rd_en                      : out   std_logic;
          TX_FIFO_wr_en                      : out   std_logic;
          N_855_i_i                          : in    std_logic;
          TX_FIFO_RST                        : out   std_logic;
          start_tx_FIFO                      : out   std_logic;
          internal_loopback                  : out   std_logic;
          external_loopback                  : out   std_logic;
          long_reset                         : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz          : in    std_logic;
          long_reset_set                     : in    std_logic;
          CommsFPGA_CCC_0_GL0                : in    std_logic;
          long_reset_i                       : in    std_logic
        );

end uP_if;

architecture DEF_ARCH of uP_if is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component Interrupts
    port( CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 1) := (others => 'U');
          i_int_mask_reg               : in    std_logic_vector(7 downto 1) := (others => 'U');
          N_799                        : in    std_logic := 'U';
          N_789                        : in    std_logic := 'U';
          N_790                        : in    std_logic := 'U';
          N_791                        : in    std_logic := 'U';
          write_reg_en                 : in    std_logic := 'U';
          CommsFPGA_top_0_INT          : out   std_logic;
          RX_packet_depth_status       : in    std_logic := 'U';
          un2_apb3_reset               : in    std_logic := 'U';
          N_385                        : out   std_logic;
          N_384                        : out   std_logic;
          N_381                        : out   std_logic;
          TX_FIFO_UNDERRUN             : in    std_logic := 'U';
          un15_int_reg_clr             : out   std_logic;
          tx_FIFO_UNDERRUN_int         : out   std_logic;
          TX_FIFO_UNDERRUN_set         : in    std_logic := 'U';
          TX_FIFO_OVERFLOW             : in    std_logic := 'U';
          un19_int_reg_clr             : out   std_logic;
          tx_FIFO_OVERFLOW_int         : out   std_logic;
          TX_FIFO_OVERFLOW_set         : in    std_logic := 'U';
          RX_FIFO_UNDERRUN             : in    std_logic := 'U';
          un23_int_reg_clr             : out   std_logic;
          RX_FIFO_UNDERRUN_set         : in    std_logic := 'U';
          RX_FIFO_OVERFLOW             : in    std_logic := 'U';
          un27_int_reg_clr             : out   std_logic;
          rx_FIFO_OVERFLOW_int         : out   std_logic;
          RX_FIFO_OVERFLOW_set         : in    std_logic := 'U';
          rx_CRC_error                 : in    std_logic := 'U';
          un31_int_reg_clr             : out   std_logic;
          rx_CRC_error_int             : out   std_logic;
          rx_CRC_error_set             : in    std_logic := 'U';
          iup_EOP                      : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic := 'U';
          tx_packet_complt             : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0          : in    std_logic := 'U';
          BIT_CLK                      : in    std_logic := 'U';
          un2_apb3_reset_i             : in    std_logic := 'U';
          un2_apb3_reset_set           : out   std_logic
        );
  end component;

    signal \iAPB3_READY[0]_net_1\, \iAPB3_READY_i[0]\, 
        \up_EOP_sync[0]_net_1\, VCC_net_1, \iup_EOP\, GND_net_1, 
        \up_EOP_sync[1]_net_1\, \up_EOP_sync[2]_net_1\, 
        \iAPB3_READYrs[0]\, un5_apb3_rst_rs, un5_apb3_rst_i, 
        CoreAPB3_0_APBmslave0_PREADYrs, 
        CoreAPB3_0_APBmslave0_PREADY, \mac_3_byte_4_reg[7]_net_1\, 
        un13_mac_3_byte_4_reg_en, \mac_3_byte_3_reg[0]_net_1\, 
        un13_mac_3_byte_3_reg_en, \mac_3_byte_3_reg[1]_net_1\, 
        \mac_3_byte_3_reg[2]_net_1\, \mac_3_byte_3_reg[3]_net_1\, 
        \mac_3_byte_3_reg[4]_net_1\, \mac_3_byte_3_reg[5]_net_1\, 
        \mac_3_byte_3_reg[6]_net_1\, \mac_3_byte_3_reg[7]_net_1\, 
        \mac_3_byte_5_reg[0]_net_1\, un13_mac_3_byte_5_reg_en, 
        \mac_3_byte_5_reg[1]_net_1\, \mac_3_byte_5_reg[2]_net_1\, 
        \mac_3_byte_5_reg[3]_net_1\, \mac_3_byte_5_reg[4]_net_1\, 
        \mac_3_byte_5_reg[5]_net_1\, \mac_3_byte_5_reg[6]_net_1\, 
        \mac_3_byte_5_reg[7]_net_1\, \mac_3_byte_4_reg[0]_net_1\, 
        \mac_3_byte_4_reg[1]_net_1\, \mac_3_byte_4_reg[2]_net_1\, 
        \mac_3_byte_4_reg[3]_net_1\, \mac_3_byte_4_reg[4]_net_1\, 
        \mac_3_byte_4_reg[5]_net_1\, \mac_3_byte_4_reg[6]_net_1\, 
        \mac_4_byte_1_reg[1]_net_1\, un13_mac_4_byte_1_reg_en, 
        \mac_4_byte_1_reg[2]_net_1\, \mac_4_byte_1_reg[3]_net_1\, 
        \mac_4_byte_1_reg[4]_net_1\, \mac_4_byte_1_reg[5]_net_1\, 
        \mac_4_byte_1_reg[6]_net_1\, \mac_4_byte_1_reg[7]_net_1\, 
        \mac_3_byte_6_reg[0]_net_1\, un13_mac_3_byte_6_reg_en, 
        \mac_3_byte_6_reg[1]_net_1\, \mac_3_byte_6_reg[2]_net_1\, 
        \mac_3_byte_6_reg[3]_net_1\, \mac_3_byte_6_reg[4]_net_1\, 
        \mac_3_byte_6_reg[5]_net_1\, \mac_3_byte_6_reg[6]_net_1\, 
        \mac_3_byte_6_reg[7]_net_1\, \mac_4_byte_3_reg[2]_net_1\, 
        un13_mac_4_byte_3_reg_en, \mac_4_byte_3_reg[3]_net_1\, 
        \mac_4_byte_3_reg[4]_net_1\, \mac_4_byte_3_reg[5]_net_1\, 
        \mac_4_byte_3_reg[6]_net_1\, \mac_4_byte_3_reg[7]_net_1\, 
        \mac_4_byte_2_reg[0]_net_1\, un13_mac_4_byte_2_reg_en, 
        \mac_4_byte_2_reg[1]_net_1\, \mac_4_byte_2_reg[2]_net_1\, 
        \mac_4_byte_2_reg[3]_net_1\, \mac_4_byte_2_reg[4]_net_1\, 
        \mac_4_byte_2_reg[5]_net_1\, \mac_4_byte_2_reg[6]_net_1\, 
        \mac_4_byte_2_reg[7]_net_1\, \mac_4_byte_1_reg[0]_net_1\, 
        \mac_4_byte_5_reg[3]_net_1\, un13_mac_4_byte_5_reg_en, 
        \mac_4_byte_5_reg[4]_net_1\, \mac_4_byte_5_reg[5]_net_1\, 
        \mac_4_byte_5_reg[6]_net_1\, \mac_4_byte_5_reg[7]_net_1\, 
        \mac_4_byte_4_reg[0]_net_1\, un13_mac_4_byte_4_reg_en, 
        \mac_4_byte_4_reg[1]_net_1\, \mac_4_byte_4_reg[2]_net_1\, 
        \mac_4_byte_4_reg[3]_net_1\, \mac_4_byte_4_reg[4]_net_1\, 
        \mac_4_byte_4_reg[5]_net_1\, \mac_4_byte_4_reg[6]_net_1\, 
        \mac_4_byte_4_reg[7]_net_1\, \mac_4_byte_3_reg[0]_net_1\, 
        \mac_4_byte_3_reg[1]_net_1\, \mac_1_byte_1_reg[4]_net_1\, 
        un13_mac_1_byte_1_reg_en, \mac_1_byte_1_reg[5]_net_1\, 
        \mac_1_byte_1_reg[6]_net_1\, \mac_1_byte_1_reg[7]_net_1\, 
        \i_int_mask_reg[0]_net_1\, N_1354_i, 
        \i_int_mask_reg[1]_net_1\, \i_int_mask_reg[2]_net_1\, 
        \i_int_mask_reg[3]_net_1\, \i_int_mask_reg[4]_net_1\, 
        \i_int_mask_reg[5]_net_1\, \i_int_mask_reg[6]_net_1\, 
        \i_int_mask_reg[7]_net_1\, \mac_4_byte_5_reg[0]_net_1\, 
        \mac_4_byte_5_reg[1]_net_1\, \mac_4_byte_5_reg[2]_net_1\, 
        \mac_1_byte_3_reg[5]_net_1\, un13_mac_1_byte_3_reg_en, 
        \mac_1_byte_3_reg[6]_net_1\, \mac_1_byte_3_reg[7]_net_1\, 
        \consumer_type1_reg[0]\, un13_mac_1_byte_2_reg_en, 
        \consumer_type1_reg[1]\, \consumer_type1_reg[2]\, 
        \consumer_type1_reg[3]\, \consumer_type1_reg[4]\, 
        \consumer_type1_reg[5]\, \consumer_type1_reg[6]\, 
        \consumer_type1_reg[7]\, \consumer_type1_reg[8]\, 
        \consumer_type1_reg[9]\, \mac_1_byte_1_reg[2]_net_1\, 
        \mac_1_byte_1_reg[3]_net_1\, \mac_1_byte_5_reg[6]_net_1\, 
        un13_mac_1_byte_5_reg_en, \mac_1_byte_5_reg[7]_net_1\, 
        \consumer_type2_reg[0]\, un13_mac_1_byte_4_reg_en, 
        \consumer_type2_reg[1]\, \consumer_type2_reg[2]\, 
        \consumer_type2_reg[3]\, \consumer_type2_reg[4]\, 
        \consumer_type2_reg[5]\, \consumer_type2_reg[6]\, 
        \consumer_type2_reg[7]\, \consumer_type2_reg[8]\, 
        \consumer_type2_reg[9]\, \mac_1_byte_3_reg[2]_net_1\, 
        \mac_1_byte_3_reg[3]_net_1\, \mac_1_byte_3_reg[4]_net_1\, 
        \mac_2_byte_1_reg[7]_net_1\, un13_mac_2_byte_1_reg_en, 
        \consumer_type3_reg[0]\, un13_mac_1_byte_6_reg_en, 
        \consumer_type3_reg[1]\, \consumer_type3_reg[2]\, 
        \consumer_type3_reg[3]\, \consumer_type3_reg[4]\, 
        \consumer_type3_reg[5]\, \consumer_type3_reg[6]\, 
        \consumer_type3_reg[7]\, \consumer_type3_reg[8]\, 
        \consumer_type3_reg[9]\, \mac_1_byte_5_reg[2]_net_1\, 
        \mac_1_byte_5_reg[3]_net_1\, \mac_1_byte_5_reg[4]_net_1\, 
        \mac_1_byte_5_reg[5]_net_1\, \consumer_type4_reg[0]\, 
        un13_mac_2_byte_2_reg_en, \consumer_type4_reg[1]\, 
        \consumer_type4_reg[2]\, \consumer_type4_reg[3]\, 
        \consumer_type4_reg[4]\, \consumer_type4_reg[5]\, 
        \consumer_type4_reg[6]\, \consumer_type4_reg[7]\, 
        \consumer_type4_reg[8]\, \consumer_type4_reg[9]\, 
        \mac_2_byte_1_reg[2]_net_1\, \mac_2_byte_1_reg[3]_net_1\, 
        \mac_2_byte_1_reg[4]_net_1\, \mac_2_byte_1_reg[5]_net_1\, 
        \mac_2_byte_1_reg[6]_net_1\, \mac_2_byte_4_reg[1]_net_1\, 
        un13_mac_2_byte_4_reg_en, \mac_2_byte_4_reg[2]_net_1\, 
        \mac_2_byte_4_reg[3]_net_1\, \mac_2_byte_4_reg[4]_net_1\, 
        \mac_2_byte_4_reg[5]_net_1\, \mac_2_byte_4_reg[6]_net_1\, 
        \mac_2_byte_4_reg[7]_net_1\, \mac_2_byte_3_reg[0]_net_1\, 
        un13_mac_2_byte_3_reg_en, \mac_2_byte_3_reg[1]_net_1\, 
        \mac_2_byte_3_reg[2]_net_1\, \mac_2_byte_3_reg[3]_net_1\, 
        \mac_2_byte_3_reg[4]_net_1\, \mac_2_byte_3_reg[5]_net_1\, 
        \mac_2_byte_3_reg[6]_net_1\, \mac_2_byte_3_reg[7]_net_1\, 
        \mac_2_byte_6_reg[2]_net_1\, un13_mac_2_byte_6_reg_en, 
        \mac_2_byte_6_reg[3]_net_1\, \mac_2_byte_6_reg[4]_net_1\, 
        \mac_2_byte_6_reg[5]_net_1\, \mac_2_byte_6_reg[6]_net_1\, 
        \mac_2_byte_6_reg[7]_net_1\, \mac_2_byte_5_reg[0]_net_1\, 
        un13_mac_2_byte_5_reg_en, \mac_2_byte_5_reg[1]_net_1\, 
        \mac_2_byte_5_reg[2]_net_1\, \mac_2_byte_5_reg[3]_net_1\, 
        \mac_2_byte_5_reg[4]_net_1\, \mac_2_byte_5_reg[5]_net_1\, 
        \mac_2_byte_5_reg[6]_net_1\, \mac_2_byte_5_reg[7]_net_1\, 
        \mac_2_byte_4_reg[0]_net_1\, \mac_3_byte_2_reg[3]_net_1\, 
        un13_mac_3_byte_2_reg_en, \mac_3_byte_2_reg[4]_net_1\, 
        \mac_3_byte_2_reg[5]_net_1\, \mac_3_byte_2_reg[6]_net_1\, 
        \mac_3_byte_2_reg[7]_net_1\, \mac_3_byte_1_reg[0]_net_1\, 
        un13_mac_3_byte_1_reg_en, \mac_3_byte_1_reg[1]_net_1\, 
        \mac_3_byte_1_reg[2]_net_1\, \mac_3_byte_1_reg[3]_net_1\, 
        \mac_3_byte_1_reg[4]_net_1\, \mac_3_byte_1_reg[5]_net_1\, 
        \mac_3_byte_1_reg[6]_net_1\, \mac_3_byte_1_reg[7]_net_1\, 
        \mac_2_byte_6_reg[0]_net_1\, \mac_2_byte_6_reg[1]_net_1\, 
        \mac_4_byte_6_reg[4]_net_1\, un13_mac_4_byte_6_reg_en, 
        \mac_4_byte_6_reg[5]_net_1\, \mac_4_byte_6_reg[6]_net_1\, 
        \mac_4_byte_6_reg[7]_net_1\, \control_reg[0]_net_1\, 
        control_reg_13, \external_loopback\, 
        \control_reg[2]_net_1\, \control_reg[3]_net_1\, 
        \internal_loopback\, \start_tx_FIFO\, \control_reg_3[5]\, 
        un1_control_reg_en_2_i_0, rx_FIFO_rst_reg, \TX_FIFO_RST\, 
        \mac_3_byte_2_reg[0]_net_1\, \mac_3_byte_2_reg[1]_net_1\, 
        \mac_3_byte_2_reg[2]_net_1\, \scratch_pad_reg[0]_net_1\, 
        \write_scratch_reg_en\, \scratch_pad_reg[1]_net_1\, 
        \scratch_pad_reg[2]_net_1\, \scratch_pad_reg[3]_net_1\, 
        \scratch_pad_reg[4]_net_1\, \scratch_pad_reg[5]_net_1\, 
        \scratch_pad_reg[6]_net_1\, \scratch_pad_reg[7]_net_1\, 
        \mac_4_byte_6_reg[0]_net_1\, \mac_4_byte_6_reg[1]_net_1\, 
        \mac_4_byte_6_reg[2]_net_1\, \mac_4_byte_6_reg[3]_net_1\, 
        \mac_4_byte_5_reg_en\, mac_4_byte_6_reg_en_1, N_357, 
        \mac_4_byte_4_reg_en\, N_356, \mac_4_byte_3_reg_en\, 
        N_355, un1_apb3_addr, N_854_i_i, N_330, 
        \mac_3_byte_2_reg_en\, N_348, \mac_3_byte_1_reg_en\, 
        N_347, \mac_2_byte_6_reg_en\, N_346, 
        \mac_2_byte_5_reg_en\, N_345, \mac_2_byte_4_reg_en\, 
        N_344, \mac_2_byte_3_reg_en\, N_343, 
        \mac_2_byte_2_reg_en\, N_342, \mac_3_byte_3_reg_en\, 
        N_349, \mac_3_byte_4_reg_en\, N_350, 
        \mac_3_byte_5_reg_en\, N_351, \mac_3_byte_6_reg_en\, 
        N_352, \mac_4_byte_1_reg_en\, N_353, 
        \mac_4_byte_2_reg_en\, N_354, \mac_4_byte_6_reg_en\, 
        N_358, N_743, N_734, N_742, N_733, \mac_1_byte_2_reg_en\, 
        N_336, \control_reg_en\, N_331, \mac_1_byte_4_reg_en\, 
        N_338, \mac_1_byte_6_reg_en\, N_340, \int_mask_reg_en\, 
        N_333, \mac_1_byte_5_reg_en\, N_339, 
        \mac_1_byte_1_reg_en\, N_335, N_329, 
        \mac_2_byte_1_reg_en\, N_341, \mac_1_byte_3_reg_en\, 
        N_337, \write_reg_en\, \read_reg_en\, un117_apb3_addr, 
        \RX_packet_depth_status\, rx_packet_depth_status2, 
        \CoreAPB3_0_APBmslave0_PRDATA[2]\, N_41_mux, 
        \APB3_RDATA_1[2]\, \CoreAPB3_0_APBmslave0_PRDATA[3]\, 
        \APB3_RDATA_1[3]\, \CoreAPB3_0_APBmslave0_PRDATA[4]\, 
        \APB3_RDATA_1[4]\, \CoreAPB3_0_APBmslave0_PRDATA[5]\, 
        \APB3_RDATA_1[5]_net_1\, 
        \CoreAPB3_0_APBmslave0_PRDATA[6]\, 
        \APB3_RDATA_1[6]_net_1\, 
        \CoreAPB3_0_APBmslave0_PRDATA[7]\, \APB3_RDATA_1[7]\, 
        \CoreAPB3_0_APBmslave0_PRDATA[0]\, \APB3_RDATA_1[0]\, 
        \CoreAPB3_0_APBmslave0_PRDATA[1]\, \APB3_RDATA_1[1]\, 
        \RX_packet_depth[0]_net_1\, \RX_packet_depth_s[0]\, 
        N_127_i, \RX_packet_depth[1]_net_1\, 
        \RX_packet_depth_s[1]\, \RX_packet_depth[2]_net_1\, 
        \RX_packet_depth_s[2]\, \RX_packet_depth[3]_net_1\, 
        \RX_packet_depth_s[3]\, \RX_packet_depth[4]_net_1\, 
        \RX_packet_depth_s[4]\, \RX_packet_depth[5]_net_1\, 
        \RX_packet_depth_s[5]\, \RX_packet_depth[6]_net_1\, 
        \RX_packet_depth_s[6]\, \RX_packet_depth[7]_net_1\, 
        \RX_packet_depth_s[7]_net_1\, 
        un12_mac_2_byte_1_reg_en_16_0_reto, 
        un12_mac_2_byte_1_reg_en_16_0, 
        un12_mac_2_byte_1_reg_en_16_1_reto, 
        un12_mac_2_byte_1_reg_en_16_1, 
        un12_mac_2_byte_1_reg_en_16_2_reto, 
        un12_mac_2_byte_1_reg_en_16_2, N_6_reto, N_6, N_335_reto, 
        N_733_reto, mac_4_byte_6_reg_en_1_reto, 
        mac_1_byte_1_reg_en_reto, RX_packet_depth_s_390_FCO, 
        \RX_packet_depth_cry[0]_net_1\, 
        \RX_packet_depth_cry[1]_net_1\, 
        \RX_packet_depth_cry[2]_net_1\, 
        \RX_packet_depth_cry[3]_net_1\, 
        \RX_packet_depth_cry[4]_net_1\, 
        \RX_packet_depth_cry[5]_net_1\, 
        \RX_packet_depth_cry[6]_net_1\, 
        \APB3_RDATA_1_25_0_wmux_0_Y[7]\, 
        \APB3_RDATA_1_25_0_0_y0[7]\, \APB3_RDATA_1_25_0_0_co0[7]\, 
        \APB3_RDATA_1_25_0_wmux_0_Y[5]\, 
        \APB3_RDATA_1_25_0_0_y0[5]\, \APB3_RDATA_1_25_0_0_co0[5]\, 
        \APB3_RDATA_1_25_0_wmux_0_Y[4]\, 
        \APB3_RDATA_1_25_0_0_y0[4]\, \APB3_RDATA_1_25_0_0_co0[4]\, 
        \APB3_RDATA_1_25_0_wmux_0_Y[3]\, 
        \APB3_RDATA_1_25_0_0_y0[3]\, \APB3_RDATA_1_25_0_0_co0[3]\, 
        \APB3_RDATA_1_14_0_wmux_0_Y[4]\, 
        \APB3_RDATA_1_14_0_0_y0[4]\, \APB3_RDATA_1_14_0_0_co0[4]\, 
        \APB3_RDATA_1_14_0_wmux_0_Y[3]\, 
        \APB3_RDATA_1_14_0_0_y0[3]\, \APB3_RDATA_1_14_0_0_co0[3]\, 
        \APB3_RDATA_1_14_0_wmux_0_Y[2]\, 
        \APB3_RDATA_1_14_0_0_y0[2]\, \APB3_RDATA_1_14_0_0_co0[2]\, 
        \APB3_RDATA_1_25_0_wmux_0_Y[2]\, 
        \APB3_RDATA_1_25_0_0_y0[2]\, \APB3_RDATA_1_25_0_0_co0[2]\, 
        \APB3_RDATA_1_0_m2_2_wmux_0_Y[0]\, 
        \APB3_RDATA_1_0_m2_2_2_y0[0]\, 
        \APB3_RDATA_1_0_m2_2_2_co0[0]\, 
        \APB3_RDATA_1_25_0_wmux_0_Y[6]\, 
        \APB3_RDATA_1_25_0_0_y0[6]\, \APB3_RDATA_1_25_0_0_co0[6]\, 
        \APB3_RDATA_1_25_0_wmux_0_Y[1]\, 
        \APB3_RDATA_1_25_0_0_y0[1]\, \APB3_RDATA_1_25_0_0_co0[1]\, 
        N_1641, \APB3_RDATA_1_21_0_0_y0[4]\, 
        \APB3_RDATA_1_21_0_0_co0[4]\, N_1643, 
        \APB3_RDATA_1_21_0_0_y0[6]\, \APB3_RDATA_1_21_0_0_co0[6]\, 
        N_1642, \APB3_RDATA_1_21_0_0_y0[5]\, 
        \APB3_RDATA_1_21_0_0_co0[5]\, N_1624, 
        \APB3_RDATA_1_19_0_0_y0[3]\, \APB3_RDATA_1_19_0_0_co0[3]\, 
        N_1627, \APB3_RDATA_1_19_0_0_y0[6]\, 
        \APB3_RDATA_1_19_0_0_co0[6]\, N_1623, 
        \APB3_RDATA_1_19_0_0_y0[2]\, \APB3_RDATA_1_19_0_0_co0[2]\, 
        N_204, \APB3_RDATA_1_18_i_m2_0_0_y0[7]\, 
        \APB3_RDATA_1_18_i_m2_0_0_co0[7]\, N_1626, 
        \APB3_RDATA_1_19_0_0_y0[5]\, \APB3_RDATA_1_19_0_0_co0[5]\, 
        N_1609, \APB3_RDATA_1_17_0_0_y0[4]\, 
        \APB3_RDATA_1_17_0_0_co0[4]\, N_1610, 
        \APB3_RDATA_1_17_0_0_y0[5]\, \APB3_RDATA_1_17_0_0_co0[5]\, 
        N_1640, \APB3_RDATA_1_21_0_0_y0[3]\, 
        \APB3_RDATA_1_21_0_0_co0[3]\, N_496, 
        \APB3_RDATA_1_24_i_m3_0_2_y0[1]\, 
        \APB3_RDATA_1_24_i_m3_0_2_co0[1]\, N_206, 
        \APB3_RDATA_1_18_i_m2_0_0_y0[5]\, 
        \APB3_RDATA_1_18_i_m2_0_0_co0[5]\, N_497, 
        \APB3_RDATA_1_24_i_m3_1_2_y0[1]\, 
        \APB3_RDATA_1_24_i_m3_1_2_co0[1]\, N_197, 
        \APB3_RDATA_1_18_i_m2_0_0_y0[0]\, 
        \APB3_RDATA_1_18_i_m2_0_0_co0[0]\, N_1611, 
        \APB3_RDATA_1_17_0_0_y0[6]\, \APB3_RDATA_1_17_0_0_co0[6]\, 
        N_1625, \APB3_RDATA_1_19_0_0_y0[4]\, 
        \APB3_RDATA_1_19_0_0_co0[4]\, N_201, 
        \APB3_RDATA_1_18_i_m2_0_0_y0[4]\, 
        \APB3_RDATA_1_18_i_m2_0_0_co0[4]\, N_593, 
        \APB3_RDATA_1_0_m2_8_2_y0[0]\, 
        \APB3_RDATA_1_0_m2_8_2_co0[0]\, N_495, 
        \APB3_RDATA_1_26_i_m3_0_2_y0[1]\, 
        \APB3_RDATA_1_26_i_m3_0_2_co0[1]\, N_1341, 
        \APB3_RDATA_1_17_i_m2_0_0_y0[3]\, 
        \APB3_RDATA_1_17_i_m2_0_0_co0[3]\, N_202, 
        \APB3_RDATA_1_21_i_m2_0_0_y0[2]\, 
        \APB3_RDATA_1_21_i_m2_0_0_co0[2]\, N_698, 
        \APB3_RDATA_1_17_i_m2_0_0_y0[0]\, 
        \APB3_RDATA_1_17_i_m2_0_0_co0[0]\, N_199, 
        \APB3_RDATA_1_18_i_m2_0_0_y0[2]\, 
        \APB3_RDATA_1_18_i_m2_0_0_co0[2]\, N_1628, 
        \APB3_RDATA_1_19_0_0_y0[7]\, \APB3_RDATA_1_19_0_0_co0[7]\, 
        N_205, \APB3_RDATA_1_18_i_m2_0_0_y0[6]\, 
        \APB3_RDATA_1_18_i_m2_0_0_co0[6]\, N_1342, 
        \APB3_RDATA_1_17_i_m2_0_0_y0[2]\, 
        \APB3_RDATA_1_17_i_m2_0_0_co0[2]\, N_200, 
        \APB3_RDATA_1_18_i_m2_0_0_y0[3]\, 
        \APB3_RDATA_1_18_i_m2_0_0_co0[3]\, N_697, 
        \APB3_RDATA_1_19_i_m2_0_0_y0[0]\, 
        \APB3_RDATA_1_19_i_m2_0_0_co0[0]\, N_1644, 
        \APB3_RDATA_1_21_0_0_y0[7]\, \APB3_RDATA_1_21_0_0_co0[7]\, 
        N_198, \APB3_RDATA_1_18_i_m2_0_0_y0[1]\, 
        \APB3_RDATA_1_18_i_m2_0_0_co0[1]\, N_1612, 
        \APB3_RDATA_1_17_0_0_y0[7]\, \APB3_RDATA_1_17_0_0_co0[7]\, 
        N_110, \APB3_RDATA_1_14_4_0_y1[1]\, 
        \APB3_RDATA_1_14_4_0_y3[1]\, \APB3_RDATA_1_14_4_co1_0[1]\, 
        \APB3_RDATA_1_14_4_y0_0[1]\, \APB3_RDATA_1_14_4_co0_0[1]\, 
        \APB3_RDATA_1_14_4_0_co1[1]\, \APB3_RDATA_1_14_4_0_y0[1]\, 
        \APB3_RDATA_1_14_4_0_co0[1]\, N_91, N_78, 
        \APB3_RDATA_1_am[1]_net_1\, \APB3_RDATA_1_bm[1]_net_1\, 
        \APB3_RDATA_1_am[2]_net_1\, \APB3_RDATA_1_bm[2]_net_1\, 
        N_1692, \APB3_RDATA_1_d_ns[5]_net_1\, N_1693, 
        \APB3_RDATA_1_d_ns[6]_net_1\, 
        \APB3_RDATA_1_0_m2_2_3[0]_net_1\, N_252, \N_817_i\, N_783, 
        N_1087, N_1496, \APB3_RDATA_1_25_3[7]_net_1\, N_51, 
        N_1494, \APB3_RDATA_1_25_3[5]_net_1\, N_50, N_1493, 
        \APB3_RDATA_1_25_3[4]_net_1\, N_49, N_1492, 
        \APB3_RDATA_1_25_3[3]_net_1\, N_48, N_1491, 
        \APB3_RDATA_1_25_3[2]_net_1\, N_52, N_1495, 
        \APB3_RDATA_1_25_3[6]_net_1\, N_137, N_1086, 
        \APB3_RDATA_1_25_3[1]_net_1\, N_3, N_577, N_1658, 
        \APB3_RDATA_1_am_1[4]_net_1\, \APB3_RDATA_1_am[4]_net_1\, 
        N_1666, N_757, N_1674, N_1655, N_1350, 
        \APB3_RDATA_1_bm_1[1]_net_1\, APB3_RDATA_1_sn_m12_i_0_0, 
        N_490, N_1656, \APB3_RDATA_1_bm_1[2]_net_1\, N_1501, 
        N_1583, APB3_RDATA_1_sn_m21_i_1, 
        \APB3_RDATA_1_0_m2_1_0[0]_net_1\, N_741, 
        \APB3_RDATA_1_29_d_bm_1_0[7]_net_1\, 
        \APB3_RDATA_1_29_d_bm[7]_net_1\, \APB3_RDATA_1_27_10\, 
        \APB3_RDATA_1_27_1[6]_net_1\, APB3_RDATA_1_sn_m12_i_0, 
        N_1595, N_1651, \APB3_RDATA_1_27_1[5]_net_1\, N_1594, 
        N_1650, \APB3_RDATA_1_23_1[7]_net_1\, \APB3_RDATA_1_23_1\, 
        \APB3_RDATA_1_23_2\, N_1661, N_385, 
        \APB3_RDATA_1_23_1[3]_net_1\, N_1657, N_381, 
        \APB3_RDATA_1_22_1_0[6]_net_1\, 
        \APB3_RDATA_1_22_1_0[5]_net_1\, 
        \APB3_RDATA_1_0_m2_6_2[0]_net_1\, N_586, 
        \APB3_RDATA_1_bm[4]_net_1\, \APB3_RDATA_1_s[3]_net_1\, 
        \APB3_RDATA_1_29_d_am[7]_net_1\, 
        \APB3_RDATA_1_29_d_ns[7]_net_1\, 
        \APB3_RDATA_1_d_bm[6]_net_1\, 
        \APB3_RDATA_1_d_am[6]_net_1\, 
        \APB3_RDATA_1_29_d_bm[3]_net_1\, 
        \APB3_RDATA_1_29_d_am[3]_net_1\, 
        \APB3_RDATA_1_29_d_ns[3]_net_1\, 
        \APB3_RDATA_1_d_bm[5]_net_1\, 
        \APB3_RDATA_1_d_am[5]_net_1\, 
        \APB3_RDATA_1_0_m2_3_am[0]_net_1\, 
        \APB3_RDATA_1_0_m2_3_bm[0]_net_1\, N_615, N_1700, 
        \APB3_RDATA_1_d_ns[3]_net_1\, N_1704, 
        \APB3_RDATA_1_d_ns[7]_net_1\, N_1677, N_1675, N_1673, 
        \APB3_RDATA_1_14_3[4]_net_1\, N_1585, 
        \APB3_RDATA_1_14_2[4]_net_1\, 
        \APB3_RDATA_1_14_3[3]_net_1\, N_1584, 
        \APB3_RDATA_1_14_2[3]_net_1\, 
        \APB3_RDATA_1_14_3[2]_net_1\, 
        \APB3_RDATA_1_14_2[2]_net_1\, N_1672, N_597, N_1676, 
        N_1671, N_790, N_801, N_732, 
        un13_mac_4_byte_5_reg_en_0_a2_0_a2_0_a2_0, 
        un13_mac_4_byte_1_reg_en_0_a2_0_a2_0_o2_0, N_802, N_796, 
        N_795, N_791, N_1357, N_1503, N_1502, N_1669, N_1682, 
        N_1667, N_1665, N_1664, N_203, N_582, N_1668, N_498, 
        N_499, un13_mac_4_byte_4_reg_en_0_a2_0_a2_0_a2_1, 
        un13_mac_4_byte_3_reg_en_0_a2_4_a2_5_a2_2, \m14_0_a3_1\, 
        un1_RX_packet_depthlto7_5, un1_RX_packet_depthlto7_4, 
        N_353_1, N_1455, N_785, N_1457, N_547, N_576, 
        tx_FIFO_UNDERRUN_int, tx_FIFO_OVERFLOW_int, N_1593, 
        rx_FIFO_OVERFLOW_int, N_186, N_384, rx_CRC_error_int, 
        N_185, APB3_RDATA_1_sn_m26_i_1, N_1649, N_1699, N_789, 
        N_234, N_1461, N_793, N_1698, N_799, N_549, N_742_0, 
        N_729, m30_0_0, N_989, \APB3_RDATA_1_0_a2_1[0]\, N_556, 
        N_8, N_10, N_570, N_561, N_726, N_581, N_1337, N_731
         : std_logic;

    for all : Interrupts
	Use entity work.Interrupts(DEF_ARCH);
begin 

    consumer_type4_reg(9) <= \consumer_type4_reg[9]\;
    consumer_type4_reg(8) <= \consumer_type4_reg[8]\;
    consumer_type4_reg(7) <= \consumer_type4_reg[7]\;
    consumer_type4_reg(6) <= \consumer_type4_reg[6]\;
    consumer_type4_reg(5) <= \consumer_type4_reg[5]\;
    consumer_type4_reg(4) <= \consumer_type4_reg[4]\;
    consumer_type4_reg(3) <= \consumer_type4_reg[3]\;
    consumer_type4_reg(2) <= \consumer_type4_reg[2]\;
    consumer_type4_reg(1) <= \consumer_type4_reg[1]\;
    consumer_type4_reg(0) <= \consumer_type4_reg[0]\;
    consumer_type3_reg(9) <= \consumer_type3_reg[9]\;
    consumer_type3_reg(8) <= \consumer_type3_reg[8]\;
    consumer_type3_reg(7) <= \consumer_type3_reg[7]\;
    consumer_type3_reg(6) <= \consumer_type3_reg[6]\;
    consumer_type3_reg(5) <= \consumer_type3_reg[5]\;
    consumer_type3_reg(4) <= \consumer_type3_reg[4]\;
    consumer_type3_reg(3) <= \consumer_type3_reg[3]\;
    consumer_type3_reg(2) <= \consumer_type3_reg[2]\;
    consumer_type3_reg(1) <= \consumer_type3_reg[1]\;
    consumer_type3_reg(0) <= \consumer_type3_reg[0]\;
    consumer_type2_reg(9) <= \consumer_type2_reg[9]\;
    consumer_type2_reg(8) <= \consumer_type2_reg[8]\;
    consumer_type2_reg(7) <= \consumer_type2_reg[7]\;
    consumer_type2_reg(6) <= \consumer_type2_reg[6]\;
    consumer_type2_reg(5) <= \consumer_type2_reg[5]\;
    consumer_type2_reg(4) <= \consumer_type2_reg[4]\;
    consumer_type2_reg(3) <= \consumer_type2_reg[3]\;
    consumer_type2_reg(2) <= \consumer_type2_reg[2]\;
    consumer_type2_reg(1) <= \consumer_type2_reg[1]\;
    consumer_type2_reg(0) <= \consumer_type2_reg[0]\;
    consumer_type1_reg(9) <= \consumer_type1_reg[9]\;
    consumer_type1_reg(8) <= \consumer_type1_reg[8]\;
    consumer_type1_reg(7) <= \consumer_type1_reg[7]\;
    consumer_type1_reg(6) <= \consumer_type1_reg[6]\;
    consumer_type1_reg(5) <= \consumer_type1_reg[5]\;
    consumer_type1_reg(4) <= \consumer_type1_reg[4]\;
    consumer_type1_reg(3) <= \consumer_type1_reg[3]\;
    consumer_type1_reg(2) <= \consumer_type1_reg[2]\;
    consumer_type1_reg(1) <= \consumer_type1_reg[1]\;
    consumer_type1_reg(0) <= \consumer_type1_reg[0]\;
    up_EOP_sync(2) <= \up_EOP_sync[2]_net_1\;
    up_EOP_sync(1) <= \up_EOP_sync[1]_net_1\;
    TX_FIFO_RST <= \TX_FIFO_RST\;
    start_tx_FIFO <= \start_tx_FIFO\;
    internal_loopback <= \internal_loopback\;
    external_loopback <= \external_loopback\;

    \READ_FIFO_ENABLE_PROC.un109_apb3_addr_0_a2_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => N_790, D => N_793, Y
         => N_330);
    
    \APB3_RDATA_1_24_i_m3_1_2_wmux[1]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => \external_loopback\, 
        D => \mac_2_byte_3_reg[1]_net_1\, FCI => VCC_net_1, S => 
        OPEN, Y => \APB3_RDATA_1_24_i_m3_1_2_y0[1]\, FCO => 
        \APB3_RDATA_1_24_i_m3_1_2_co0[1]\);
    
    \mac_3_byte_1_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_1_reg[7]_net_1\);
    
    \mac_2_byte_4_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_4_reg[3]_net_1\);
    
    \APB3_RDATA_1_19_0_wmux_0[7]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_19_0_0_y0[7]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \mac_2_byte_5_reg[7]_net_1\, D => 
        \mac_4_byte_1_reg[7]_net_1\, FCI => 
        \APB3_RDATA_1_19_0_0_co0[7]\, S => OPEN, Y => N_1628, FCO
         => OPEN);
    
    \mac_2_byte_3_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_3_reg[4]_net_1\);
    
    \mac_2_byte_2_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type4_reg[3]\);
    
    \APB3_RDATA_1_25_3[3]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_49, B => CoreAPB3_0_APBmslave0_PADDR(3), C
         => N_1492, Y => \APB3_RDATA_1_25_3[3]_net_1\);
    
    \i_int_mask_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_1354_i, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \i_int_mask_reg[3]_net_1\);
    
    iRX_FIFO_rd_en : SLE
      port map(D => \iAPB3_READY_i[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_330, ALn => N_854_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => RX_FIFO_rd_en);
    
    \mac_3_byte_2_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_2_reg[0]_net_1\);
    
    \APB3_RDATA_1_14_4_wmux_3[1]\ : ARI1
      generic map(INIT => x"0EC2C")

      port map(A => \APB3_RDATA_1_14_4_0_y3[1]\, B => 
        \APB3_RDATA_1_14_4_0_y1[1]\, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), D => VCC_net_1, FCI => 
        \APB3_RDATA_1_14_4_co1_0[1]\, S => OPEN, Y => N_110, FCO
         => OPEN);
    
    \REG_WRITE_PROC.un13_mac_4_byte_3_reg_en_0_a2_4_a2_5_a2_2\ : 
        CFG4
      generic map(INIT => x"0100")

      port map(A => \int_mask_reg_en\, B => \mac_4_byte_2_reg_en\, 
        C => N_743, D => \mac_4_byte_3_reg_en\, Y => 
        un13_mac_4_byte_3_reg_en_0_a2_4_a2_5_a2_2);
    
    \WRITE_REGISTER_ENABLE_PROC.un97_apb3_addr_0_a2\ : CFG3
      generic map(INIT => x"80")

      port map(A => N_801, B => CoreAPB3_0_APBmslave0_PADDR(7), C
         => N_791, Y => N_356);
    
    \APB3_RDATA_1_bm[2]\ : CFG4
      generic map(INIT => x"8F88")

      port map(A => N_1656, B => N_1350, C => \N_817_i\, D => 
        \APB3_RDATA_1_bm_1[2]_net_1\, Y => 
        \APB3_RDATA_1_bm[2]_net_1\);
    
    \i_int_mask_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_1354_i, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \i_int_mask_reg[4]_net_1\);
    
    \APB3_RDATA_1_26_i_m3_0_2_wmux[1]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_2_byte_4_reg[1]_net_1\, D => 
        \mac_2_byte_6_reg[1]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_26_i_m3_0_2_y0[1]\, FCO => 
        \APB3_RDATA_1_26_i_m3_0_2_co0[1]\);
    
    \mac_2_byte_3_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_3_reg[3]_net_1\);
    
    \mac_2_byte_2_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type4_reg[4]\);
    
    \APB3_RDATA_1_29_d_am[3]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_1640, B => N_200, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => 
        \APB3_RDATA_1_29_d_am[3]_net_1\);
    
    \APB3_RDATA_1_14_0_0_wmux[3]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => ReadFIFO_Read_Ptr(0), B => 
        ReadFIFO_Read_Ptr(1), C => N_652, D => N_659, FCI => 
        VCC_net_1, S => OPEN, Y => \APB3_RDATA_1_14_0_0_y0[3]\, 
        FCO => \APB3_RDATA_1_14_0_0_co0[3]\);
    
    \RX_packet_depth_cry[1]\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \RX_packet_depth[1]_net_1\, B => 
        rx_packet_complt, C => GND_net_1, D => GND_net_1, FCI => 
        \RX_packet_depth_cry[0]_net_1\, S => 
        \RX_packet_depth_s[1]\, Y => OPEN, FCO => 
        \RX_packet_depth_cry[1]_net_1\);
    
    \APB3_RDATA_RNIDFI5[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        \CoreAPB3_0_APBmslave0_PRDATA[0]\, Y => 
        CoreAPB3_0_APBmslave0_PRDATA_m(0));
    
    \RX_packet_depth_cry[5]\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \RX_packet_depth[5]_net_1\, B => 
        rx_packet_complt, C => GND_net_1, D => GND_net_1, FCI => 
        \RX_packet_depth_cry[4]_net_1\, S => 
        \RX_packet_depth_s[5]\, Y => OPEN, FCO => 
        \RX_packet_depth_cry[5]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_4_byte_1_reg_en_0_a2_0_a2_0_o2_0_0\ : 
        CFG2
      generic map(INIT => x"E")

      port map(A => \mac_3_byte_3_reg_en\, B => 
        \mac_3_byte_4_reg_en\, Y => 
        un13_mac_4_byte_1_reg_en_0_a2_0_a2_0_o2_0);
    
    \APB3_RDATA_1_19_0_0_wmux[7]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \i_int_mask_reg[7]_net_1\, D => 
        \mac_1_byte_3_reg[7]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_19_0_0_y0[7]\, FCO => 
        \APB3_RDATA_1_19_0_0_co0[7]\);
    
    \mac_4_byte_5_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_5_reg[7]_net_1\);
    
    \mac_3_byte_3_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_3_reg[0]_net_1\);
    
    \APB3_RDATA_1_18_i_m2_0_wmux_0[0]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_18_i_m2_0_0_y0[0]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_5_reg[0]_net_1\, D => 
        \mac_4_byte_6_reg[0]_net_1\, FCI => 
        \APB3_RDATA_1_18_i_m2_0_0_co0[0]\, S => OPEN, Y => N_197, 
        FCO => OPEN);
    
    \up_EOP_sync[2]\ : SLE
      port map(D => \up_EOP_sync[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \up_EOP_sync[2]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.apb3_addr_0_a2\ : CFG3
      generic map(INIT => x"80")

      port map(A => N_790, B => N_793, C => N_791, Y => N_329);
    
    \APB3_RDATA_1_26[4]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_1641, B => N_201, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_1682);
    
    \APB3_RDATA_1_29_d_bm_RNO[3]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \APB3_RDATA_1_14_0_wmux_0_Y[3]\, B => 
        \APB3_RDATA_1_14_3[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_1584);
    
    \APB3_RDATA_1_am_1[4]\ : CFG3
      generic map(INIT => x"47")

      port map(A => N_1666, B => N_757, C => N_1674, Y => 
        \APB3_RDATA_1_am_1[4]_net_1\);
    
    \REG_WRITE_PROC.control_reg_3[5]\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(5), B => 
        \control_reg_en\, Y => \control_reg_3[5]\);
    
    \mac_4_byte_5_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_5_reg[4]_net_1\);
    
    control_reg_en_0 : CFG4
      generic map(INIT => x"7430")

      port map(A => CoreAPB3_0_APBmslave0_PREADY, B => N_331, C
         => \control_reg_en\, D => \iAPB3_READY[0]_net_1\, Y => 
        N_3);
    
    \APB3_RDATA_1_17_i_m2_0_0_wmux[0]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \control_reg[0]_net_1\, D => \mac_2_byte_3_reg[0]_net_1\, 
        FCI => VCC_net_1, S => OPEN, Y => 
        \APB3_RDATA_1_17_i_m2_0_0_y0[0]\, FCO => 
        \APB3_RDATA_1_17_i_m2_0_0_co0[0]\);
    
    \APB3_RDATA_1_18_i_m2_0_0_wmux[6]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_3_reg[6]_net_1\, D => 
        \mac_4_byte_4_reg[6]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_18_i_m2_0_0_y0[6]\, FCO => 
        \APB3_RDATA_1_18_i_m2_0_0_co0[6]\);
    
    \mac_2_byte_2_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type4_reg[2]\);
    
    \APB3_RDATA_1_19_0_0_wmux[4]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \i_int_mask_reg[4]_net_1\, D => 
        \mac_1_byte_3_reg[4]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_19_0_0_y0[4]\, FCO => 
        \APB3_RDATA_1_19_0_0_co0[4]\);
    
    \control_reg[5]\ : SLE
      port map(D => \control_reg_3[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un1_control_reg_en_2_i_0, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \start_tx_FIFO\);
    
    \mac_2_byte_3_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_3_reg[2]_net_1\);
    
    \mac_3_byte_5_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_5_reg[3]_net_1\);
    
    mac_1_byte_3_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_337, ALn => N_855_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_1_byte_3_reg_en\);
    
    \WRITE_REGISTER_ENABLE_PROC.un65_apb3_addr_0_a2_0_RNIU8TB1\ : 
        CFG4
      generic map(INIT => x"5073")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => N_791, D => N_757, Y
         => APB3_RDATA_1_sn_m26_i_1);
    
    \APB3_RDATA_1_bm_1_RNO[2]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \APB3_RDATA_1_14_0_wmux_0_Y[2]\, B => 
        \APB3_RDATA_1_14_3[2]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_1583);
    
    \APB3_RDATA_1_25_0_wmux_0[3]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_25_0_0_y0[3]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_1_reg[3]_net_1\, D => 
        \mac_3_byte_3_reg[3]_net_1\, FCI => 
        \APB3_RDATA_1_25_0_0_co0[3]\, S => OPEN, Y => 
        \APB3_RDATA_1_25_0_wmux_0_Y[3]\, FCO => OPEN);
    
    \mac_4_byte_6_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_6_reg[6]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_3_byte_1_reg_en_0_a2_1_a2_0_o2\ : 
        CFG3
      generic map(INIT => x"FE")

      port map(A => \mac_2_byte_6_reg_en\, B => 
        \mac_2_byte_5_reg_en\, C => N_547, Y => N_549);
    
    read_reg_en_RNIG54T2 : CFG4
      generic map(INIT => x"FBFF")

      port map(A => N_252, B => \read_reg_en\, C => \N_817_i\, D
         => N_783, Y => N_78);
    
    mac_4_byte_6_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_358, ALn => N_855_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_4_byte_6_reg_en\);
    
    \APB3_RDATA_RNIFHI5[2]\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        \CoreAPB3_0_APBmslave0_PRDATA[2]\, Y => 
        CoreAPB3_0_APBmslave0_PRDATA_m(2));
    
    \APB3_RDATA_1_18_i_m2_0_wmux_0[1]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_18_i_m2_0_0_y0[1]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_5_reg[1]_net_1\, D => 
        \mac_4_byte_6_reg[1]_net_1\, FCI => 
        \APB3_RDATA_1_18_i_m2_0_0_co0[1]\, S => OPEN, Y => N_198, 
        FCO => OPEN);
    
    \mac_3_byte_5_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_5_reg[6]_net_1\);
    
    \mac_1_byte_5_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type3_reg[8]\);
    
    mac_1_byte_2_reg_en_0 : CFG4
      generic map(INIT => x"CAAA")

      port map(A => \mac_1_byte_2_reg_en\, B => 
        mac_4_byte_6_reg_en_1, C => N_802, D => N_799, Y => N_6);
    
    \mac_2_byte_5_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_5_reg[2]_net_1\);
    
    \APB3_RDATA_1_3[6]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \consumer_type4_reg[6]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_4_reg[6]_net_1\, Y => N_1495);
    
    mac_1_byte_2_reg_en_ret_1 : SLE
      port map(D => N_6, CLK => m2s010_som_sb_0_CCC_71MHz, EN => 
        VCC_net_1, ALn => N_855_i_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        N_6_reto);
    
    \APB3_RDATA_1_am[4]\ : CFG3
      generic map(INIT => x"8B")

      port map(A => N_1658, B => N_91, C => 
        \APB3_RDATA_1_am_1[4]_net_1\, Y => 
        \APB3_RDATA_1_am[4]_net_1\);
    
    \mac_4_byte_4_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_4_reg[2]_net_1\);
    
    \APB3_RDATA_1_19_i_m2_0_wmux_0[0]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_19_i_m2_0_0_y0[0]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \mac_2_byte_5_reg[0]_net_1\, D => 
        \mac_4_byte_1_reg[0]_net_1\, FCI => 
        \APB3_RDATA_1_19_i_m2_0_0_co0[0]\, S => OPEN, Y => N_697, 
        FCO => OPEN);
    
    \APB3_RDATA_1_19_0_wmux_0[5]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_19_0_0_y0[5]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \mac_2_byte_5_reg[5]_net_1\, D => 
        \mac_4_byte_1_reg[5]_net_1\, FCI => 
        \APB3_RDATA_1_19_0_0_co0[5]\, S => OPEN, Y => N_1626, FCO
         => OPEN);
    
    \APB3_RDATA[5]\ : SLE
      port map(D => \APB3_RDATA_1[5]_net_1\, CLK => N_41_mux, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        \CoreAPB3_0_APBmslave0_PRDATA[5]\);
    
    \mac_4_byte_3_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_3_reg[5]_net_1\);
    
    \APB3_RDATA_1_14_2[3]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => ReadFIFO_Read_Ptr(1), B => TX_FIFO_Full, C
         => ReadFIFO_Read_Ptr(0), Y => 
        \APB3_RDATA_1_14_2[3]_net_1\);
    
    \APB3_RDATA_1_14_2[2]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => ReadFIFO_Read_Ptr(1), B => TX_FIFO_Empty, C
         => ReadFIFO_Read_Ptr(0), Y => 
        \APB3_RDATA_1_14_2[2]_net_1\);
    
    \APB3_RDATA_1_24[6]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_1611, B => CoreAPB3_0_APBmslave0_PADDR(3), 
        C => N_1627, Y => N_1668);
    
    \WRITE_REGISTER_ENABLE_PROC.un57_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_789, D => N_795, Y
         => N_346);
    
    \mac_4_byte_5_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_5_reg[5]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_4_byte_6_reg_en_0_a2_4_a2_3_o2\ : 
        CFG4
      generic map(INIT => x"FFFE")

      port map(A => \mac_4_byte_5_reg_en\, B => 
        \mac_4_byte_4_reg_en\, C => \mac_4_byte_3_reg_en\, D => 
        \mac_4_byte_2_reg_en\, Y => N_577);
    
    \APB3_RDATA_1_19_0_wmux_0[3]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_19_0_0_y0[3]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \mac_2_byte_5_reg[3]_net_1\, D => 
        \mac_4_byte_1_reg[3]_net_1\, FCI => 
        \APB3_RDATA_1_19_0_0_co0[3]\, S => OPEN, Y => N_1624, FCO
         => OPEN);
    
    \APB3_RDATA_1_17_i_m2_0_wmux_0[0]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_17_i_m2_0_0_y0[0]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \consumer_type1_reg[8]\, D => \mac_3_byte_5_reg[0]_net_1\, 
        FCI => \APB3_RDATA_1_17_i_m2_0_0_co0[0]\, S => OPEN, Y
         => N_698, FCO => OPEN);
    
    \APB3_RDATA_1_25_0_0_wmux[7]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_1_byte_5_reg[7]_net_1\, D => 
        \mac_2_byte_1_reg[7]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_25_0_0_y0[7]\, FCO => 
        \APB3_RDATA_1_25_0_0_co0[7]\);
    
    \APB3_RDATA_1_22_i_m3_0[1]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \consumer_type3_reg[1]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \scratch_pad_reg[1]_net_1\, Y => N_490);
    
    \APB3_RDATA_1_19_0_wmux_0[2]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_19_0_0_y0[2]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \mac_2_byte_5_reg[2]_net_1\, D => 
        \mac_4_byte_1_reg[2]_net_1\, FCI => 
        \APB3_RDATA_1_19_0_0_co0[2]\, S => OPEN, Y => N_1623, FCO
         => OPEN);
    
    \REG_WRITE_PROC.un13_mac_2_byte_1_reg_en_0_a2_2_a2_1_a2\ : 
        CFG4
      generic map(INIT => x"4000")

      port map(A => \mac_1_byte_6_reg_en\, B => 
        \mac_2_byte_1_reg_en\, C => N_1461, D => N_1457, Y => 
        un13_mac_2_byte_1_reg_en);
    
    \APB3_RDATA_1_19_0_wmux_0[4]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_19_0_0_y0[4]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \mac_2_byte_5_reg[4]_net_1\, D => 
        \mac_4_byte_1_reg[4]_net_1\, FCI => 
        \APB3_RDATA_1_19_0_0_co0[4]\, S => OPEN, Y => N_1625, FCO
         => OPEN);
    
    \scratch_pad_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \write_scratch_reg_en\, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \scratch_pad_reg[3]_net_1\);
    
    \APB3_RDATA_1_22[4]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => N_1503, 
        C => N_1585, Y => N_1649);
    
    \APB3_RDATA_1_bm[4]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N_1682, B => N_1649, C => N_78, Y => 
        \APB3_RDATA_1_bm[4]_net_1\);
    
    \mac_1_byte_5_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_5_reg[7]_net_1\);
    
    control_reg_en_ret_RNID0IJ : CFG2
      generic map(INIT => x"2")

      port map(A => \int_mask_reg_en\, B => N_743, Y => N_1354_i);
    
    \APB3_RDATA_1_19_0_wmux_0[6]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_19_0_0_y0[6]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \mac_2_byte_5_reg[6]_net_1\, D => 
        \mac_4_byte_1_reg[6]_net_1\, FCI => 
        \APB3_RDATA_1_19_0_0_co0[6]\, S => OPEN, Y => N_1627, FCO
         => OPEN);
    
    \WRITE_REGISTER_ENABLE_PROC.un53_apb3_addr_0_a2_0_a2_0\ : 
        CFG2
      generic map(INIT => x"4")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), Y => N_795);
    
    \mac_2_byte_1_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_1_reg[4]_net_1\);
    
    \mac_1_byte_5_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_5_reg[4]_net_1\);
    
    \APB3_RDATA_1_17_0_0_wmux[6]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => rx_FIFO_rst_reg, D
         => \mac_2_byte_3_reg[6]_net_1\, FCI => VCC_net_1, S => 
        OPEN, Y => \APB3_RDATA_1_17_0_0_y0[6]\, FCO => 
        \APB3_RDATA_1_17_0_0_co0[6]\);
    
    \mac_3_byte_2_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_2_reg[7]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_1_byte_6_reg_en_0_a2_1_a2_1_a2_0\ : 
        CFG3
      generic map(INIT => x"01")

      port map(A => \mac_1_byte_5_reg_en\, B => 
        \mac_1_byte_4_reg_en\, C => \mac_1_byte_3_reg_en\, Y => 
        N_1457);
    
    \WRITE_REGISTER_ENABLE_PROC.un105_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(7), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => N_801, Y => N_358);
    
    \REG_WRITE_PROC.un12_mac_2_byte_1_reg_en_16_1\ : CFG4
      generic map(INIT => x"FFCA")

      port map(A => \mac_2_byte_1_reg_en\, B => 
        mac_4_byte_6_reg_en_1, C => N_341, D => N_8, Y => 
        un12_mac_2_byte_1_reg_en_16_1);
    
    \APB3_RDATA_1_19_i_m2_0_0_wmux[0]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \i_int_mask_reg[0]_net_1\, D => \consumer_type2_reg[8]\, 
        FCI => VCC_net_1, S => OPEN, Y => 
        \APB3_RDATA_1_19_i_m2_0_0_y0[0]\, FCO => 
        \APB3_RDATA_1_19_i_m2_0_0_co0[0]\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \APB3_RDATA_1_18_i_m2_0_0_wmux[7]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_3_reg[7]_net_1\, D => 
        \mac_4_byte_4_reg[7]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_18_i_m2_0_0_y0[7]\, FCO => 
        \APB3_RDATA_1_18_i_m2_0_0_co0[7]\);
    
    \APB3_RDATA_1_18_i_m2_0_wmux_0[4]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_18_i_m2_0_0_y0[4]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_5_reg[4]_net_1\, D => 
        \mac_4_byte_6_reg[4]_net_1\, FCI => 
        \APB3_RDATA_1_18_i_m2_0_0_co0[4]\, S => OPEN, Y => N_201, 
        FCO => OPEN);
    
    \mac_4_byte_1_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_1_reg[1]_net_1\);
    
    mac_1_byte_6_reg_en_0 : CFG3
      generic map(INIT => x"CA")

      port map(A => \mac_1_byte_6_reg_en\, B => 
        mac_4_byte_6_reg_en_1, C => N_340, Y => N_10);
    
    control_reg_en_ret_0 : SLE
      port map(D => N_733, CLK => m2s010_som_sb_0_CCC_71MHz, EN
         => VCC_net_1, ALn => N_855_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        N_742);
    
    \WRITE_REGISTER_ENABLE_PROC.apb3_addr_0_a2_1_0_a2\ : CFG4
      generic map(INIT => x"0001")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => 
        CoreAPB3_0_APBmslave0_PADDR(7), C => 
        CoreAPB3_0_APBmslave0_PADDR(0), D => 
        CoreAPB3_0_APBmslave0_PADDR(1), Y => N_793);
    
    \APB3_RDATA[7]\ : SLE
      port map(D => \APB3_RDATA_1[7]\, CLK => N_41_mux, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        \CoreAPB3_0_APBmslave0_PRDATA[7]\);
    
    \mac_4_byte_5_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_5_reg[1]_net_1\);
    
    \APB3_RDATA_1_25_0_wmux_0[7]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_25_0_0_y0[7]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_1_reg[7]_net_1\, D => 
        \mac_3_byte_3_reg[7]_net_1\, FCI => 
        \APB3_RDATA_1_25_0_0_co0[7]\, S => OPEN, Y => 
        \APB3_RDATA_1_25_0_wmux_0_Y[7]\, FCO => OPEN);
    
    \mac_2_byte_6_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_6_reg[1]_net_1\);
    
    \mac_2_byte_1_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type4_reg[8]\);
    
    \APB3_RDATA_1_14_2[4]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => ReadFIFO_Read_Ptr(1), B => 
        \RX_packet_depth_status\, C => ReadFIFO_Read_Ptr(0), Y
         => \APB3_RDATA_1_14_2[4]_net_1\);
    
    \mac_3_byte_3_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_3_reg[7]_net_1\);
    
    \mac_1_byte_6_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type3_reg[6]\);
    
    \APB3_RDATA_1_25_0_0_wmux[5]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_1_byte_5_reg[5]_net_1\, D => 
        \mac_2_byte_1_reg[5]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_25_0_0_y0[5]\, FCO => 
        \APB3_RDATA_1_25_0_0_co0[5]\);
    
    \mac_2_byte_6_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_6_reg[7]_net_1\);
    
    \mac_3_byte_3_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_3_reg[1]_net_1\);
    
    \REG_WRITE_PROC.un12_mac_1_byte_2_reg_en_20\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_732, B => N_6_reto, Y => N_731);
    
    \REG_WRITE_PROC.un13_mac_4_byte_3_reg_en_0_a2_4_a2_5_a2\ : 
        CFG4
      generic map(INIT => x"1000")

      port map(A => \mac_1_byte_2_reg_en\, B => 
        \mac_1_byte_1_reg_en\, C => 
        un13_mac_4_byte_3_reg_en_0_a2_4_a2_5_a2_2, D => N_1337, Y
         => un13_mac_4_byte_3_reg_en);
    
    mac_3_byte_6_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_352, ALn => N_855_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_3_byte_6_reg_en\);
    
    \APB3_RDATA_1_d_bm[6]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_1643, B => N_205, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => 
        \APB3_RDATA_1_d_bm[6]_net_1\);
    
    \APB3_RDATA_1_15[6]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \mac_4_byte_2_reg[6]_net_1\, B => N_384, C
         => CoreAPB3_0_APBmslave0_PADDR(3), Y => N_1595);
    
    \mac_1_byte_4_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type2_reg[2]\);
    
    \mac_2_byte_2_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type4_reg[5]\);
    
    \mac_4_byte_4_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_4_reg[7]_net_1\);
    
    \mac_1_byte_3_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_3_reg[5]_net_1\);
    
    \mac_4_byte_4_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_4_reg[6]_net_1\);
    
    \mac_4_byte_3_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_3_reg[6]_net_1\);
    
    \APB3_RDATA_1_23_1[7]\ : CFG4
      generic map(INIT => x"0C0A")

      port map(A => N_385, B => \mac_4_byte_2_reg[7]_net_1\, C
         => APB3_RDATA_1_sn_m12_i_0, D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => 
        \APB3_RDATA_1_23_1[7]_net_1\);
    
    \mac_2_byte_1_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_1_reg[6]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_1_byte_4_reg_en_0_a2_0_a2_0_a2\ : 
        CFG3
      generic map(INIT => x"20")

      port map(A => \mac_1_byte_4_reg_en\, B => 
        \mac_1_byte_3_reg_en\, C => N_1461, Y => 
        un13_mac_1_byte_4_reg_en);
    
    \REG_WRITE_PROC.un12_mac_2_byte_1_reg_en_16_2\ : CFG4
      generic map(INIT => x"FFCA")

      port map(A => \mac_1_byte_3_reg_en\, B => 
        mac_4_byte_6_reg_en_1, C => N_337, D => N_6, Y => 
        un12_mac_2_byte_1_reg_en_16_2);
    
    \i_int_mask_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_1354_i, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \i_int_mask_reg[7]_net_1\);
    
    \APB3_RDATA_1_3[3]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \consumer_type4_reg[3]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_4_reg[3]_net_1\, Y => N_1492);
    
    \mac_1_byte_5_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_5_reg[5]_net_1\);
    
    \RX_packet_depth_cry[0]\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \RX_packet_depth[0]_net_1\, B => 
        rx_packet_complt, C => GND_net_1, D => GND_net_1, FCI => 
        RX_packet_depth_s_390_FCO, S => \RX_packet_depth_s[0]\, Y
         => OPEN, FCO => \RX_packet_depth_cry[0]_net_1\);
    
    APB3_RDATA_1_sn_m26_i_a2_0 : CFG3
      generic map(INIT => x"80")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => N_785);
    
    \lfsr_c_i_i[4]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rx_crc_data_calc(11), B => 
        rx_crc_data_calc(10), C => RX_FIFO_DIN(3), D => 
        RX_FIFO_DIN(2), Y => lfsr_c_i_i_0);
    
    \mac_4_byte_4_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_4_reg[3]_net_1\);
    
    \APB3_RDATA_1_23[7]\ : CFG4
      generic map(INIT => x"FFF4")

      port map(A => \N_817_i\, B => \APB3_RDATA_1_23_1[7]_net_1\, 
        C => \APB3_RDATA_1_23_1\, D => \APB3_RDATA_1_23_2\, Y => 
        N_1661);
    
    \mac_4_byte_3_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_3_reg[4]_net_1\);
    
    \mac_4_byte_2_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_2_reg[3]_net_1\);
    
    \APB3_RDATA_1_19_0_0_wmux[6]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \i_int_mask_reg[6]_net_1\, D => 
        \mac_1_byte_3_reg[6]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_19_0_0_y0[6]\, FCO => 
        \APB3_RDATA_1_19_0_0_co0[6]\);
    
    \APB3_RDATA_1_0_m2_3_am[0]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \mac_3_byte_6_reg[0]_net_1\, B => 
        \mac_3_byte_2_reg[0]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => 
        \APB3_RDATA_1_0_m2_3_am[0]_net_1\);
    
    RX_packet_depth_s_390 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => rx_packet_complt, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => RX_packet_depth_s_390_FCO);
    
    \mac_2_byte_6_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_6_reg[4]_net_1\);
    
    
        \WRITE_REGISTER_ENABLE_PROC.un9_apb3_addr_0_a2_0_a2_0_a2_RNIDDPT_0\ : 
        CFG4
      generic map(INIT => x"0100")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => 
        CoreAPB3_0_APBmslave0_PADDR(0), C => 
        CoreAPB3_0_APBmslave0_PADDR(1), D => N_790, Y => N_801);
    
    \APB3_RDATA_1_14_4_wmux_0[1]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_14_4_0_y0[1]\, B => 
        ReadFIFO_Read_Ptr(1), C => RX_FIFO_DOUT_2_0, D => 
        RX_FIFO_DOUT_3_0, FCI => \APB3_RDATA_1_14_4_0_co0[1]\, S
         => OPEN, Y => \APB3_RDATA_1_14_4_0_y1[1]\, FCO => 
        \APB3_RDATA_1_14_4_0_co1[1]\);
    
    \APB3_RDATA_1_28[2]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => N_1664, B => N_757, C => N_1672, Y => N_1699);
    
    \SYNC2_APB3_CLK_PROC.RX_FIFO_RST_1\ : CFG2
      generic map(INIT => x"E")

      port map(A => RX_EarlyTerm, B => rx_FIFO_rst_reg, Y => 
        RX_FIFO_RST_1);
    
    \APB3_RDATA_1_s[3]\ : CFG3
      generic map(INIT => x"2A")

      port map(A => N_91, B => N_1350, C => N_78, Y => 
        \APB3_RDATA_1_s[3]_net_1\);
    
    mac_2_byte_4_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_344, ALn => N_855_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_2_byte_4_reg_en\);
    
    \mac_4_byte_3_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_3_reg[3]_net_1\);
    
    \mac_4_byte_2_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_2_reg[4]_net_1\);
    
    \APB3_RDATA_1_14_3[2]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => ReadFIFO_Read_Ptr(1), B => 
        \APB3_RDATA_1_14_2[2]_net_1\, C => TX_FIFO_Empty, Y => 
        \APB3_RDATA_1_14_3[2]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_4_byte_5_reg_en_0_a2_0_a2_0_a2_0\ : 
        CFG2
      generic map(INIT => x"4")

      port map(A => N_732, B => \mac_4_byte_5_reg_en\, Y => 
        un13_mac_4_byte_5_reg_en_0_a2_0_a2_0_a2_0);
    
    \APB3_RDATA_1_18_i_m2_0_wmux_0[6]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_18_i_m2_0_0_y0[6]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_5_reg[6]_net_1\, D => 
        \mac_4_byte_6_reg[6]_net_1\, FCI => 
        \APB3_RDATA_1_18_i_m2_0_0_co0[6]\, S => OPEN, Y => N_205, 
        FCO => OPEN);
    
    \mac_1_byte_1_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type1_reg[9]\);
    
    \REG_WRITE_PROC.un13_mac_4_byte_1_reg_en_0_a2_0_a2_0_o2_0\ : 
        CFG2
      generic map(INIT => x"E")

      port map(A => \mac_3_byte_5_reg_en\, B => 
        \mac_3_byte_6_reg_en\, Y => N_1357);
    
    N_854_i : CFG4
      generic map(INIT => x"0040")

      port map(A => CoreAPB3_0_APBmslave0_PWRITE, B => 
        CoreAPB3_0_APBmslave0_PSELx, C => 
        CoreAPB3_0_APBmslave0_PENABLE, D => long_reset, Y => 
        N_854_i_i);
    
    \mac_1_byte_5_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type3_reg[9]\);
    
    \REG_WRITE_PROC.un13_mac_4_byte_1_reg_en_0_a2_0_a2_0_o2\ : 
        CFG4
      generic map(INIT => x"FFFE")

      port map(A => \mac_3_byte_2_reg_en\, B => 
        \mac_3_byte_1_reg_en\, C => 
        un13_mac_4_byte_1_reg_en_0_a2_0_a2_0_o2_0, D => N_549, Y
         => N_561);
    
    \APB3_RDATA_1_21_0_0_wmux[7]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_2_byte_4_reg[7]_net_1\, D => 
        \mac_2_byte_6_reg[7]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_21_0_0_y0[7]\, FCO => 
        \APB3_RDATA_1_21_0_0_co0[7]\);
    
    \WRITE_REGISTER_ENABLE_PROC.un49_apb3_addr_0_a2_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_789, B => N_791, Y => N_799);
    
    \APB3_RDATA_1_d_bm[5]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_1642, B => N_206, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => 
        \APB3_RDATA_1_d_bm[5]_net_1\);
    
    \APB3_RDATA_1_17_i_m2_0_wmux_0[3]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_17_i_m2_0_0_y0[3]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_1_byte_1_reg[3]_net_1\, D => 
        \mac_3_byte_5_reg[3]_net_1\, FCI => 
        \APB3_RDATA_1_17_i_m2_0_0_co0[3]\, S => OPEN, Y => N_1341, 
        FCO => OPEN);
    
    \mac_2_byte_6_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_6_reg[2]_net_1\);
    
    \APB3_RDATA_1_25_0_wmux_0[5]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_25_0_0_y0[5]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_1_reg[5]_net_1\, D => 
        \mac_3_byte_3_reg[5]_net_1\, FCI => 
        \APB3_RDATA_1_25_0_0_co0[5]\, S => OPEN, Y => 
        \APB3_RDATA_1_25_0_wmux_0_Y[5]\, FCO => OPEN);
    
    \scratch_pad_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \write_scratch_reg_en\, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \scratch_pad_reg[5]_net_1\);
    
    \APB3_RDATA_1_28_RNO[7]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \APB3_RDATA_1_25_0_wmux_0_Y[7]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \APB3_RDATA_1_25_3[7]_net_1\, Y => N_1677);
    
    \mac_4_byte_2_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_2_reg[2]_net_1\);
    
    \mac_3_byte_5_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_5_reg[0]_net_1\);
    
    \mac_4_byte_3_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_3_reg[2]_net_1\);
    
    \APB3_RDATA_1_d_ns[7]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_1661, B => N_1704, C => N_91, Y => 
        \APB3_RDATA_1_d_ns[7]_net_1\);
    
    \APB3_RDATA_1_21_0_wmux_0[3]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_21_0_0_y0[3]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \consumer_type1_reg[3]\, D => \consumer_type2_reg[3]\, 
        FCI => \APB3_RDATA_1_21_0_0_co0[3]\, S => OPEN, Y => 
        N_1640, FCO => OPEN);
    
    \PROCESSOR_EOP_READ_PROC.un117_apb3_addr_0_a2_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \read_reg_en\, B => 
        CoreAPB3_0_APBmslave0_PREADY, C => N_712, D => N_330, Y
         => un117_apb3_addr);
    
    \mac_1_byte_4_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type2_reg[7]\);
    
    \mac_1_byte_4_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type2_reg[6]\);
    
    \mac_2_byte_2_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type4_reg[6]\);
    
    \mac_1_byte_3_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_3_reg[6]_net_1\);
    
    \mac_2_byte_2_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type4_reg[1]\);
    
    mac_1_byte_6_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_340, ALn => N_855_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_1_byte_6_reg_en\);
    
    \APB3_RDATA_1_ns[4]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \APB3_RDATA_1_bm[4]_net_1\, B => 
        \APB3_RDATA_1_s[3]_net_1\, C => 
        \APB3_RDATA_1_am[4]_net_1\, Y => \APB3_RDATA_1[4]\);
    
    \WRITE_REGISTER_ENABLE_PROC.un9_apb3_addr_0_a2_0_a2\ : CFG4
      generic map(INIT => x"2000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_789, D => N_790, Y
         => N_333);
    
    \RX_PACKET_DEPTH_STATUS_PROC.un1_RX_packet_depthlto7_4\ : 
        CFG4
      generic map(INIT => x"0001")

      port map(A => \RX_packet_depth[7]_net_1\, B => 
        \RX_packet_depth[6]_net_1\, C => 
        \RX_packet_depth[5]_net_1\, D => 
        \RX_packet_depth[4]_net_1\, Y => 
        un1_RX_packet_depthlto7_4);
    
    \mac_4_byte_5_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_5_reg[2]_net_1\);
    
    \mac_2_byte_1_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_1_reg[3]_net_1\);
    
    mac_1_byte_4_reg_en_0 : CFG3
      generic map(INIT => x"CA")

      port map(A => \mac_1_byte_4_reg_en\, B => 
        mac_4_byte_6_reg_en_1, C => N_338, Y => N_8);
    
    \APB3_RDATA_1_21_0_0_wmux[5]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_2_byte_4_reg[5]_net_1\, D => 
        \mac_2_byte_6_reg[5]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_21_0_0_y0[5]\, FCO => 
        \APB3_RDATA_1_21_0_0_co0[5]\);
    
    \APB3_RDATA_RNIJLI5[6]\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        \CoreAPB3_0_APBmslave0_PRDATA[6]\, Y => 
        CoreAPB3_0_APBmslave0_PRDATA_m(6));
    
    \APB3_RDATA_1_25_3[5]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_51, B => CoreAPB3_0_APBmslave0_PADDR(3), C
         => N_1494, Y => \APB3_RDATA_1_25_3[5]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un41_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_793, D => N_795, Y
         => N_342);
    
    \mac_1_byte_4_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type2_reg[3]\);
    
    \APB3_RDATA_1_24[3]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_1624, B => N_1341, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => N_1665);
    
    \APB3_RDATA_1_14_3[4]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => ReadFIFO_Read_Ptr(1), B => 
        \APB3_RDATA_1_14_2[4]_net_1\, C => 
        \RX_packet_depth_status\, Y => 
        \APB3_RDATA_1_14_3[4]_net_1\);
    
    \APB3_RDATA_1_d_am_RNO[5]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \APB3_RDATA_1_25_0_wmux_0_Y[5]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \APB3_RDATA_1_25_3[5]_net_1\, Y => N_1675);
    
    \mac_1_byte_3_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_3_reg[4]_net_1\);
    
    \mac_1_byte_2_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type1_reg[3]\);
    
    mac_2_byte_1_reg_en_ret_4 : SLE
      port map(D => un12_mac_2_byte_1_reg_en_16_2, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        N_855_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        un12_mac_2_byte_1_reg_en_16_2_reto);
    
    \RX_packet_depth[5]\ : SLE
      port map(D => \RX_packet_depth_s[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_127_i, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RX_packet_depth[5]_net_1\);
    
    read_reg_en_RNI3S732 : CFG3
      generic map(INIT => x"F7")

      port map(A => N_783, B => \read_reg_en\, C => N_252, Y => 
        APB3_RDATA_1_sn_m21_i_1);
    
    \REG_WRITE_PROC.un13_mac_1_byte_3_reg_en_0_a2_0_a2_1_a2\ : 
        CFG2
      generic map(INIT => x"8")

      port map(A => N_1461, B => \mac_1_byte_3_reg_en\, Y => 
        un13_mac_1_byte_3_reg_en);
    
    \REG_WRITE_PROC.un12_mac_1_byte_1_reg_en_20\ : CFG4
      generic map(INIT => x"FCFA")

      port map(A => mac_1_byte_1_reg_en_reto, B => 
        mac_4_byte_6_reg_en_1_reto, C => N_733_reto, D => 
        N_335_reto, Y => N_732);
    
    \APB3_RDATA_1_ns[7]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \APB3_RDATA_1_29_d_ns[7]_net_1\, B => 
        \APB3_RDATA_1_s[3]_net_1\, C => 
        \APB3_RDATA_1_d_ns[7]_net_1\, Y => \APB3_RDATA_1[7]\);
    
    \mac_3_byte_5_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_5_reg[7]_net_1\);
    
    \APB3_RDATA_1_22[5]\ : CFG4
      generic map(INIT => x"2075")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => RX_FIFO_DOUT(5), D
         => \APB3_RDATA_1_22_1_0[5]_net_1\, Y => N_1650);
    
    mac_4_byte_4_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_356, ALn => N_855_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_4_byte_4_reg_en\);
    
    \mac_2_byte_6_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_6_reg[5]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_2_byte_3_reg_en_0_a2_0_a2_0_a2\ : 
        CFG3
      generic map(INIT => x"20")

      port map(A => \mac_2_byte_3_reg_en\, B => 
        \mac_2_byte_2_reg_en\, C => N_989, Y => 
        un13_mac_2_byte_3_reg_en);
    
    \RX_packet_depth_cry[6]\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \RX_packet_depth[6]_net_1\, B => 
        rx_packet_complt, C => GND_net_1, D => GND_net_1, FCI => 
        \RX_packet_depth_cry[5]_net_1\, S => 
        \RX_packet_depth_s[6]\, Y => OPEN, FCO => 
        \RX_packet_depth_cry[6]_net_1\);
    
    \mac_1_byte_3_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_3_reg[3]_net_1\);
    
    \mac_1_byte_2_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type1_reg[4]\);
    
    \mac_3_byte_5_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_5_reg[4]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_3_byte_3_reg_en_0_a2_1_a2_0_a2\ : 
        CFG3
      generic map(INIT => x"08")

      port map(A => N_989, B => \mac_3_byte_3_reg_en\, C => N_556, 
        Y => un13_mac_3_byte_3_reg_en);
    
    \mac_2_byte_4_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_4_reg[4]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un5_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"1000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_789, D => N_790, Y
         => N_331);
    
    \mac_2_byte_6_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_6_reg[0]_net_1\);
    
    \APB3_RDATA_1_24[7]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_1612, B => CoreAPB3_0_APBmslave0_PADDR(3), 
        C => N_1628, Y => N_1669);
    
    \mac_2_byte_1_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_1_reg[5]_net_1\);
    
    \scratch_pad_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \write_scratch_reg_en\, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \scratch_pad_reg[7]_net_1\);
    
    \APB3_RDATA_1_25_0_0_wmux[6]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_1_byte_5_reg[6]_net_1\, D => 
        \mac_2_byte_1_reg[6]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_25_0_0_y0[6]\, FCO => 
        \APB3_RDATA_1_25_0_0_co0[6]\);
    
    \mac_4_byte_1_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_1_reg[4]_net_1\);
    
    \APB3_RDATA_1_28_RNO[3]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \APB3_RDATA_1_25_0_wmux_0_Y[3]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \APB3_RDATA_1_25_3[3]_net_1\, Y => N_1673);
    
    \mac_3_byte_6_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_6_reg[6]_net_1\);
    
    \APB3_RDATA_1_28_RNO[1]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \APB3_RDATA_1_25_0_wmux_0_Y[1]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \APB3_RDATA_1_25_3[1]_net_1\, Y => N_1671);
    
    \APB3_RDATA_1_am[1]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_1698, B => N_91, C => N_499, Y => 
        \APB3_RDATA_1_am[1]_net_1\);
    
    \APB3_RDATA_1_21_0_wmux_0[7]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_21_0_0_y0[7]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \consumer_type1_reg[7]\, D => \consumer_type2_reg[7]\, 
        FCI => \APB3_RDATA_1_21_0_0_co0[7]\, S => OPEN, Y => 
        N_1644, FCO => OPEN);
    
    \mac_2_byte_1_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_1_reg[2]_net_1\);
    
    \mac_1_byte_2_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type1_reg[2]\);
    
    \APB3_RDATA_1_ns[3]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \APB3_RDATA_1_29_d_ns[3]_net_1\, B => 
        \APB3_RDATA_1_s[3]_net_1\, C => 
        \APB3_RDATA_1_d_ns[3]_net_1\, Y => \APB3_RDATA_1[3]\);
    
    \APB3_RDATA_1_25_0_wmux_0[4]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_25_0_0_y0[4]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_1_reg[4]_net_1\, D => 
        \mac_3_byte_3_reg[4]_net_1\, FCI => 
        \APB3_RDATA_1_25_0_0_co0[4]\, S => OPEN, Y => 
        \APB3_RDATA_1_25_0_wmux_0_Y[4]\, FCO => OPEN);
    
    \APB3_RDATA_1_0_m2_6_2[0]\ : CFG3
      generic map(INIT => x"27")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        \mac_4_byte_2_reg[0]_net_1\, C => N_693, Y => 
        \APB3_RDATA_1_0_m2_6_2[0]_net_1\);
    
    \mac_1_byte_3_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_3_reg[2]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un101_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"2000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(7), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => N_801, Y => N_357);
    
    \mac_4_byte_6_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_6_reg[1]_net_1\);
    
    \mac_4_byte_1_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_1_reg[0]_net_1\);
    
    \mac_3_byte_4_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_4_reg[2]_net_1\);
    
    \mac_2_byte_4_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_4_reg[1]_net_1\);
    
    \mac_2_byte_4_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_4_reg[0]_net_1\);
    
    \mac_4_byte_6_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_6_reg[7]_net_1\);
    
    \RX_packet_depth[1]\ : SLE
      port map(D => \RX_packet_depth_s[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_127_i, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RX_packet_depth[1]_net_1\);
    
    \APB3_RDATA_1_d_am_RNO[6]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \APB3_RDATA_1_25_0_wmux_0_Y[6]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \APB3_RDATA_1_25_3[6]_net_1\, Y => N_1676);
    
    \APB3_RDATA_RNIIKI5[5]\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        \CoreAPB3_0_APBmslave0_PRDATA[5]\, Y => 
        CoreAPB3_0_APBmslave0_PRDATA_m(5));
    
    \mac_3_byte_3_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_3_reg[5]_net_1\);
    
    \APB3_RDATA_1_4[4]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \consumer_type3_reg[4]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \scratch_pad_reg[4]_net_1\, Y => N_1503);
    
    \APB3_RDATA_1_18_i_m2_0_wmux_0[3]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_18_i_m2_0_0_y0[3]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_5_reg[3]_net_1\, D => 
        \mac_4_byte_6_reg[3]_net_1\, FCI => 
        \APB3_RDATA_1_18_i_m2_0_0_co0[3]\, S => OPEN, Y => N_200, 
        FCO => OPEN);
    
    \APB3_RDATA_1_0_m2_1[0]\ : CFG4
      generic map(INIT => x"CFDF")

      port map(A => APB3_RDATA_1_sn_m21_i_1, B => \N_817_i\, C
         => \read_reg_en\, D => \APB3_RDATA_1_0_m2_1_0[0]_net_1\, 
        Y => N_741);
    
    \APB3_RDATA_1_0_m2_0[0]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => N_615, C
         => N_597, Y => N_729);
    
    \mac_1_byte_5_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_5_reg[2]_net_1\);
    
    \APB3_RDATA_1_3[5]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \consumer_type4_reg[5]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_4_reg[5]_net_1\, Y => N_1494);
    
    mac_2_byte_1_reg_en_ret_8 : SLE
      port map(D => \mac_1_byte_1_reg_en\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        N_855_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        mac_1_byte_1_reg_en_reto);
    
    \REG_WRITE_PROC.un13_mac_3_byte_6_reg_en_0_a2_1_a2_0_a2\ : 
        CFG4
      generic map(INIT => x"0040")

      port map(A => \mac_3_byte_5_reg_en\, B => 
        \mac_3_byte_6_reg_en\, C => N_989, D => N_561, Y => 
        un13_mac_3_byte_6_reg_en);
    
    \mac_2_byte_4_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_4_reg[5]_net_1\);
    
    \mac_4_byte_2_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_2_reg[5]_net_1\);
    
    \APB3_RDATA_1_3[7]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \consumer_type4_reg[7]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_4_reg[7]_net_1\, Y => N_1496);
    
    mac_2_byte_1_reg_en_ret_5 : SLE
      port map(D => N_335, CLK => m2s010_som_sb_0_CCC_71MHz, EN
         => VCC_net_1, ALn => N_855_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        N_335_reto);
    
    \mac_3_byte_5_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_5_reg[5]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_4_byte_5_reg_en_0_a2_0_a2_0_o2\ : 
        CFG3
      generic map(INIT => x"FE")

      port map(A => \mac_4_byte_4_reg_en\, B => 
        \mac_4_byte_3_reg_en\, C => \mac_4_byte_2_reg_en\, Y => 
        N_576);
    
    \APB3_RDATA_1_29_d_am[7]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_1644, B => N_204, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => 
        \APB3_RDATA_1_29_d_am[7]_net_1\);
    
    \APB3_RDATA_1_bm[1]\ : CFG4
      generic map(INIT => x"8F88")

      port map(A => N_1655, B => N_1350, C => \N_817_i\, D => 
        \APB3_RDATA_1_bm_1[1]_net_1\, Y => 
        \APB3_RDATA_1_bm[1]_net_1\);
    
    \mac_2_byte_6_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_6_reg[3]_net_1\);
    
    \mac_4_byte_1_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_1_reg[6]_net_1\);
    
    mac_2_byte_2_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_342, ALn => N_855_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_2_byte_2_reg_en\);
    
    \APB3_RDATA_1_24_i_m3_1_wmux_0[1]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_24_i_m3_1_2_y0[1]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \consumer_type1_reg[9]\, D => \mac_3_byte_5_reg[1]_net_1\, 
        FCI => \APB3_RDATA_1_24_i_m3_1_2_co0[1]\, S => OPEN, Y
         => N_497, FCO => OPEN);
    
    \N_41_i\ : CFG3
      generic map(INIT => x"A8")

      port map(A => N_535, B => rx_crc_HighByte_en, C => 
        RX_FIFO_DIN_pipe_0, Y => N_41_i);
    
    \APB3_RDATA[4]\ : SLE
      port map(D => \APB3_RDATA_1[4]\, CLK => N_41_mux, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        \CoreAPB3_0_APBmslave0_PRDATA[4]\);
    
    mac_3_byte_4_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_350, ALn => N_855_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_3_byte_4_reg_en\);
    
    \APB3_RDATA_1_25_3[4]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_50, B => CoreAPB3_0_APBmslave0_PADDR(3), C
         => N_1493, Y => \APB3_RDATA_1_25_3[4]_net_1\);
    
    \APB3_RDATA_RNIEGI5[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        \CoreAPB3_0_APBmslave0_PRDATA[1]\, Y => 
        CoreAPB3_0_APBmslave0_PRDATA_m(1));
    
    control_reg_en_ret : SLE
      port map(D => N_734, CLK => m2s010_som_sb_0_CCC_71MHz, EN
         => VCC_net_1, ALn => N_855_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        N_743);
    
    \WRITE_REGISTER_ENABLE_PROC.un53_apb3_addr_0_a2_0_a2\ : CFG4
      generic map(INIT => x"2000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_789, D => N_795, Y
         => N_345);
    
    \APB3_RDATA_1_25_3[1]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => N_137, C
         => N_1086, Y => \APB3_RDATA_1_25_3[1]_net_1\);
    
    APB3_RDATA_1_sn_m21_i_a2 : CFG4
      generic map(INIT => x"C040")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(5), Y => N_252);
    
    iup_EOP : SLE
      port map(D => un117_apb3_addr, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \iup_EOP\);
    
    \mac_4_byte_6_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_6_reg[4]_net_1\);
    
    \mac_3_byte_1_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_1_reg[1]_net_1\);
    
    \iAPB3_READY_RNIV0ML[0]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \iAPB3_READYrs[0]\, B => un5_apb3_rst_rs, C
         => long_reset_set, Y => \iAPB3_READY[0]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_4_byte_4_reg_en_0_a2_0_a2_0_a2_1\ : 
        CFG4
      generic map(INIT => x"0100")

      port map(A => \mac_4_byte_3_reg_en\, B => 
        \mac_4_byte_2_reg_en\, C => N_742, D => 
        \mac_4_byte_4_reg_en\, Y => 
        un13_mac_4_byte_4_reg_en_0_a2_0_a2_0_a2_1);
    
    \mac_3_byte_5_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_5_reg[1]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_3_byte_2_reg_en_0_a2_1_a2_0_a2\ : 
        CFG4
      generic map(INIT => x"0040")

      port map(A => \mac_3_byte_1_reg_en\, B => 
        \mac_3_byte_2_reg_en\, C => N_989, D => N_549, Y => 
        un13_mac_3_byte_2_reg_en);
    
    \APB3_RDATA_1_24[5]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_1610, B => CoreAPB3_0_APBmslave0_PADDR(3), 
        C => N_1626, Y => N_1667);
    
    \mac_1_byte_1_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_1_reg[4]_net_1\);
    
    \mac_2_byte_1_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_1_reg[7]_net_1\);
    
    \APB3_RDATA_1_19_0_0_wmux[3]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \i_int_mask_reg[3]_net_1\, D => 
        \mac_1_byte_3_reg[3]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_19_0_0_y0[3]\, FCO => 
        \APB3_RDATA_1_19_0_0_co0[3]\);
    
    \REG_WRITE_PROC.un12_control_reg_en_0\ : CFG4
      generic map(INIT => x"FFCA")

      port map(A => \write_scratch_reg_en\, B => 
        mac_4_byte_6_reg_en_1, C => N_329, D => N_3, Y => N_734);
    
    APB3_RDATA_1_sn_m13_0_o2_i_a2 : CFG2
      generic map(INIT => x"4")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_757);
    
    mac_2_byte_5_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_345, ALn => N_855_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_2_byte_5_reg_en\);
    
    \WRITE_REGISTER_ENABLE_PROC.un49_apb3_addr_0_a2\ : CFG3
      generic map(INIT => x"80")

      port map(A => N_795, B => N_791, C => N_789, Y => N_344);
    
    \APB3_RDATA_1[5]\ : CFG4
      generic map(INIT => x"F780")

      port map(A => N_78, B => N_91, C => N_1692, D => 
        \APB3_RDATA_1_d_ns[5]_net_1\, Y => 
        \APB3_RDATA_1[5]_net_1\);
    
    \APB3_RDATA_1_21_0_wmux_0[5]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_21_0_0_y0[5]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \consumer_type1_reg[5]\, D => \consumer_type2_reg[5]\, 
        FCI => \APB3_RDATA_1_21_0_0_co0[5]\, S => OPEN, Y => 
        N_1642, FCO => OPEN);
    
    \RX_packet_depth[7]\ : SLE
      port map(D => \RX_packet_depth_s[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_127_i, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RX_packet_depth[7]_net_1\);
    
    \mac_2_byte_2_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type4_reg[0]\);
    
    \mac_1_byte_6_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type3_reg[1]\);
    
    \mac_1_byte_1_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type1_reg[8]\);
    
    \mac_4_byte_6_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_6_reg[2]_net_1\);
    
    \i_int_mask_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_1354_i, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \i_int_mask_reg[5]_net_1\);
    
    read_reg_en_RNINPBI4 : CFG4
      generic map(INIT => x"FFFD")

      port map(A => \read_reg_en\, B => m30_0_0, C => \N_817_i\, 
        D => N_234, Y => N_41_mux);
    
    m14_0_a3_1 : CFG3
      generic map(INIT => x"02")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(7), C => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => N_353_1);
    
    \iAPB3_READY_RNID89P[1]\ : CFG2
      generic map(INIT => x"D")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        CoreAPB3_0_APBmslave0_PREADY, Y => 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i);
    
    \mac_1_byte_6_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type3_reg[7]\);
    
    \WRITE_REGISTER_ENABLE_PROC.un45_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"1000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_789, D => N_795, Y
         => N_343);
    
    \APB3_RDATA_1_0_m2_3_bm[0]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \consumer_type4_reg[0]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_4_reg[0]_net_1\, Y => 
        \APB3_RDATA_1_0_m2_3_bm[0]_net_1\);
    
    \mac_3_byte_4_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_4_reg[7]_net_1\);
    
    \mac_3_byte_4_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_4_reg[6]_net_1\);
    
    \mac_3_byte_3_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_3_reg[6]_net_1\);
    
    \APB3_RDATA_1_am_1_RNO[4]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \APB3_RDATA_1_25_0_wmux_0_Y[4]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \APB3_RDATA_1_25_3[4]_net_1\, Y => N_1674);
    
    \APB3_RDATA_1_14_0_0_wmux[2]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => ReadFIFO_Read_Ptr(0), B => 
        ReadFIFO_Read_Ptr(1), C => N_651, D => N_658, FCI => 
        VCC_net_1, S => OPEN, Y => \APB3_RDATA_1_14_0_0_y0[2]\, 
        FCO => \APB3_RDATA_1_14_0_0_co0[2]\);
    
    \APB3_RDATA_1_21_0_0_wmux[6]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_2_byte_4_reg[6]_net_1\, D => 
        \mac_2_byte_6_reg[6]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_21_0_0_y0[6]\, FCO => 
        \APB3_RDATA_1_21_0_0_co0[6]\);
    
    \APB3_RDATA_1_0_m2_6[0]\ : CFG4
      generic map(INIT => x"555C")

      port map(A => \APB3_RDATA_1_0_m2_6_2[0]_net_1\, B => N_678, 
        C => CoreAPB3_0_APBmslave0_PADDR(4), D => 
        CoreAPB3_0_APBmslave0_PADDR(5), Y => N_586);
    
    \APB3_RDATA[1]\ : SLE
      port map(D => \APB3_RDATA_1[1]\, CLK => N_41_mux, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        \CoreAPB3_0_APBmslave0_PRDATA[1]\);
    
    \APB3_RDATA_1_0_m2_2_3[0]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => N_697, C
         => N_698, Y => \APB3_RDATA_1_0_m2_2_3[0]_net_1\);
    
    \APB3_RDATA_1_25_3[7]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_1087, B => CoreAPB3_0_APBmslave0_PADDR(3), 
        C => N_1496, Y => \APB3_RDATA_1_25_3[7]_net_1\);
    
    \APB3_RDATA_1_18_i_m2_0_wmux_0[7]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_18_i_m2_0_0_y0[7]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_5_reg[7]_net_1\, D => 
        \mac_4_byte_6_reg[7]_net_1\, FCI => 
        \APB3_RDATA_1_18_i_m2_0_0_co0[7]\, S => OPEN, Y => N_204, 
        FCO => OPEN);
    
    \i_int_mask_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_1354_i, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \i_int_mask_reg[2]_net_1\);
    
    read_reg_en_RNI0LK33 : CFG4
      generic map(INIT => x"FFEF")

      port map(A => APB3_RDATA_1_sn_m26_i_1, B => \N_817_i\, C
         => \read_reg_en\, D => N_785, Y => N_91);
    
    \APB3_RDATA_1_4[3]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \consumer_type3_reg[3]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \scratch_pad_reg[3]_net_1\, Y => N_1502);
    
    \mac_2_byte_3_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_3_reg[0]_net_1\);
    
    \APB3_RDATA_1_25_0_wmux_0[1]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_25_0_0_y0[1]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_1_reg[1]_net_1\, D => 
        \mac_3_byte_3_reg[1]_net_1\, FCI => 
        \APB3_RDATA_1_25_0_0_co0[1]\, S => OPEN, Y => 
        \APB3_RDATA_1_25_0_wmux_0_Y[1]\, FCO => OPEN);
    
    \REG_WRITE_PROC.un13_mac_4_byte_2_reg_en_0_a2_3_a2_2_o2\ : 
        CFG4
      generic map(INIT => x"FFFE")

      port map(A => \mac_4_byte_1_reg_en\, B => N_1357, C => 
        un13_mac_4_byte_1_reg_en_0_a2_0_a2_0_o2_0, D => N_556, Y
         => N_570);
    
    \WRITE_REGISTER_ENABLE_PROC.un65_apb3_addr_0_a2_0\ : CFG2
      generic map(INIT => x"4")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => N_791);
    
    \mac_1_byte_2_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type1_reg[5]\);
    
    \APB3_RDATA_1_17_i_m2_0_wmux_0[2]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_17_i_m2_0_0_y0[2]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_1_byte_1_reg[2]_net_1\, D => 
        \mac_3_byte_5_reg[2]_net_1\, FCI => 
        \APB3_RDATA_1_17_i_m2_0_0_co0[2]\, S => OPEN, Y => N_1342, 
        FCO => OPEN);
    
    \APB3_RDATA_1_14_0_wmux_0[3]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_14_0_0_y0[3]\, B => 
        ReadFIFO_Read_Ptr(1), C => N_666, D => N_673, FCI => 
        \APB3_RDATA_1_14_0_0_co0[3]\, S => OPEN, Y => 
        \APB3_RDATA_1_14_0_wmux_0_Y[3]\, FCO => OPEN);
    
    \mac_3_byte_4_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_4_reg[3]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un33_apb3_addr_0_a2\ : CFG3
      generic map(INIT => x"80")

      port map(A => N_793, B => N_795, C => N_791, Y => N_340);
    
    \mac_4_byte_2_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_2_reg[6]_net_1\);
    
    \APB3_RDATA_1_14_0_wmux_0[2]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_14_0_0_y0[2]\, B => 
        ReadFIFO_Read_Ptr(1), C => N_665, D => N_672, FCI => 
        \APB3_RDATA_1_14_0_0_co0[2]\, S => OPEN, Y => 
        \APB3_RDATA_1_14_0_wmux_0_Y[2]\, FCO => OPEN);
    
    \mac_4_byte_2_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_2_reg[1]_net_1\);
    
    mac_4_byte_2_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_354, ALn => N_855_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_4_byte_2_reg_en\);
    
    \mac_3_byte_3_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_3_reg[4]_net_1\);
    
    \mac_3_byte_2_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_2_reg[3]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.mac_4_byte_6_reg_en_1\ : CFG2
      generic map(INIT => x"2")

      port map(A => \iAPB3_READY[0]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PREADY, Y => mac_4_byte_6_reg_en_1);
    
    \APB3_RDATA_1_15[4]\ : CFG4
      generic map(INIT => x"AA30")

      port map(A => \mac_4_byte_2_reg[4]_net_1\, B => 
        \i_int_mask_reg[4]_net_1\, C => tx_FIFO_OVERFLOW_int, D
         => CoreAPB3_0_APBmslave0_PADDR(3), Y => N_1593);
    
    \APB3_RDATA_1_14_0_wmux_0[4]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_14_0_0_y0[4]\, B => 
        ReadFIFO_Read_Ptr(1), C => N_667, D => N_674, FCI => 
        \APB3_RDATA_1_14_0_0_co0[4]\, S => OPEN, Y => 
        \APB3_RDATA_1_14_0_wmux_0_Y[4]\, FCO => OPEN);
    
    \mac_1_byte_1_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_1_reg[6]_net_1\);
    
    \RX_packet_depth[4]\ : SLE
      port map(D => \RX_packet_depth_s[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_127_i, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RX_packet_depth[4]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un13_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"1000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_789, D => N_802, Y
         => N_335);
    
    \mac_4_byte_1_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_1_reg[3]_net_1\);
    
    \APB3_RDATA_1_25_0_0_wmux[1]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \consumer_type3_reg[9]\, D => \consumer_type4_reg[9]\, 
        FCI => VCC_net_1, S => OPEN, Y => 
        \APB3_RDATA_1_25_0_0_y0[1]\, FCO => 
        \APB3_RDATA_1_25_0_0_co0[1]\);
    
    \iAPB3_READY[1]\ : SLE
      port map(D => \iAPB3_READY[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        un5_apb3_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAPB3_0_APBmslave0_PREADYrs);
    
    \REG_WRITE_PROC.un13_mac_1_byte_6_reg_en_0_a2_1_a2_1_a2\ : 
        CFG3
      generic map(INIT => x"80")

      port map(A => N_1461, B => \mac_1_byte_6_reg_en\, C => 
        N_1457, Y => un13_mac_1_byte_6_reg_en);
    
    \mac_2_byte_5_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_5_reg[3]_net_1\);
    
    \APB3_RDATA_1_29_d_bm_1_0[7]\ : CFG3
      generic map(INIT => x"47")

      port map(A => \consumer_type3_reg[7]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \scratch_pad_reg[7]_net_1\, Y => 
        \APB3_RDATA_1_29_d_bm_1_0[7]_net_1\);
    
    \control_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => control_reg_13, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => rx_FIFO_rst_reg);
    
    \APB3_RDATA_1_20_i_m3_0_i_m2[1]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \consumer_type4_reg[1]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_4_reg[1]_net_1\, Y => N_137);
    
    \APB3_RDATA_1_18_i_m2_0_0_wmux[5]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_3_reg[5]_net_1\, D => 
        \mac_4_byte_4_reg[5]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_18_i_m2_0_0_y0[5]\, FCO => 
        \APB3_RDATA_1_18_i_m2_0_0_co0[5]\);
    
    \APB3_RDATA_1_ns[1]\ : CFG4
      generic map(INIT => x"F870")

      port map(A => N_91, B => N_78, C => 
        \APB3_RDATA_1_am[1]_net_1\, D => 
        \APB3_RDATA_1_bm[1]_net_1\, Y => \APB3_RDATA_1[1]\);
    
    \REG_WRITE_PROC.un13_mac_3_byte_4_reg_en_0_a2_1_a2_0_a2\ : 
        CFG4
      generic map(INIT => x"0040")

      port map(A => \mac_3_byte_3_reg_en\, B => 
        \mac_3_byte_4_reg_en\, C => N_989, D => N_556, Y => 
        un13_mac_3_byte_4_reg_en);
    
    \mac_3_byte_3_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_3_reg[3]_net_1\);
    
    \mac_3_byte_2_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_2_reg[4]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_2_byte_6_reg_en_0_a2_1_a2_0_a2\ : 
        CFG4
      generic map(INIT => x"0040")

      port map(A => \mac_2_byte_5_reg_en\, B => 
        \mac_2_byte_6_reg_en\, C => N_989, D => N_547, Y => 
        un13_mac_2_byte_6_reg_en);
    
    iRX_FIFO_rd_en_RNO : CFG1
      generic map(INIT => "01")

      port map(A => \iAPB3_READY[0]_net_1\, Y => 
        \iAPB3_READY_i[0]\);
    
    \APB3_RDATA_1_0_m2_8_2_wmux[0]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_2_byte_4_reg[0]_net_1\, D => 
        \mac_2_byte_6_reg[0]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_0_m2_8_2_y0[0]\, FCO => 
        \APB3_RDATA_1_0_m2_8_2_co0[0]\);
    
    \mac_1_byte_6_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type3_reg[4]\);
    
    \APB3_RDATA_1_25_0_wmux_0[6]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_25_0_0_y0[6]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_1_reg[6]_net_1\, D => 
        \mac_3_byte_3_reg[6]_net_1\, FCI => 
        \APB3_RDATA_1_25_0_0_co0[6]\, S => OPEN, Y => 
        \APB3_RDATA_1_25_0_wmux_0_Y[6]\, FCO => OPEN);
    
    \APB3_RDATA_1_18_i_m2_0_0_wmux[4]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_3_reg[4]_net_1\, D => 
        \mac_4_byte_4_reg[4]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_18_i_m2_0_0_y0[4]\, FCO => 
        \APB3_RDATA_1_18_i_m2_0_0_co0[4]\);
    
    \APB3_RDATA_1_14_4_0_wmux[1]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => ReadFIFO_Read_Ptr(0), B => 
        ReadFIFO_Read_Ptr(1), C => RX_FIFO_DOUT_0_0, D => 
        RX_FIFO_DOUT_1_0, FCI => VCC_net_1, S => OPEN, Y => 
        \APB3_RDATA_1_14_4_0_y0[1]\, FCO => 
        \APB3_RDATA_1_14_4_0_co0[1]\);
    
    \mac_2_byte_5_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_5_reg[6]_net_1\);
    
    \RX_packet_depth_cry[2]\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \RX_packet_depth[2]_net_1\, B => 
        rx_packet_complt, C => GND_net_1, D => GND_net_1, FCI => 
        \RX_packet_depth_cry[1]_net_1\, S => 
        \RX_packet_depth_s[2]\, Y => OPEN, FCO => 
        \RX_packet_depth_cry[2]_net_1\);
    
    \APB3_RDATA_1_ns[2]\ : CFG4
      generic map(INIT => x"F870")

      port map(A => N_91, B => N_78, C => 
        \APB3_RDATA_1_am[2]_net_1\, D => 
        \APB3_RDATA_1_bm[2]_net_1\, Y => \APB3_RDATA_1[2]\);
    
    
        \WRITE_REGISTER_ENABLE_PROC.un9_apb3_addr_0_a2_0_a2_0_0_a2_RNIDDPT\ : 
        CFG4
      generic map(INIT => x"2EAA")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(7), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => N_790, D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => N_783);
    
    \RX_packet_depth[0]\ : SLE
      port map(D => \RX_packet_depth_s[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_127_i, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RX_packet_depth[0]_net_1\);
    
    \mac_4_byte_6_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_6_reg[5]_net_1\);
    
    N_817_i : CFG4
      generic map(INIT => x"CC4C")

      port map(A => CoreAPB3_0_APBmslave0_PENABLE, B => 
        long_reset, C => CoreAPB3_0_APBmslave0_PSELx, D => 
        CoreAPB3_0_APBmslave0_PWRITE, Y => \N_817_i\);
    
    mac_1_byte_4_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_338, ALn => N_855_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_1_byte_4_reg_en\);
    
    read_reg_en_RNI3OAV1 : CFG2
      generic map(INIT => x"E")

      port map(A => \N_817_i\, B => APB3_RDATA_1_sn_m12_i_0_0, Y
         => N_1350);
    
    mac_4_byte_5_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_357, ALn => N_855_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_4_byte_5_reg_en\);
    
    APB3_RDATA_1_27_10 : CFG2
      generic map(INIT => x"B")

      port map(A => \N_817_i\, B => \read_reg_en\, Y => 
        \APB3_RDATA_1_27_10\);
    
    \mac_4_byte_4_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_4_reg[4]_net_1\);
    
    \APB3_RDATA_1_27_1[5]\ : CFG4
      generic map(INIT => x"44F0")

      port map(A => APB3_RDATA_1_sn_m12_i_0, B => N_1594, C => 
        N_1650, D => APB3_RDATA_1_sn_m12_i_0_0, Y => 
        \APB3_RDATA_1_27_1[5]_net_1\);
    
    \mac_4_byte_6_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_6_reg[0]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un9_apb3_addr_0_a2_0_a2_0_0_a2\ : 
        CFG2
      generic map(INIT => x"1")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), Y => N_790);
    
    \APB3_RDATA_1_27[6]\ : CFG3
      generic map(INIT => x"BA")

      port map(A => \APB3_RDATA_1_27_10\, B => \N_817_i\, C => 
        \APB3_RDATA_1_27_1[6]_net_1\, Y => N_1693);
    
    \APB3_RDATA_1_15[5]\ : CFG4
      generic map(INIT => x"AA30")

      port map(A => \mac_4_byte_2_reg[5]_net_1\, B => 
        \i_int_mask_reg[5]_net_1\, C => tx_FIFO_UNDERRUN_int, D
         => CoreAPB3_0_APBmslave0_PADDR(3), Y => N_1594);
    
    \mac_3_byte_2_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_2_reg[2]_net_1\);
    
    \APB3_RDATA_1_29_d_bm[3]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => N_1502, 
        C => N_1584, Y => \APB3_RDATA_1_29_d_bm[3]_net_1\);
    
    \mac_4_byte_1_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_1_reg[5]_net_1\);
    
    \mac_1_byte_6_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type3_reg[2]\);
    
    \APB3_RDATA_1_29_d_ns[7]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \APB3_RDATA_1_29_d_bm[7]_net_1\, B => N_78, C
         => \APB3_RDATA_1_29_d_am[7]_net_1\, Y => 
        \APB3_RDATA_1_29_d_ns[7]_net_1\);
    
    \mac_3_byte_3_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_3_reg[2]_net_1\);
    
    \APB3_RDATA_1_27_1[6]\ : CFG4
      generic map(INIT => x"44F0")

      port map(A => APB3_RDATA_1_sn_m12_i_0, B => N_1595, C => 
        N_1651, D => APB3_RDATA_1_sn_m12_i_0_0, Y => 
        \APB3_RDATA_1_27_1[6]_net_1\);
    
    mac_2_byte_1_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_341, ALn => N_855_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_2_byte_1_reg_en\);
    
    \WRITE_REGISTER_ENABLE_PROC.un61_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"1000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_793, D => N_796, Y
         => N_347);
    
    \APB3_RDATA_RNIGII5[3]\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        \CoreAPB3_0_APBmslave0_PRDATA[3]\, Y => 
        CoreAPB3_0_APBmslave0_PRDATA_m(3));
    
    \APB3_RDATA_1_23[4]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \N_817_i\, B => N_1593, C => 
        APB3_RDATA_1_sn_m12_i_0, Y => N_1658);
    
    \REG_WRITE_PROC.un13_mac_4_byte_6_reg_en_0_a2_4_a2_3_a2_0\ : 
        CFG4
      generic map(INIT => x"0010")

      port map(A => \mac_2_byte_1_reg_en\, B => 
        \mac_1_byte_6_reg_en\, C => N_1457, D => N_570, Y => 
        N_1337);
    
    \APB3_RDATA_1_21_0_wmux_0[4]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_21_0_0_y0[4]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \consumer_type1_reg[4]\, D => \consumer_type2_reg[4]\, 
        FCI => \APB3_RDATA_1_21_0_0_co0[4]\, S => OPEN, Y => 
        N_1641, FCO => OPEN);
    
    \mac_4_byte_1_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_1_reg[2]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un81_apb3_addr_0_a2\ : CFG3
      generic map(INIT => x"80")

      port map(A => N_796, B => N_791, C => N_789, Y => N_352);
    
    \mac_3_byte_5_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_5_reg[2]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_4_byte_1_reg_en_0_a2_0_a2_0_a2\ : 
        CFG4
      generic map(INIT => x"0040")

      port map(A => N_1357, B => \mac_4_byte_1_reg_en\, C => 
        N_989, D => N_561, Y => un13_mac_4_byte_1_reg_en);
    
    \APB3_RDATA_1_14_0_0_wmux[4]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => ReadFIFO_Read_Ptr(0), B => 
        ReadFIFO_Read_Ptr(1), C => N_653, D => N_660, FCI => 
        VCC_net_1, S => OPEN, Y => \APB3_RDATA_1_14_0_0_y0[4]\, 
        FCO => \APB3_RDATA_1_14_0_0_co0[4]\);
    
    \mac_4_byte_4_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_4_reg[1]_net_1\);
    
    \APB3_RDATA_1_0_m2_3_ns[0]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \APB3_RDATA_1_0_m2_3_am[0]_net_1\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \APB3_RDATA_1_0_m2_3_bm[0]_net_1\, Y => N_615);
    
    \APB3_RDATA_1_0[0]\ : CFG4
      generic map(INIT => x"FDA8")

      port map(A => N_91, B => N_741, C => 
        \APB3_RDATA_1_0_a2_1[0]\, D => N_729, Y => 
        \APB3_RDATA_1[0]\);
    
    write_scratch_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_329, ALn => N_855_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \write_scratch_reg_en\);
    
    \mac_4_byte_4_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_4_reg[0]_net_1\);
    
    control_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_331, ALn => N_855_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \control_reg_en\);
    
    \APB3_RDATA_1_d_am[6]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => N_1668, B => N_757, C => N_1676, Y => 
        \APB3_RDATA_1_d_am[6]_net_1\);
    
    mac_4_byte_1_reg_en_RNO : CFG4
      generic map(INIT => x"1000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(1), B => 
        CoreAPB3_0_APBmslave0_PADDR(0), C => N_353_1, D => 
        \m14_0_a3_1\, Y => N_353);
    
    \mac_2_byte_2_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type4_reg[7]\);
    
    \mac_1_byte_2_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type1_reg[6]\);
    
    \mac_1_byte_2_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type1_reg[1]\);
    
    \APB3_RDATA_1_0_m2_0_RNO[0]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => 
        \APB3_RDATA_1_0_m2_2_wmux_0_Y[0]\, C => 
        \APB3_RDATA_1_0_m2_2_3[0]_net_1\, Y => N_597);
    
    \REG_WRITE_PROC.un13_mac_3_byte_5_reg_en_0_a2_1_a2_0_a2\ : 
        CFG4
      generic map(INIT => x"0040")

      port map(A => un13_mac_4_byte_1_reg_en_0_a2_0_a2_0_o2_0, B
         => \mac_3_byte_5_reg_en\, C => N_989, D => N_556, Y => 
        un13_mac_3_byte_5_reg_en);
    
    mac_3_byte_2_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_348, ALn => N_855_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_3_byte_2_reg_en\);
    
    write_reg_en : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => N_855_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \write_reg_en\);
    
    
        \WRITE_REGISTER_ENABLE_PROC.un9_apb3_addr_0_a2_0_a2_0_0_a2_RNIK11J2\ : 
        CFG3
      generic map(INIT => x"F4")

      port map(A => N_353_1, B => N_801, C => N_789, Y => m30_0_0);
    
    \mac_1_byte_1_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_1_reg[3]_net_1\);
    
    \mac_4_byte_4_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_4_reg[5]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_1_byte_2_reg_en_0_a2_0_a2_2_a2\ : 
        CFG3
      generic map(INIT => x"20")

      port map(A => \mac_1_byte_2_reg_en\, B => 
        \mac_1_byte_1_reg_en\, C => N_1455, Y => 
        un13_mac_1_byte_2_reg_en);
    
    \APB3_RDATA_1_22_1_0[5]\ : CFG3
      generic map(INIT => x"47")

      port map(A => \consumer_type3_reg[5]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \scratch_pad_reg[5]_net_1\, Y => 
        \APB3_RDATA_1_22_1_0[5]_net_1\);
    
    \RX_PACKET_DEPTH_STATUS_PROC.un1_RX_packet_depthlto7_5\ : 
        CFG4
      generic map(INIT => x"0001")

      port map(A => \RX_packet_depth[3]_net_1\, B => 
        \RX_packet_depth[2]_net_1\, C => 
        \RX_packet_depth[1]_net_1\, D => 
        \RX_packet_depth[0]_net_1\, Y => 
        un1_RX_packet_depthlto7_5);
    
    \REG_WRITE_PROC.un12_int_mask_reg_en\ : CFG4
      generic map(INIT => x"FAFC")

      port map(A => mac_4_byte_6_reg_en_1, B => \int_mask_reg_en\, 
        C => N_734, D => N_333, Y => N_733);
    
    \i_int_mask_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_1354_i, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \i_int_mask_reg[6]_net_1\);
    
    \mac_2_byte_3_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_3_reg[7]_net_1\);
    
    \iAPB3_READY_RNI02ML[1]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => CoreAPB3_0_APBmslave0_PREADYrs, B => 
        un5_apb3_rst_rs, C => long_reset_set, Y => 
        CoreAPB3_0_APBmslave0_PREADY);
    
    \REG_WRITE_PROC.un13_mac_3_byte_4_reg_en_0_a2_1_a2_0_o2\ : 
        CFG3
      generic map(INIT => x"FE")

      port map(A => \mac_3_byte_2_reg_en\, B => 
        \mac_3_byte_1_reg_en\, C => N_549, Y => N_556);
    
    \APB3_RDATA_1_17_0_wmux_0[7]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_17_0_0_y0[7]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_1_byte_1_reg[7]_net_1\, D => 
        \mac_3_byte_5_reg[7]_net_1\, FCI => 
        \APB3_RDATA_1_17_0_0_co0[7]\, S => OPEN, Y => N_1612, FCO
         => OPEN);
    
    \mac_4_byte_6_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_6_reg[3]_net_1\);
    
    \mac_2_byte_3_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_3_reg[1]_net_1\);
    
    \RX_PACKET_DEPTH_STATUS_PROC.rx_packet_depth_status2\ : CFG4
      generic map(INIT => x"7707")

      port map(A => un1_RX_packet_depthlto7_4, B => 
        un1_RX_packet_depthlto7_5, C => \iup_EOP\, D => 
        \RX_packet_depth_status\, Y => rx_packet_depth_status2);
    
    \APB3_RDATA_1_18_i_m2_0_0_wmux[2]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_3_reg[2]_net_1\, D => 
        \mac_4_byte_4_reg[2]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_18_i_m2_0_0_y0[2]\, FCO => 
        \APB3_RDATA_1_18_i_m2_0_0_co0[2]\);
    
    \WRITE_REGISTER_ENABLE_PROC.un89_apb3_addr_0_a2_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_789, D => N_796, Y
         => N_354);
    
    \mac_1_byte_6_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type3_reg[5]\);
    
    \REG_WRITE_PROC.un13_mac_1_byte_1_reg_en_0_a2_2_a2_0_a2_0\ : 
        CFG3
      generic map(INIT => x"01")

      port map(A => \control_reg_en\, B => \write_scratch_reg_en\, 
        C => \int_mask_reg_en\, Y => N_1455);
    
    mac_2_byte_1_reg_en_ret_7 : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        N_855_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        mac_4_byte_6_reg_en_1_reto);
    
    \up_EOP_sync[1]\ : SLE
      port map(D => \up_EOP_sync[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \up_EOP_sync[1]_net_1\);
    
    read_reg_en_RNIJAKE : CFG2
      generic map(INIT => x"7")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \read_reg_en\, Y => APB3_RDATA_1_sn_m12_i_0);
    
    \mac_3_byte_1_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_1_reg[4]_net_1\);
    
    \i_int_mask_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_1354_i, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \i_int_mask_reg[0]_net_1\);
    
    \APB3_RDATA_1_22_1_0[6]\ : CFG3
      generic map(INIT => x"47")

      port map(A => \consumer_type3_reg[6]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \scratch_pad_reg[6]_net_1\, Y => 
        \APB3_RDATA_1_22_1_0[6]_net_1\);
    
    APB3_RDATA_1_23_1 : CFG3
      generic map(INIT => x"0B")

      port map(A => \N_817_i\, B => \read_reg_en\, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => \APB3_RDATA_1_23_1\);
    
    \APB3_RDATA_1_25_0_0_wmux[3]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_1_byte_5_reg[3]_net_1\, D => 
        \mac_2_byte_1_reg[3]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_25_0_0_y0[3]\, FCO => 
        \APB3_RDATA_1_25_0_0_co0[3]\);
    
    \mac_1_byte_4_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type2_reg[4]\);
    
    \APB3_RDATA_1_14_3[3]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => ReadFIFO_Read_Ptr(1), B => 
        \APB3_RDATA_1_14_2[3]_net_1\, C => TX_FIFO_Full, Y => 
        \APB3_RDATA_1_14_3[3]_net_1\);
    
    mac_3_byte_5_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_351, ALn => N_855_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_3_byte_5_reg_en\);
    
    \APB3_RDATA_1_28[7]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => N_1669, B => N_757, C => N_1677, Y => N_1704);
    
    \mac_1_byte_6_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type3_reg[0]\);
    
    \APB3_RDATA[0]\ : SLE
      port map(D => \APB3_RDATA_1[0]\, CLK => N_41_mux, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        \CoreAPB3_0_APBmslave0_PRDATA[0]\);
    
    \REG_WRITE_PROC.un13_mac_2_byte_1_reg_en_0_a2_2_a2_1_a2_1\ : 
        CFG3
      generic map(INIT => x"10")

      port map(A => \mac_1_byte_2_reg_en\, B => 
        \mac_1_byte_1_reg_en\, C => N_1455, Y => N_1461);
    
    \APB3_RDATA_1_14_4_wmux_2[1]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_14_4_y0_0[1]\, B => 
        ReadFIFO_Read_Ptr(1), C => iRX_FIFO_Full(2), D => 
        iRX_FIFO_Full(3), FCI => \APB3_RDATA_1_14_4_co0_0[1]\, S
         => OPEN, Y => \APB3_RDATA_1_14_4_0_y3[1]\, FCO => 
        \APB3_RDATA_1_14_4_co1_0[1]\);
    
    \REG_WRITE_PROC.un13_mac_2_byte_4_reg_en_0_a2_1_a2_0_a2\ : 
        CFG4
      generic map(INIT => x"0200")

      port map(A => \mac_2_byte_4_reg_en\, B => 
        \mac_2_byte_3_reg_en\, C => \mac_2_byte_2_reg_en\, D => 
        N_989, Y => un13_mac_2_byte_4_reg_en);
    
    \mac_1_byte_1_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_1_reg[5]_net_1\);
    
    \APB3_RDATA_1_22[6]\ : CFG4
      generic map(INIT => x"2075")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => RX_FIFO_DOUT(6), D
         => \APB3_RDATA_1_22_1_0[6]_net_1\, Y => N_1651);
    
    mac_4_byte_1_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_353, ALn => N_855_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_4_byte_1_reg_en\);
    
    \mac_3_byte_6_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_6_reg[1]_net_1\);
    
    \mac_3_byte_1_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_1_reg[0]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un37_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"2000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_793, D => N_795, Y
         => N_341);
    
    \scratch_pad_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \write_scratch_reg_en\, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \scratch_pad_reg[6]_net_1\);
    
    \mac_4_byte_1_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_1_reg[7]_net_1\);
    
    \APB3_RDATA_1_bm_1[1]\ : CFG4
      generic map(INIT => x"4540")

      port map(A => APB3_RDATA_1_sn_m12_i_0_0, B => N_110, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => N_490, Y => 
        \APB3_RDATA_1_bm_1[1]_net_1\);
    
    \REG_WRITE_PROC.un12_mac_2_byte_1_reg_en_16_0\ : CFG4
      generic map(INIT => x"FFCA")

      port map(A => \mac_1_byte_5_reg_en\, B => 
        mac_4_byte_6_reg_en_1, C => N_339, D => N_10, Y => 
        un12_mac_2_byte_1_reg_en_16_0);
    
    \mac_3_byte_6_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_6_reg[7]_net_1\);
    
    \APB3_RDATA_1_25_0_0_wmux[4]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_1_byte_5_reg[4]_net_1\, D => 
        \mac_2_byte_1_reg[4]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_25_0_0_y0[4]\, FCO => 
        \APB3_RDATA_1_25_0_0_co0[4]\);
    
    \APB3_RDATA_1_d_am[5]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => N_1667, B => N_757, C => N_1675, Y => 
        \APB3_RDATA_1_d_am[5]_net_1\);
    
    \APB3_RDATA_1_0_m2_2_wmux_0[0]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_0_m2_2_2_y0[0]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_1_reg[0]_net_1\, D => 
        \mac_3_byte_3_reg[0]_net_1\, FCI => 
        \APB3_RDATA_1_0_m2_2_2_co0[0]\, S => OPEN, Y => 
        \APB3_RDATA_1_0_m2_2_wmux_0_Y[0]\, FCO => OPEN);
    
    \WRITE_REGISTER_ENABLE_PROC.un17_apb3_addr_0_a2\ : CFG3
      generic map(INIT => x"80")

      port map(A => N_802, B => N_791, C => N_789, Y => N_336);
    
    \APB3_RDATA_1_23_0_m2[1]\ : CFG4
      generic map(INIT => x"AA30")

      port map(A => \mac_4_byte_2_reg[1]_net_1\, B => 
        \i_int_mask_reg[1]_net_1\, C => rx_CRC_error_int, D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => N_185);
    
    \mac_1_byte_1_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_1_reg[2]_net_1\);
    
    \APB3_RDATA_1_23_0[2]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => N_186, B => APB3_RDATA_1_sn_m12_i_0, C => 
        \N_817_i\, Y => N_1656);
    
    control_reg_13_0_0_a2_0_0 : CFG4
      generic map(INIT => x"0C88")

      port map(A => TX_PreAmble, B => \control_reg_en\, C => 
        \write_scratch_reg_en\, D => N_581, Y => control_reg_13);
    
    \mac_4_byte_2_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_2_reg[0]_net_1\);
    
    \APB3_RDATA_1_1[3]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \mac_3_byte_6_reg[3]_net_1\, B => 
        \mac_3_byte_2_reg[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_49);
    
    \mac_1_byte_4_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type2_reg[1]\);
    
    \WRITE_REGISTER_ENABLE_PROC.un21_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"2000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_789, D => N_802, Y
         => N_337);
    
    \mac_3_byte_2_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_2_reg[5]_net_1\);
    
    \APB3_RDATA_1_29_d_ns[3]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \APB3_RDATA_1_29_d_bm[3]_net_1\, B => N_78, C
         => \APB3_RDATA_1_29_d_am[3]_net_1\, Y => 
        \APB3_RDATA_1_29_d_ns[3]_net_1\);
    
    \mac_1_byte_4_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type2_reg[0]\);
    
    \APB3_RDATA_1_23_0_m2[2]\ : CFG4
      generic map(INIT => x"AA30")

      port map(A => \mac_4_byte_2_reg[2]_net_1\, B => 
        \i_int_mask_reg[2]_net_1\, C => rx_FIFO_OVERFLOW_int, D
         => CoreAPB3_0_APBmslave0_PADDR(3), Y => N_186);
    
    \APB3_RDATA_1_18_i_m2_0_0_wmux[1]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_3_reg[1]_net_1\, D => 
        \mac_4_byte_4_reg[1]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_18_i_m2_0_0_y0[1]\, FCO => 
        \APB3_RDATA_1_18_i_m2_0_0_co0[1]\);
    
    \RX_packet_depth[6]\ : SLE
      port map(D => \RX_packet_depth_s[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_127_i, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RX_packet_depth[6]_net_1\);
    
    mac_2_byte_1_reg_en_ret_3 : SLE
      port map(D => un12_mac_2_byte_1_reg_en_16_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        N_855_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        un12_mac_2_byte_1_reg_en_16_1_reto);
    
    \mac_3_byte_1_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_1_reg[6]_net_1\);
    
    \N_855_i\ : CFG4
      generic map(INIT => x"0080")

      port map(A => CoreAPB3_0_APBmslave0_PWRITE, B => 
        CoreAPB3_0_APBmslave0_PSELx, C => 
        CoreAPB3_0_APBmslave0_PENABLE, D => long_reset, Y => 
        N_855_i);
    
    \mac_4_byte_3_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_3_reg[0]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \mac_1_byte_4_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type2_reg[5]\);
    
    APB3_RDATA_1_23_2 : CFG3
      generic map(INIT => x"B0")

      port map(A => \N_817_i\, B => \read_reg_en\, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => \APB3_RDATA_1_23_2\);
    
    \APB3_RDATA_1_0_a2_1_0[0]\ : CFG4
      generic map(INIT => x"C080")

      port map(A => \N_817_i\, B => N_742_0, C => 
        CoreAPB3_0_APBmslave0_PADDR(2), D => 
        APB3_RDATA_1_sn_m21_i_1, Y => \APB3_RDATA_1_0_a2_1[0]\);
    
    \RX_packet_depth[2]\ : SLE
      port map(D => \RX_packet_depth_s[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_127_i, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RX_packet_depth[2]_net_1\);
    
    mac_2_byte_1_reg_en_ret_2 : SLE
      port map(D => un12_mac_2_byte_1_reg_en_16_0, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        N_855_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        un12_mac_2_byte_1_reg_en_16_0_reto);
    
    \APB3_RDATA_1_17_0_wmux_0[5]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_17_0_0_y0[5]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_1_byte_1_reg[5]_net_1\, D => 
        \mac_3_byte_5_reg[5]_net_1\, FCI => 
        \APB3_RDATA_1_17_0_0_co0[5]\, S => OPEN, Y => N_1610, FCO
         => OPEN);
    
    mac_2_byte_3_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_343, ALn => N_855_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_2_byte_3_reg_en\);
    
    \iAPB3_READY[0]\ : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => un5_apb3_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \iAPB3_READYrs[0]\);
    
    \APB3_RDATA_1_18_i_m2_0_0_wmux[0]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_3_reg[0]_net_1\, D => 
        \mac_4_byte_4_reg[0]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_18_i_m2_0_0_y0[0]\, FCO => 
        \APB3_RDATA_1_18_i_m2_0_0_co0[0]\);
    
    \mac_1_byte_6_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type3_reg[3]\);
    
    mac_1_byte_2_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_336, ALn => N_855_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_1_byte_2_reg_en\);
    
    \REG_WRITE_PROC.un13_mac_1_byte_5_reg_en_0_a2_1_a2_1_a2\ : 
        CFG4
      generic map(INIT => x"0200")

      port map(A => \mac_1_byte_5_reg_en\, B => 
        \mac_1_byte_4_reg_en\, C => \mac_1_byte_3_reg_en\, D => 
        N_1461, Y => un13_mac_1_byte_5_reg_en);
    
    \RX_packet_depth_cry[4]\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \RX_packet_depth[4]_net_1\, B => 
        rx_packet_complt, C => GND_net_1, D => GND_net_1, FCI => 
        \RX_packet_depth_cry[3]_net_1\, S => 
        \RX_packet_depth_s[4]\, Y => OPEN, FCO => 
        \RX_packet_depth_cry[4]_net_1\);
    
    \mac_3_byte_6_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_6_reg[4]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un25_apb3_addr_0_a2_0\ : CFG2
      generic map(INIT => x"2")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), Y => N_802);
    
    \APB3_RDATA_1_1[1]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \mac_3_byte_6_reg[1]_net_1\, B => 
        \mac_3_byte_2_reg[1]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_1086);
    
    \mac_2_byte_5_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_5_reg[0]_net_1\);
    
    \control_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => control_reg_13, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \control_reg[3]_net_1\);
    
    \APB3_RDATA_1_d_ns[6]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \APB3_RDATA_1_d_bm[6]_net_1\, B => 
        \APB3_RDATA_1_d_am[6]_net_1\, C => N_91, Y => 
        \APB3_RDATA_1_d_ns[6]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_4_byte_4_reg_en_0_a2_0_a2_0_a2\ : 
        CFG4
      generic map(INIT => x"1000")

      port map(A => \mac_1_byte_2_reg_en\, B => 
        \mac_1_byte_1_reg_en\, C => 
        un13_mac_4_byte_4_reg_en_0_a2_0_a2_0_a2_1, D => N_1337, Y
         => un13_mac_4_byte_4_reg_en);
    
    \control_reg_RNO[5]\ : CFG4
      generic map(INIT => x"0CAA")

      port map(A => TX_PreAmble, B => \control_reg_en\, C => 
        \write_scratch_reg_en\, D => N_581, Y => 
        un1_control_reg_en_2_i_0);
    
    \WRITE_REGISTER_ENABLE_PROC.un69_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"2000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_793, D => N_796, Y
         => N_349);
    
    \mac_4_byte_5_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_5_reg[3]_net_1\);
    
    \i_int_mask_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_1354_i, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \i_int_mask_reg[1]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_2_byte_5_reg_en_0_a2_1_a2_0_a2\ : 
        CFG3
      generic map(INIT => x"08")

      port map(A => N_989, B => \mac_2_byte_5_reg_en\, C => N_547, 
        Y => un13_mac_2_byte_5_reg_en);
    
    \APB3_RDATA_1_28[3]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => N_1665, B => N_757, C => N_1673, Y => N_1700);
    
    \REG_WRITE_PROC.un13_mac_4_byte_5_reg_en_0_a2_0_a2_0_a2\ : 
        CFG4
      generic map(INIT => x"0008")

      port map(A => un13_mac_4_byte_5_reg_en_0_a2_0_a2_0_a2_0, B
         => N_1337, C => \mac_1_byte_2_reg_en\, D => N_576, Y => 
        un13_mac_4_byte_5_reg_en);
    
    \APB3_RDATA_1_0_o2[0]\ : CFG4
      generic map(INIT => x"B1A0")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => N_586, D => N_582, Y
         => N_742_0);
    
    \APB3_RDATA_1_21_0_wmux_0[6]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_21_0_0_y0[6]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \consumer_type1_reg[6]\, D => \consumer_type2_reg[6]\, 
        FCI => \APB3_RDATA_1_21_0_0_co0[6]\, S => OPEN, Y => 
        N_1643, FCO => OPEN);
    
    \APB3_RDATA_1_28[1]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => N_1671, B => N_498, C => N_757, Y => N_1698);
    
    \APB3_RDATA_1_26_i_m3_0_wmux_0[1]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_26_i_m3_0_2_y0[1]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \consumer_type1_reg[1]\, D => \consumer_type2_reg[1]\, 
        FCI => \APB3_RDATA_1_26_i_m3_0_2_co0[1]\, S => OPEN, Y
         => N_495, FCO => OPEN);
    
    \WRITE_REGISTER_ENABLE_PROC.un65_apb3_addr_0_a2\ : CFG3
      generic map(INIT => x"80")

      port map(A => N_793, B => N_796, C => N_791, Y => N_348);
    
    \mac_4_byte_5_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_5_reg[6]_net_1\);
    
    \APB3_RDATA_1_24_i_m3_0_2_wmux[1]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \i_int_mask_reg[1]_net_1\, D => \consumer_type2_reg[9]\, 
        FCI => VCC_net_1, S => OPEN, Y => 
        \APB3_RDATA_1_24_i_m3_0_2_y0[1]\, FCO => 
        \APB3_RDATA_1_24_i_m3_0_2_co0[1]\);
    
    \APB3_RDATA_1_17_0_wmux_0[4]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_17_0_0_y0[4]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_1_byte_1_reg[4]_net_1\, D => 
        \mac_3_byte_5_reg[4]_net_1\, FCI => 
        \APB3_RDATA_1_17_0_0_co0[4]\, S => OPEN, Y => N_1609, FCO
         => OPEN);
    
    \APB3_RDATA_1_26_i_m3[1]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => N_495, C
         => N_198, Y => N_499);
    
    \APB3_RDATA_1_17_i_m2_0_0_wmux[2]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \control_reg[2]_net_1\, D => \mac_2_byte_3_reg[2]_net_1\, 
        FCI => VCC_net_1, S => OPEN, Y => 
        \APB3_RDATA_1_17_i_m2_0_0_y0[2]\, FCO => 
        \APB3_RDATA_1_17_i_m2_0_0_co0[2]\);
    
    \APB3_RDATA[3]\ : SLE
      port map(D => \APB3_RDATA_1[3]\, CLK => N_41_mux, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        \CoreAPB3_0_APBmslave0_PRDATA[3]\);
    
    \mac_3_byte_6_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_6_reg[2]_net_1\);
    
    \APB3_RDATA_1_17_0_wmux_0[6]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_17_0_0_y0[6]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_1_byte_1_reg[6]_net_1\, D => 
        \mac_3_byte_5_reg[6]_net_1\, FCI => 
        \APB3_RDATA_1_17_0_0_co0[6]\, S => OPEN, Y => N_1611, FCO
         => OPEN);
    
    \mac_1_byte_1_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_1_reg[7]_net_1\);
    
    \REG_WRITE_PROC.un12_mac_2_byte_1_reg_en_16\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => un12_mac_2_byte_1_reg_en_16_2_reto, B => 
        un12_mac_2_byte_1_reg_en_16_1_reto, C => 
        un12_mac_2_byte_1_reg_en_16_0_reto, D => N_732, Y => 
        N_726);
    
    mac_3_byte_1_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_347, ALn => N_855_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_3_byte_1_reg_en\);
    
    \APB3_RDATA_RNIKMI5[7]\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        \CoreAPB3_0_APBmslave0_PRDATA[7]\, Y => 
        CoreAPB3_0_APBmslave0_PRDATA_m(7));
    
    \APB3_RDATA_1_d_ns[5]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \APB3_RDATA_1_d_bm[5]_net_1\, B => 
        \APB3_RDATA_1_d_am[5]_net_1\, C => N_91, Y => 
        \APB3_RDATA_1_d_ns[5]_net_1\);
    
    mac_1_byte_5_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_339, ALn => N_855_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_1_byte_5_reg_en\);
    
    \APB3_RDATA_1_24[2]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_1623, B => N_1342, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => N_1664);
    
    \APB3_RDATA[6]\ : SLE
      port map(D => \APB3_RDATA_1[6]_net_1\, CLK => N_41_mux, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        \CoreAPB3_0_APBmslave0_PRDATA[6]\);
    
    \REG_WRITE_PROC.un13_mac_1_byte_1_reg_en_0_a2_2_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"8")

      port map(A => N_1455, B => \mac_1_byte_1_reg_en\, Y => 
        un13_mac_1_byte_1_reg_en);
    
    \APB3_RDATA_1_23_1[3]\ : CFG4
      generic map(INIT => x"0C0A")

      port map(A => N_381, B => \mac_4_byte_2_reg[3]_net_1\, C
         => APB3_RDATA_1_sn_m12_i_0, D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => 
        \APB3_RDATA_1_23_1[3]_net_1\);
    
    \mac_1_byte_2_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type1_reg[0]\);
    
    \mac_2_byte_5_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_5_reg[7]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_2_byte_2_reg_en_0_a2_0_a2_0_a2\ : 
        CFG2
      generic map(INIT => x"8")

      port map(A => N_989, B => \mac_2_byte_2_reg_en\, Y => 
        un13_mac_2_byte_2_reg_en);
    
    \APB3_RDATA_1_21_0_0_wmux[3]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_2_byte_4_reg[3]_net_1\, D => 
        \mac_2_byte_6_reg[3]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_21_0_0_y0[3]\, FCO => 
        \APB3_RDATA_1_21_0_0_co0[3]\);
    
    \APB3_RDATA_1_17_0_0_wmux[5]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => \start_tx_FIFO\, D
         => \mac_2_byte_3_reg[5]_net_1\, FCI => VCC_net_1, S => 
        OPEN, Y => \APB3_RDATA_1_17_0_0_y0[5]\, FCO => 
        \APB3_RDATA_1_17_0_0_co0[5]\);
    
    \scratch_pad_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \write_scratch_reg_en\, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \scratch_pad_reg[1]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un73_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_793, D => N_796, Y
         => N_350);
    
    \RX_packet_depth_s[7]\ : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \RX_packet_depth[7]_net_1\, C
         => rx_packet_complt, D => GND_net_1, FCI => 
        \RX_packet_depth_cry[6]_net_1\, S => 
        \RX_packet_depth_s[7]_net_1\, Y => OPEN, FCO => OPEN);
    
    \control_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => control_reg_13, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \TX_FIFO_RST\);
    
    \APB3_RDATA_1_24_i_m3_0_wmux_0[1]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_24_i_m3_0_2_y0[1]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \mac_2_byte_5_reg[1]_net_1\, D => 
        \mac_4_byte_1_reg[1]_net_1\, FCI => 
        \APB3_RDATA_1_24_i_m3_0_2_co0[1]\, S => OPEN, Y => N_496, 
        FCO => OPEN);
    
    \WRITE_REGISTER_ENABLE_PROC.un89_apb3_addr_0_a2_0_a2_0\ : 
        CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), Y => N_796);
    
    \mac_2_byte_5_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_5_reg[4]_net_1\);
    
    \APB3_RDATA_1_1[2]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \mac_3_byte_6_reg[2]_net_1\, B => 
        \mac_3_byte_2_reg[2]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_48);
    
    \mac_3_byte_2_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_2_reg[6]_net_1\);
    
    \mac_3_byte_2_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_2_reg[1]_net_1\);
    
    \APB3_RDATA_1_14_4_wmux_1[1]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => ReadFIFO_Read_Ptr(0), B => 
        ReadFIFO_Read_Ptr(1), C => iRX_FIFO_Full(0), D => 
        iRX_FIFO_Full(1), FCI => \APB3_RDATA_1_14_4_0_co1[1]\, S
         => OPEN, Y => \APB3_RDATA_1_14_4_y0_0[1]\, FCO => 
        \APB3_RDATA_1_14_4_co0_0[1]\);
    
    \mac_1_byte_3_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type2_reg[8]\);
    
    \APB3_RDATA_1_1[4]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \mac_3_byte_6_reg[4]_net_1\, B => 
        \mac_3_byte_2_reg[4]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_50);
    
    \APB3_RDATA_1_28_RNO[2]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \APB3_RDATA_1_25_0_wmux_0_Y[2]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \APB3_RDATA_1_25_3[2]_net_1\, Y => N_1672);
    
    \mac_3_byte_1_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_1_reg[3]_net_1\);
    
    mac_4_byte_3_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_355, ALn => N_855_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_4_byte_3_reg_en\);
    
    \APB3_RDATA_1_21_0_0_wmux[4]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_2_byte_4_reg[4]_net_1\, D => 
        \mac_2_byte_6_reg[4]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_21_0_0_y0[4]\, FCO => 
        \APB3_RDATA_1_21_0_0_co0[4]\);
    
    \APB3_RDATA_1_25_3[6]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_52, B => CoreAPB3_0_APBmslave0_PADDR(3), C
         => N_1495, Y => \APB3_RDATA_1_25_3[6]_net_1\);
    
    \APB3_RDATA_1_24[4]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_1609, B => CoreAPB3_0_APBmslave0_PADDR(3), 
        C => N_1625, Y => N_1666);
    
    \APB3_RDATA_1_22_RNO[4]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \APB3_RDATA_1_14_0_wmux_0_Y[4]\, B => 
        \APB3_RDATA_1_14_3[4]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_1585);
    
    \APB3_RDATA_1_0_m2_1_0[0]\ : CFG3
      generic map(INIT => x"27")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => N_593, C
         => N_197, Y => \APB3_RDATA_1_0_m2_1_0[0]_net_1\);
    
    \mac_4_byte_2_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_2_reg[7]_net_1\);
    
    \APB3_RDATA_1_3[2]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \consumer_type4_reg[2]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_4_reg[2]_net_1\, Y => N_1491);
    
    \mac_2_byte_6_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_6_reg[6]_net_1\);
    
    \APB3_RDATA_1_0_m2_5[0]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \consumer_type3_reg[0]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \scratch_pad_reg[0]_net_1\, Y => N_582);
    
    \WRITE_REGISTER_ENABLE_PROC.un93_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"0200")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(7), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => N_801, Y => N_355);
    
    int_mask_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_333, ALn => N_855_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \int_mask_reg_en\);
    
    \READY_DELAY_PROC.un5_apb3_rst_rs\ : SLE
      port map(D => VCC_net_1, CLK => long_reset, EN => VCC_net_1, 
        ALn => un5_apb3_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => VCC_net_1, Q => un5_apb3_rst_rs);
    
    \REG_WRITE_PROC.un13_mac_4_byte_6_reg_en_0_a2_4_a2_3_a2\ : 
        CFG4
      generic map(INIT => x"0040")

      port map(A => N_731, B => N_1337, C => 
        \mac_4_byte_6_reg_en\, D => N_577, Y => 
        un13_mac_4_byte_6_reg_en);
    
    \APB3_RDATA_1_d_ns[3]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_1657, B => N_1700, C => N_91, Y => 
        \APB3_RDATA_1_d_ns[3]_net_1\);
    
    \scratch_pad_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \write_scratch_reg_en\, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \scratch_pad_reg[0]_net_1\);
    
    \mac_1_byte_5_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_5_reg[3]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_4_byte_2_reg_en_0_a2_3_a2_2_a2\ : 
        CFG3
      generic map(INIT => x"08")

      port map(A => \mac_4_byte_2_reg_en\, B => N_989, C => N_570, 
        Y => un13_mac_4_byte_2_reg_en);
    
    \mac_3_byte_6_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_6_reg[5]_net_1\);
    
    \mac_2_byte_4_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_4_reg[2]_net_1\);
    
    \control_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => control_reg_13, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \control_reg[0]_net_1\);
    
    \APB3_RDATA_1_23[3]\ : CFG4
      generic map(INIT => x"FFF4")

      port map(A => \N_817_i\, B => \APB3_RDATA_1_23_1[3]_net_1\, 
        C => \APB3_RDATA_1_23_1\, D => \APB3_RDATA_1_23_2\, Y => 
        N_1657);
    
    \APB3_RDATA_1_25_0_0_wmux[2]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_1_byte_5_reg[2]_net_1\, D => 
        \mac_2_byte_1_reg[2]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_25_0_0_y0[2]\, FCO => 
        \APB3_RDATA_1_25_0_0_co0[2]\);
    
    \mac_4_byte_3_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_3_reg[7]_net_1\);
    
    \APB3_RDATA_1_1[5]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \mac_3_byte_6_reg[5]_net_1\, B => 
        \mac_3_byte_2_reg[5]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_51);
    
    iTX_FIFO_wr_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un1_apb3_addr, ALn => 
        N_855_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => TX_FIFO_wr_en);
    
    m30_0_a2 : CFG4
      generic map(INIT => x"0004")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(7), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        CoreAPB3_0_APBmslave0_PADDR(1), D => 
        CoreAPB3_0_APBmslave0_PADDR(0), Y => N_234);
    
    \control_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => control_reg_13, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \external_loopback\);
    
    \RX_packet_depth_cry[3]\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \RX_packet_depth[3]_net_1\, B => 
        rx_packet_complt, C => GND_net_1, D => GND_net_1, FCI => 
        \RX_packet_depth_cry[2]_net_1\, S => 
        \RX_packet_depth_s[3]\, Y => OPEN, FCO => 
        \RX_packet_depth_cry[3]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_4_byte_1_reg_en_0_a2_0_a2_0_a2_0\ : 
        CFG4
      generic map(INIT => x"1000")

      port map(A => \mac_1_byte_6_reg_en\, B => 
        \mac_2_byte_1_reg_en\, C => N_1461, D => N_1457, Y => 
        N_989);
    
    \mac_4_byte_3_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_3_reg[1]_net_1\);
    
    \APB3_RDATA_1[6]\ : CFG4
      generic map(INIT => x"F780")

      port map(A => N_78, B => N_91, C => N_1693, D => 
        \APB3_RDATA_1_d_ns[6]_net_1\, Y => 
        \APB3_RDATA_1[6]_net_1\);
    
    \control_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => control_reg_13, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \control_reg[2]_net_1\);
    
    \mac_2_byte_3_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_3_reg[5]_net_1\);
    
    \mac_3_byte_4_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_4_reg[4]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un29_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"1000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_793, D => N_795, Y
         => N_339);
    
    \mac_1_byte_5_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_5_reg[6]_net_1\);
    
    \mac_3_byte_6_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_6_reg[0]_net_1\);
    
    \APB3_RDATA_RNIHJI5[4]\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        \CoreAPB3_0_APBmslave0_PRDATA[4]\, Y => 
        CoreAPB3_0_APBmslave0_PRDATA_m(4));
    
    \APB3_RDATA_1_27[5]\ : CFG3
      generic map(INIT => x"BA")

      port map(A => \APB3_RDATA_1_27_10\, B => \N_817_i\, C => 
        \APB3_RDATA_1_27_1[5]_net_1\, Y => N_1692);
    
    \APB3_RDATA_1_3[4]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \consumer_type4_reg[4]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_4_reg[4]_net_1\, Y => N_1493);
    
    \mac_3_byte_1_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_1_reg[5]_net_1\);
    
    \APB3_RDATA_1_19_0_0_wmux[5]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \i_int_mask_reg[5]_net_1\, D => 
        \mac_1_byte_3_reg[5]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_19_0_0_y0[5]\, FCO => 
        \APB3_RDATA_1_19_0_0_co0[5]\);
    
    \mac_2_byte_5_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_5_reg[5]_net_1\);
    
    \APB3_RDATA_1_26_i_m2[2]\ : CFG3
      generic map(INIT => x"D8")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => N_202, C
         => N_199, Y => N_203);
    
    \WRITE_REGISTER_ENABLE_PROC.un25_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_789, D => N_802, Y
         => N_338);
    
    mac_4_byte_1_reg_en_RNO_0 : CFG3
      generic map(INIT => x"80")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => 
        CoreAPB3_0_APBmslave0_PADDR(6), Y => \m14_0_a3_1\);
    
    \APB3_RDATA_1_25_0_wmux_0[2]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_25_0_0_y0[2]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_1_reg[2]_net_1\, D => 
        \mac_3_byte_3_reg[2]_net_1\, FCI => 
        \APB3_RDATA_1_25_0_0_co0[2]\, S => OPEN, Y => 
        \APB3_RDATA_1_25_0_wmux_0_Y[2]\, FCO => OPEN);
    
    \READY_DELAY_PROC.un5_apb3_rst_0_a2_0_a2\ : CFG3
      generic map(INIT => x"F8")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        CoreAPB3_0_APBmslave0_PENABLE, C => long_reset, Y => 
        un5_apb3_rst_i);
    
    \APB3_RDATA_1_1[6]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \mac_3_byte_6_reg[6]_net_1\, B => 
        \mac_3_byte_2_reg[6]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_52);
    
    \mac_3_byte_1_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_1_reg[2]_net_1\);
    
    read_reg_en_RNIMEE51 : CFG4
      generic map(INIT => x"FEDC")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        APB3_RDATA_1_sn_m12_i_0, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), D => 
        CoreAPB3_0_APBmslave0_PADDR(5), Y => 
        APB3_RDATA_1_sn_m12_i_0_0);
    
    \APB3_RDATA[2]\ : SLE
      port map(D => \APB3_RDATA_1[2]\, CLK => N_41_mux, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        \CoreAPB3_0_APBmslave0_PRDATA[2]\);
    
    \mac_3_byte_4_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_4_reg[1]_net_1\);
    
    mac_1_byte_1_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_335, ALn => N_855_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_1_byte_1_reg_en\);
    
    \APB3_RDATA_1_24_i_m3[1]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_497, B => CoreAPB3_0_APBmslave0_PADDR(3), C
         => N_496, Y => N_498);
    
    \APB3_RDATA_1_21_i_m2_0_0_wmux[2]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_2_byte_4_reg[2]_net_1\, D => 
        \mac_2_byte_6_reg[2]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_21_i_m2_0_0_y0[2]\, FCO => 
        \APB3_RDATA_1_21_i_m2_0_0_co0[2]\);
    
    \N_993_i\ : CFG3
      generic map(INIT => x"80")

      port map(A => SM_advance_i, B => rx_crc_HighByte_en, C => 
        sampler_clk1x_en, Y => N_993_i);
    
    \mac_3_byte_4_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_4_reg[0]_net_1\);
    
    \APB3_RDATA_1_4[2]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \consumer_type3_reg[2]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \scratch_pad_reg[2]_net_1\, Y => N_1501);
    
    \scratch_pad_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \write_scratch_reg_en\, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \scratch_pad_reg[2]_net_1\);
    
    \APB3_RDATA_1_bm_1[2]\ : CFG4
      generic map(INIT => x"0E04")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => N_1501, 
        C => APB3_RDATA_1_sn_m12_i_0_0, D => N_1583, Y => 
        \APB3_RDATA_1_bm_1[2]_net_1\);
    
    \APB3_RDATA_1_0_m2_8_wmux_0[0]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_0_m2_8_2_y0[0]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \consumer_type1_reg[0]\, D => \consumer_type2_reg[0]\, 
        FCI => \APB3_RDATA_1_0_m2_8_2_co0[0]\, S => OPEN, Y => 
        N_593, FCO => OPEN);
    
    \up_EOP_sync_RNIOGPQ[2]\ : CFG3
      generic map(INIT => x"9C")

      port map(A => \up_EOP_sync[1]_net_1\, B => rx_packet_complt, 
        C => \up_EOP_sync[2]_net_1\, Y => N_127_i);
    
    \RX_packet_depth[3]\ : SLE
      port map(D => \RX_packet_depth_s[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_127_i, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RX_packet_depth[3]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un1_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"4000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => N_790, D => N_793, Y
         => un1_apb3_addr);
    
    \mac_2_byte_1_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type4_reg[9]\);
    
    read_reg_en : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => N_854_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \read_reg_en\);
    
    INTERRUPT_INST : Interrupts
      port map(CoreAPB3_0_APBmslave0_PWDATA(7) => 
        CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), i_int_mask_reg(7) => 
        \i_int_mask_reg[7]_net_1\, i_int_mask_reg(6) => 
        \i_int_mask_reg[6]_net_1\, i_int_mask_reg(5) => 
        \i_int_mask_reg[5]_net_1\, i_int_mask_reg(4) => 
        \i_int_mask_reg[4]_net_1\, i_int_mask_reg(3) => 
        \i_int_mask_reg[3]_net_1\, i_int_mask_reg(2) => 
        \i_int_mask_reg[2]_net_1\, i_int_mask_reg(1) => 
        \i_int_mask_reg[1]_net_1\, N_799 => N_799, N_789 => N_789, 
        N_790 => N_790, N_791 => N_791, write_reg_en => 
        \write_reg_en\, CommsFPGA_top_0_INT => 
        CommsFPGA_top_0_INT, RX_packet_depth_status => 
        \RX_packet_depth_status\, un2_apb3_reset => 
        un2_apb3_reset, N_385 => N_385, N_384 => N_384, N_381 => 
        N_381, TX_FIFO_UNDERRUN => TX_FIFO_UNDERRUN, 
        un15_int_reg_clr => un15_int_reg_clr, 
        tx_FIFO_UNDERRUN_int => tx_FIFO_UNDERRUN_int, 
        TX_FIFO_UNDERRUN_set => TX_FIFO_UNDERRUN_set, 
        TX_FIFO_OVERFLOW => TX_FIFO_OVERFLOW, un19_int_reg_clr
         => un19_int_reg_clr, tx_FIFO_OVERFLOW_int => 
        tx_FIFO_OVERFLOW_int, TX_FIFO_OVERFLOW_set => 
        TX_FIFO_OVERFLOW_set, RX_FIFO_UNDERRUN => 
        RX_FIFO_UNDERRUN, un23_int_reg_clr => un23_int_reg_clr, 
        RX_FIFO_UNDERRUN_set => RX_FIFO_UNDERRUN_set, 
        RX_FIFO_OVERFLOW => RX_FIFO_OVERFLOW, un27_int_reg_clr
         => un27_int_reg_clr, rx_FIFO_OVERFLOW_int => 
        rx_FIFO_OVERFLOW_int, RX_FIFO_OVERFLOW_set => 
        RX_FIFO_OVERFLOW_set, rx_CRC_error => rx_CRC_error, 
        un31_int_reg_clr => un31_int_reg_clr, rx_CRC_error_int
         => rx_CRC_error_int, rx_CRC_error_set => 
        rx_CRC_error_set, iup_EOP => \iup_EOP\, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz, 
        tx_packet_complt => tx_packet_complt, CommsFPGA_CCC_0_GL0
         => CommsFPGA_CCC_0_GL0, BIT_CLK => BIT_CLK, 
        un2_apb3_reset_i => un2_apb3_reset_i, un2_apb3_reset_set
         => un2_apb3_reset_set);
    
    \APB3_RDATA_1_23_0[1]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => N_185, B => APB3_RDATA_1_sn_m12_i_0, C => 
        \N_817_i\, Y => N_1655);
    
    \mac_2_byte_5_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_5_reg[1]_net_1\);
    
    \mac_3_byte_4_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_4_reg[5]_net_1\);
    
    mac_3_byte_3_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_349, ALn => N_855_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_3_byte_3_reg_en\);
    
    \mac_1_byte_2_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type1_reg[7]\);
    
    RX_packet_depth_status : SLE
      port map(D => rx_packet_depth_status2, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \RX_packet_depth_status\);
    
    control_reg_13_0_0_a2_0_0_o2 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \mac_4_byte_6_reg_en\, B => N_577, C => N_726, 
        D => N_570, Y => N_581);
    
    \APB3_RDATA_1_21_i_m2_0_wmux_0[2]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_21_i_m2_0_0_y0[2]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \consumer_type1_reg[2]\, D => \consumer_type2_reg[2]\, 
        FCI => \APB3_RDATA_1_21_i_m2_0_0_co0[2]\, S => OPEN, Y
         => N_202, FCO => OPEN);
    
    \APB3_RDATA_1_1[7]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \mac_3_byte_6_reg[7]_net_1\, B => 
        \mac_3_byte_2_reg[7]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_1087);
    
    \APB3_RDATA_1_19_0_0_wmux[2]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \i_int_mask_reg[2]_net_1\, D => 
        \mac_1_byte_3_reg[2]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_19_0_0_y0[2]\, FCO => 
        \APB3_RDATA_1_19_0_0_co0[2]\);
    
    \mac_3_byte_6_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_6_reg[3]_net_1\);
    
    \APB3_RDATA_1_17_0_0_wmux[7]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => \TX_FIFO_RST\, D => 
        \mac_2_byte_3_reg[7]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_17_0_0_y0[7]\, FCO => 
        \APB3_RDATA_1_17_0_0_co0[7]\);
    
    m30_0_a2_1 : CFG4
      generic map(INIT => x"0002")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(4), B => 
        CoreAPB3_0_APBmslave0_PADDR(7), C => 
        CoreAPB3_0_APBmslave0_PADDR(0), D => 
        CoreAPB3_0_APBmslave0_PADDR(1), Y => N_789);
    
    \REG_WRITE_PROC.un13_mac_2_byte_5_reg_en_0_a2_1_a2_0_o2\ : 
        CFG3
      generic map(INIT => x"FE")

      port map(A => \mac_2_byte_4_reg_en\, B => 
        \mac_2_byte_3_reg_en\, C => \mac_2_byte_2_reg_en\, Y => 
        N_547);
    
    \scratch_pad_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \write_scratch_reg_en\, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \scratch_pad_reg[4]_net_1\);
    
    \APB3_RDATA_1_18_i_m2_0_wmux_0[5]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_18_i_m2_0_0_y0[5]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_5_reg[5]_net_1\, D => 
        \mac_4_byte_6_reg[5]_net_1\, FCI => 
        \APB3_RDATA_1_18_i_m2_0_0_co0[5]\, S => OPEN, Y => N_206, 
        FCO => OPEN);
    
    \APB3_RDATA_1_25_3[2]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_48, B => CoreAPB3_0_APBmslave0_PADDR(3), C
         => N_1491, Y => \APB3_RDATA_1_25_3[2]_net_1\);
    
    \mac_1_byte_3_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_3_reg[7]_net_1\);
    
    \control_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => control_reg_13, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \internal_loopback\);
    
    \APB3_RDATA_1_17_i_m2_0_0_wmux[3]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \control_reg[3]_net_1\, D => \mac_2_byte_3_reg[3]_net_1\, 
        FCI => VCC_net_1, S => OPEN, Y => 
        \APB3_RDATA_1_17_i_m2_0_0_y0[3]\, FCO => 
        \APB3_RDATA_1_17_i_m2_0_0_co0[3]\);
    
    \APB3_RDATA_1_18_i_m2_0_0_wmux[3]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_3_reg[3]_net_1\, D => 
        \mac_4_byte_4_reg[3]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_18_i_m2_0_0_y0[3]\, FCO => 
        \APB3_RDATA_1_18_i_m2_0_0_co0[3]\);
    
    \APB3_RDATA_1_0_m2_2_2_wmux[0]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \consumer_type3_reg[8]\, D => \consumer_type4_reg[8]\, 
        FCI => VCC_net_1, S => OPEN, Y => 
        \APB3_RDATA_1_0_m2_2_2_y0[0]\, FCO => 
        \APB3_RDATA_1_0_m2_2_2_co0[0]\);
    
    \mac_1_byte_3_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type2_reg[9]\);
    
    \REG_WRITE_PROC.un13_mac_3_byte_1_reg_en_0_a2_1_a2_0_a2\ : 
        CFG3
      generic map(INIT => x"08")

      port map(A => N_989, B => \mac_3_byte_1_reg_en\, C => N_549, 
        Y => un13_mac_3_byte_1_reg_en);
    
    \mac_2_byte_4_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_4_reg[7]_net_1\);
    
    \mac_2_byte_4_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_4_reg[6]_net_1\);
    
    mac_2_byte_1_reg_en_ret_6 : SLE
      port map(D => N_733, CLK => m2s010_som_sb_0_CCC_71MHz, EN
         => VCC_net_1, ALn => N_855_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        N_733_reto);
    
    \APB3_RDATA_1_am[2]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_1699, B => N_91, C => N_203, Y => 
        \APB3_RDATA_1_am[2]_net_1\);
    
    \mac_2_byte_3_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_3_reg[6]_net_1\);
    
    mac_2_byte_6_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_346, ALn => N_855_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_2_byte_6_reg_en\);
    
    \up_EOP_sync[0]\ : SLE
      port map(D => \iup_EOP\, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => long_reset_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \up_EOP_sync[0]_net_1\);
    
    \APB3_RDATA_1_17_0_0_wmux[4]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => \internal_loopback\, 
        D => \mac_2_byte_3_reg[4]_net_1\, FCI => VCC_net_1, S => 
        OPEN, Y => \APB3_RDATA_1_17_0_0_y0[4]\, FCO => 
        \APB3_RDATA_1_17_0_0_co0[4]\);
    
    \mac_4_byte_5_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_5_reg[0]_net_1\);
    
    \APB3_RDATA_1_29_d_bm[7]\ : CFG4
      generic map(INIT => x"2075")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => RX_FIFO_DOUT(7), D
         => \APB3_RDATA_1_29_d_bm_1_0[7]_net_1\, Y => 
        \APB3_RDATA_1_29_d_bm[7]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un77_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"1000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_789, D => N_796, Y
         => N_351);
    
    \APB3_RDATA_1_18_i_m2_0_wmux_0[2]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_18_i_m2_0_0_y0[2]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_5_reg[2]_net_1\, D => 
        \mac_4_byte_6_reg[2]_net_1\, FCI => 
        \APB3_RDATA_1_18_i_m2_0_0_co0[2]\, S => OPEN, Y => N_199, 
        FCO => OPEN);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CommsFPGA_top is

    port( CoreAPB3_0_APBmslave0_PWDATA       : in    std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PRDATA_m     : out   std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PADDR        : in    std_logic_vector(7 downto 0);
          DEBOUNCE_IN_c                      : in    std_logic_vector(2 downto 0);
          Y_net_0                            : in    std_logic_vector(3 downto 1);
          DEBOUNCE_OUT_net_0_0               : out   std_logic;
          MANCHESTER_IN_c                    : in    std_logic;
          MANCH_OUT_P_c                      : out   std_logic;
          MANCH_OUT_P_c_i                    : out   std_logic;
          DRVR_EN_c                          : out   std_logic;
          N_855_i_i                          : in    std_logic;
          CoreAPB3_0_APBmslave0_PSELx        : in    std_logic;
          CoreAPB3_0_APBmslave0_PENABLE      : in    std_logic;
          CoreAPB3_0_APBmslave0_PREADY_i_m_i : out   std_logic;
          CoreAPB3_0_APBmslave0_PWRITE       : in    std_logic;
          N_855_i                            : out   std_logic;
          CommsFPGA_top_0_INT                : out   std_logic;
          DEBOUNCE_OUT_1_c                   : out   std_logic;
          DEBOUNCE_OUT_2_c                   : out   std_logic;
          CommsFPGA_top_0_CAMERA_NODE        : out   std_logic;
          m2s010_som_sb_0_POWER_ON_RESET_N   : in    std_logic;
          m2s010_som_sb_0_GPIO_28_SW_RESET   : in    std_logic;
          CommsFPGA_CCC_0_LOCK               : in    std_logic;
          CommsFPGA_CCC_0_GL1                : in    std_logic;
          CommsFPGA_CCC_0_GL0                : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz          : in    std_logic
        );

end CommsFPGA_top;

architecture DEF_ARCH of CommsFPGA_top is 

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component TriDebounce
    port( DEBOUNCE_IN_c        : in    std_logic_vector(2 downto 0) := (others => 'U');
          DEBOUNCE_OUT_net_0_0 : out   std_logic;
          DEBOUNCE_OUT_2_c     : out   std_logic;
          DEBOUNCE_OUT_1_c     : out   std_logic;
          BIT_CLK              : in    std_logic := 'U';
          un2_apb3_reset_set   : in    std_logic := 'U';
          un2_apb3_reset       : in    std_logic := 'U'
        );
  end component;

  component ManchesEncoder
    port( manches_in_dly                  : in    std_logic_vector(1 downto 0) := (others => 'U');
          start_tx_FIFO                   : in    std_logic := 'U';
          un1_tx_packet_length_0_sqmuxa_o : out   std_logic;
          TX_DataEn_1_o                   : out   std_logic;
          TX_FIFO_Empty                   : in    std_logic := 'U';
          idle_line5                      : out   std_logic;
          tx_col_detect_en                : out   std_logic;
          CommsFPGA_CCC_0_GL0             : in    std_logic := 'U';
          DRVR_EN_c                       : out   std_logic;
          internal_loopback               : in    std_logic := 'U';
          external_loopback               : in    std_logic := 'U';
          tx_packet_complt                : out   std_logic;
          un2_apb3_reset                  : in    std_logic := 'U';
          N_706                           : in    std_logic := 'U';
          N_704                           : in    std_logic := 'U';
          N_709                           : in    std_logic := 'U';
          N_708                           : in    std_logic := 'U';
          N_707                           : in    std_logic := 'U';
          N_710                           : in    std_logic := 'U';
          N_711                           : in    std_logic := 'U';
          N_705                           : in    std_logic := 'U';
          TX_PreAmble                     : out   std_logic;
          CommsFPGA_CCC_0_GL1             : in    std_logic := 'U';
          byte_clk_en                     : in    std_logic := 'U';
          BIT_CLK                         : in    std_logic := 'U';
          un2_apb3_reset_i                : in    std_logic := 'U';
          MANCH_OUT_P_c_i                 : out   std_logic;
          MANCH_OUT_P_c                   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component ManchesDecoder
    port( RX_FIFO_DIN_pipe    : out   std_logic_vector(8 downto 0);
          rx_crc_data_calc    : out   std_logic_vector(11 downto 10);
          consumer_type1_reg  : in    std_logic_vector(9 downto 0) := (others => 'U');
          consumer_type3_reg  : in    std_logic_vector(9 downto 0) := (others => 'U');
          consumer_type4_reg  : in    std_logic_vector(9 downto 0) := (others => 'U');
          consumer_type2_reg  : in    std_logic_vector(9 downto 0) := (others => 'U');
          manches_in_dly      : out   std_logic_vector(1 downto 0);
          RX_FIFO_DIN         : out   std_logic_vector(3 downto 2);
          lfsr_c_i_i_0        : in    std_logic := 'U';
          rx_CRC_error        : out   std_logic;
          rx_CRC_error_i      : out   std_logic;
          N_993_i             : in    std_logic := 'U';
          N_41_i              : in    std_logic := 'U';
          iRX_FIFO_wr_en      : out   std_logic;
          rx_crc_HighByte_en  : out   std_logic;
          SM_advance_i        : out   std_logic;
          N_535               : out   std_logic;
          rx_packet_complt    : out   std_logic;
          RX_InProcess_d1     : out   std_logic;
          tx_col_detect_en    : in    std_logic := 'U';
          DRVR_EN_c           : in    std_logic := 'U';
          RX_EarlyTerm        : out   std_logic;
          un2_apb3_reset_i    : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          sampler_clk1x_en    : out   std_logic;
          MANCH_OUT_P_c       : in    std_logic := 'U';
          MANCHESTER_IN_c     : in    std_logic := 'U';
          internal_loopback   : in    std_logic := 'U';
          un2_apb3_reset      : in    std_logic := 'U';
          idle_line5          : in    std_logic := 'U'
        );
  end component;

  component FIFOs
    port( iRX_FIFO_Full                   : out   std_logic_vector(3 downto 0);
          RX_FIFO_DIN_pipe                : in    std_logic_vector(8 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PWDATA    : in    std_logic_vector(7 downto 0) := (others => 'U');
          up_EOP_sync                     : in    std_logic_vector(2 downto 1) := (others => 'U');
          RX_FIFO_DOUT                    : out   std_logic_vector(7 downto 5);
          ReadFIFO_Read_Ptr               : out   std_logic_vector(1 downto 0);
          RX_FIFO_DOUT_3_0                : out   std_logic;
          RX_FIFO_DOUT_2_0                : out   std_logic;
          RX_FIFO_DOUT_1_0                : out   std_logic;
          RX_FIFO_DOUT_0_0                : out   std_logic;
          N_674                           : out   std_logic;
          N_673                           : out   std_logic;
          N_672                           : out   std_logic;
          N_667                           : out   std_logic;
          N_666                           : out   std_logic;
          N_665                           : out   std_logic;
          N_660                           : out   std_logic;
          N_659                           : out   std_logic;
          N_658                           : out   std_logic;
          iRX_FIFO_wr_en                  : in    std_logic := 'U';
          sampler_clk1x_en                : in    std_logic := 'U';
          RX_InProcess_d1                 : in    std_logic := 'U';
          tx_col_detect_en                : in    std_logic := 'U';
          N_653                           : out   std_logic;
          N_652                           : out   std_logic;
          N_651                           : out   std_logic;
          TX_FIFO_UNDERRUN                : out   std_logic;
          TX_FIFO_UNDERRUN_i              : out   std_logic;
          TX_FIFO_OVERFLOW                : out   std_logic;
          TX_FIFO_OVERFLOW_i              : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz       : in    std_logic := 'U';
          TX_FIFO_Full                    : out   std_logic;
          TX_FIFO_wr_en                   : in    std_logic := 'U';
          un1_tx_packet_length_0_sqmuxa_o : in    std_logic := 'U';
          TX_DataEn_1_o                   : in    std_logic := 'U';
          TX_PreAmble                     : in    std_logic := 'U';
          N_704                           : out   std_logic;
          N_705                           : out   std_logic;
          N_706                           : out   std_logic;
          N_707                           : out   std_logic;
          N_708                           : out   std_logic;
          N_709                           : out   std_logic;
          N_710                           : out   std_logic;
          N_711                           : out   std_logic;
          byte_clk_en                     : in    std_logic := 'U';
          TX_FIFO_Empty                   : out   std_logic;
          BIT_CLK                         : in    std_logic := 'U';
          RX_FIFO_RST                     : in    std_logic := 'U';
          RX_FIFO_rd_en                   : in    std_logic := 'U';
          TX_FIFO_RST                     : in    std_logic := 'U';
          un2_apb3_reset                  : in    std_logic := 'U';
          rx_packet_complt                : in    std_logic := 'U';
          N_678                           : out   std_logic;
          N_712                           : out   std_logic;
          N_693                           : out   std_logic;
          CommsFPGA_CCC_0_GL0             : in    std_logic := 'U';
          RX_FIFO_OVERFLOW_i              : out   std_logic;
          RX_FIFO_OVERFLOW                : out   std_logic;
          RX_FIFO_UNDERRUN_i              : out   std_logic;
          RX_FIFO_UNDERRUN                : out   std_logic
        );
  end component;

  component uP_if
    port( RX_FIFO_DIN                        : in    std_logic_vector(3 downto 2) := (others => 'U');
          rx_crc_data_calc                   : in    std_logic_vector(11 downto 10) := (others => 'U');
          CoreAPB3_0_APBmslave0_PADDR        : in    std_logic_vector(7 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PRDATA_m     : out   std_logic_vector(7 downto 0);
          RX_FIFO_DOUT                       : in    std_logic_vector(7 downto 5) := (others => 'U');
          iRX_FIFO_Full                      : in    std_logic_vector(3 downto 0) := (others => 'U');
          ReadFIFO_Read_Ptr                  : in    std_logic_vector(1 downto 0) := (others => 'U');
          consumer_type4_reg                 : out   std_logic_vector(9 downto 0);
          consumer_type3_reg                 : out   std_logic_vector(9 downto 0);
          consumer_type2_reg                 : out   std_logic_vector(9 downto 0);
          consumer_type1_reg                 : out   std_logic_vector(9 downto 0);
          CoreAPB3_0_APBmslave0_PWDATA       : in    std_logic_vector(7 downto 0) := (others => 'U');
          up_EOP_sync                        : out   std_logic_vector(2 downto 1);
          lfsr_c_i_i_0                       : out   std_logic;
          RX_FIFO_DIN_pipe_0                 : in    std_logic := 'U';
          RX_FIFO_DOUT_1_0                   : in    std_logic := 'U';
          RX_FIFO_DOUT_0_0                   : in    std_logic := 'U';
          RX_FIFO_DOUT_3_0                   : in    std_logic := 'U';
          RX_FIFO_DOUT_2_0                   : in    std_logic := 'U';
          un2_apb3_reset_set                 : out   std_logic;
          un2_apb3_reset_i                   : in    std_logic := 'U';
          BIT_CLK                            : in    std_logic := 'U';
          tx_packet_complt                   : in    std_logic := 'U';
          rx_CRC_error_set                   : in    std_logic := 'U';
          un31_int_reg_clr                   : out   std_logic;
          rx_CRC_error                       : in    std_logic := 'U';
          RX_FIFO_OVERFLOW_set               : in    std_logic := 'U';
          un27_int_reg_clr                   : out   std_logic;
          RX_FIFO_OVERFLOW                   : in    std_logic := 'U';
          RX_FIFO_UNDERRUN_set               : in    std_logic := 'U';
          un23_int_reg_clr                   : out   std_logic;
          RX_FIFO_UNDERRUN                   : in    std_logic := 'U';
          TX_FIFO_OVERFLOW_set               : in    std_logic := 'U';
          un19_int_reg_clr                   : out   std_logic;
          TX_FIFO_OVERFLOW                   : in    std_logic := 'U';
          TX_FIFO_UNDERRUN_set               : in    std_logic := 'U';
          un15_int_reg_clr                   : out   std_logic;
          TX_FIFO_UNDERRUN                   : in    std_logic := 'U';
          un2_apb3_reset                     : in    std_logic := 'U';
          CommsFPGA_top_0_INT                : out   std_logic;
          TX_PreAmble                        : in    std_logic := 'U';
          N_712                              : in    std_logic := 'U';
          N_855_i                            : out   std_logic;
          CoreAPB3_0_APBmslave0_PWRITE       : in    std_logic := 'U';
          N_993_i                            : out   std_logic;
          sampler_clk1x_en                   : in    std_logic := 'U';
          SM_advance_i                       : in    std_logic := 'U';
          N_41_i                             : out   std_logic;
          rx_crc_HighByte_en                 : in    std_logic := 'U';
          N_535                              : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PREADY_i_m_i : out   std_logic;
          CoreAPB3_0_APBmslave0_PENABLE      : in    std_logic := 'U';
          RX_FIFO_RST_1                      : out   std_logic;
          RX_EarlyTerm                       : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PSELx        : in    std_logic := 'U';
          TX_FIFO_Empty                      : in    std_logic := 'U';
          TX_FIFO_Full                       : in    std_logic := 'U';
          N_693                              : in    std_logic := 'U';
          N_678                              : in    std_logic := 'U';
          N_658                              : in    std_logic := 'U';
          N_651                              : in    std_logic := 'U';
          N_672                              : in    std_logic := 'U';
          N_665                              : in    std_logic := 'U';
          N_659                              : in    std_logic := 'U';
          N_652                              : in    std_logic := 'U';
          N_673                              : in    std_logic := 'U';
          N_666                              : in    std_logic := 'U';
          N_660                              : in    std_logic := 'U';
          N_653                              : in    std_logic := 'U';
          N_674                              : in    std_logic := 'U';
          N_667                              : in    std_logic := 'U';
          rx_packet_complt                   : in    std_logic := 'U';
          RX_FIFO_rd_en                      : out   std_logic;
          TX_FIFO_wr_en                      : out   std_logic;
          N_855_i_i                          : in    std_logic := 'U';
          TX_FIFO_RST                        : out   std_logic;
          start_tx_FIFO                      : out   std_logic;
          internal_loopback                  : out   std_logic;
          external_loopback                  : out   std_logic;
          long_reset                         : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz          : in    std_logic := 'U';
          long_reset_set                     : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0                : in    std_logic := 'U';
          long_reset_i                       : in    std_logic := 'U'
        );
  end component;

    signal bd_reset_i, \bd_reset\, \long_reset\, long_reset_0, 
        \BIT_CLK\, BIT_CLK_0, un2_apb3_reset, \RESET\, 
        \ClkDivider[0]_net_1\, \ClkDivider_i[0]\, BIT_CLK_i_i, 
        un2_apb3_reset_i, long_reset_i, \long_reset_set\, 
        GND_net_1, VCC_net_1, \rx_CRC_error_set\, rx_CRC_error_i, 
        un31_int_reg_clr, \RX_FIFO_OVERFLOW_set\, 
        RX_FIFO_OVERFLOW_i, un27_int_reg_clr, 
        \RX_FIFO_UNDERRUN_set\, RX_FIFO_UNDERRUN_i, 
        un23_int_reg_clr, \TX_FIFO_OVERFLOW_set\, 
        TX_FIFO_OVERFLOW_i, un19_int_reg_clr, 
        \TX_FIFO_UNDERRUN_set\, TX_FIFO_UNDERRUN_i, 
        un15_int_reg_clr, \ClkDivider[1]_net_1\, 
        \ClkDivider_RNO[1]_net_1\, \ClkDivider[2]_net_1\, 
        \ClkDivider_RNO[2]_net_1\, \long_reset_cntr[0]_net_1\, 
        \long_reset_cntr_3[0]_net_1\, \long_reset_cntr[1]_net_1\, 
        \long_reset_cntr_3[1]_net_1\, \long_reset_cntr[2]_net_1\, 
        \long_reset_cntr_3[2]_net_1\, \long_reset_cntr[3]_net_1\, 
        \long_reset_cntr_3[3]_net_1\, \long_reset_cntr[4]_net_1\, 
        \long_reset_cntr_3[4]_net_1\, \long_reset_cntr[5]_net_1\, 
        \long_reset_cntr_3[5]_net_1\, \long_reset_cntr[6]_net_1\, 
        un4_long_reset_cntr_cry_6_S, \long_reset_cntr[7]_net_1\, 
        un4_long_reset_cntr_s_7_S, un2_long_reset_cntr_i, 
        \RX_FIFO_RST\, RX_FIFO_RST_1, \byte_clk_en\, 
        byte_clk_en_1, un4_long_reset_cntr_s_1_396_FCO, 
        \un4_long_reset_cntr_cry_1\, un4_long_reset_cntr_cry_1_S, 
        \un4_long_reset_cntr_cry_2\, un4_long_reset_cntr_cry_2_S, 
        \un4_long_reset_cntr_cry_3\, un4_long_reset_cntr_cry_3_S, 
        \un4_long_reset_cntr_cry_4\, un4_long_reset_cntr_cry_4_S, 
        \un4_long_reset_cntr_cry_5\, un4_long_reset_cntr_cry_5_S, 
        \un4_long_reset_cntr_cry_6\, un2_long_reset_cntr_5, 
        un2_long_reset_cntr_4, un2_apb3_reset_set, 
        \lfsr_c_i_i[4]\, \RX_FIFO_DIN[2]\, \RX_FIFO_DIN[3]\, 
        \rx_crc_data_calc[10]\, \rx_crc_data_calc[11]\, 
        \RX_FIFO_DIN_pipe[8]\, \RX_FIFO_DOUT[5]\, 
        \RX_FIFO_DOUT[6]\, \RX_FIFO_DOUT[7]\, \RX_FIFO_DOUT_1[1]\, 
        \RX_FIFO_DOUT_0[1]\, \RX_FIFO_DOUT_3[1]\, 
        \RX_FIFO_DOUT_2[1]\, \iRX_FIFO_Full[0]\, 
        \iRX_FIFO_Full[1]\, \iRX_FIFO_Full[2]\, 
        \iRX_FIFO_Full[3]\, \ReadFIFO_Read_Ptr[0]\, 
        \ReadFIFO_Read_Ptr[1]\, \consumer_type4_reg[0]\, 
        \consumer_type4_reg[1]\, \consumer_type4_reg[2]\, 
        \consumer_type4_reg[3]\, \consumer_type4_reg[4]\, 
        \consumer_type4_reg[5]\, \consumer_type4_reg[6]\, 
        \consumer_type4_reg[7]\, \consumer_type4_reg[8]\, 
        \consumer_type4_reg[9]\, \consumer_type3_reg[0]\, 
        \consumer_type3_reg[1]\, \consumer_type3_reg[2]\, 
        \consumer_type3_reg[3]\, \consumer_type3_reg[4]\, 
        \consumer_type3_reg[5]\, \consumer_type3_reg[6]\, 
        \consumer_type3_reg[7]\, \consumer_type3_reg[8]\, 
        \consumer_type3_reg[9]\, \consumer_type2_reg[0]\, 
        \consumer_type2_reg[1]\, \consumer_type2_reg[2]\, 
        \consumer_type2_reg[3]\, \consumer_type2_reg[4]\, 
        \consumer_type2_reg[5]\, \consumer_type2_reg[6]\, 
        \consumer_type2_reg[7]\, \consumer_type2_reg[8]\, 
        \consumer_type2_reg[9]\, \consumer_type1_reg[0]\, 
        \consumer_type1_reg[1]\, \consumer_type1_reg[2]\, 
        \consumer_type1_reg[3]\, \consumer_type1_reg[4]\, 
        \consumer_type1_reg[5]\, \consumer_type1_reg[6]\, 
        \consumer_type1_reg[7]\, \consumer_type1_reg[8]\, 
        \consumer_type1_reg[9]\, \up_EOP_sync[1]\, 
        \up_EOP_sync[2]\, tx_packet_complt, rx_CRC_error, 
        RX_FIFO_OVERFLOW, RX_FIFO_UNDERRUN, TX_FIFO_OVERFLOW, 
        TX_FIFO_UNDERRUN, TX_PreAmble, N_712, N_993_i, 
        sampler_clk1x_en, SM_advance_i, N_41_i, 
        rx_crc_HighByte_en, N_535, RX_EarlyTerm, TX_FIFO_Empty, 
        TX_FIFO_Full, N_693, N_678, N_658, N_651, N_672, N_665, 
        N_659, N_652, N_673, N_666, N_660, N_653, N_674, N_667, 
        rx_packet_complt, RX_FIFO_rd_en, TX_FIFO_wr_en, 
        TX_FIFO_RST, start_tx_FIFO, internal_loopback, 
        external_loopback, \RX_FIFO_DIN_pipe[0]\, 
        \RX_FIFO_DIN_pipe[1]\, \RX_FIFO_DIN_pipe[2]\, 
        \RX_FIFO_DIN_pipe[3]\, \RX_FIFO_DIN_pipe[4]\, 
        \RX_FIFO_DIN_pipe[5]\, \RX_FIFO_DIN_pipe[6]\, 
        \RX_FIFO_DIN_pipe[7]\, iRX_FIFO_wr_en, RX_InProcess_d1, 
        tx_col_detect_en, un1_tx_packet_length_0_sqmuxa_o, 
        TX_DataEn_1_o, N_704, N_705, N_706, N_707, N_708, N_709, 
        N_710, N_711, \manches_in_dly[0]\, \manches_in_dly[1]\, 
        idle_line5, \DRVR_EN_c\, \MANCH_OUT_P_c\ : std_logic;

    for all : TriDebounce
	Use entity work.TriDebounce(DEF_ARCH);
    for all : ManchesEncoder
	Use entity work.ManchesEncoder(DEF_ARCH);
    for all : ManchesDecoder
	Use entity work.ManchesDecoder(DEF_ARCH);
    for all : FIFOs
	Use entity work.FIFOs(DEF_ARCH);
    for all : uP_if
	Use entity work.uP_if(DEF_ARCH);
begin 

    MANCH_OUT_P_c <= \MANCH_OUT_P_c\;
    DRVR_EN_c <= \DRVR_EN_c\;

    BIT_CLK_inferred_clock_RNIT9E2 : CLKINT
      port map(A => BIT_CLK_0, Y => \BIT_CLK\);
    
    \long_reset_cntr_3[3]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => un2_long_reset_cntr_4, B => 
        un2_long_reset_cntr_5, C => un4_long_reset_cntr_cry_3_S, 
        Y => \long_reset_cntr_3[3]_net_1\);
    
    bd_reset : CFG2
      generic map(INIT => x"4")

      port map(A => m2s010_som_sb_0_GPIO_28_SW_RESET, B => 
        m2s010_som_sb_0_POWER_ON_RESET_N, Y => \bd_reset\);
    
    \long_reset_cntr[3]\ : SLE
      port map(D => \long_reset_cntr_3[3]_net_1\, CLK => 
        \BIT_CLK\, EN => VCC_net_1, ALn => bd_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \long_reset_cntr[3]_net_1\);
    
    \RESET_DELAY_PROC.un2_long_reset_cntr_4\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \long_reset_cntr[4]_net_1\, B => 
        \long_reset_cntr[3]_net_1\, C => 
        \long_reset_cntr[2]_net_1\, D => 
        \long_reset_cntr[1]_net_1\, Y => un2_long_reset_cntr_4);
    
    \long_reset_cntr[6]\ : SLE
      port map(D => un4_long_reset_cntr_cry_6_S, CLK => \BIT_CLK\, 
        EN => VCC_net_1, ALn => bd_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \long_reset_cntr[6]_net_1\);
    
    \ClkDivider_RNO[2]\ : CFG3
      generic map(INIT => x"6A")

      port map(A => \ClkDivider[2]_net_1\, B => 
        \ClkDivider[1]_net_1\, C => \ClkDivider[0]_net_1\, Y => 
        \ClkDivider_RNO[2]_net_1\);
    
    byte_clk_en : SLE
      port map(D => byte_clk_en_1, CLK => \BIT_CLK\, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \byte_clk_en\);
    
    long_reset_set : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => long_reset_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \long_reset_set\);
    
    \ClkDivider_RNO[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \ClkDivider[0]_net_1\, B => 
        \ClkDivider[1]_net_1\, Y => \ClkDivider_RNO[1]_net_1\);
    
    \RESET_DELAY_PROC.un2_long_reset_cntr_5\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \long_reset_cntr[7]_net_1\, B => 
        \long_reset_cntr[6]_net_1\, C => 
        \long_reset_cntr[5]_net_1\, D => 
        \long_reset_cntr[0]_net_1\, Y => un2_long_reset_cntr_5);
    
    un4_long_reset_cntr_cry_2 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \long_reset_cntr[2]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un4_long_reset_cntr_cry_1\, S => 
        un4_long_reset_cntr_cry_2_S, Y => OPEN, FCO => 
        \un4_long_reset_cntr_cry_2\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \ID_RES_DECODE_PROC.un4_id_res\ : CFG3
      generic map(INIT => x"08")

      port map(A => Y_net_0(3), B => Y_net_0(2), C => Y_net_0(1), 
        Y => CommsFPGA_top_0_CAMERA_NODE);
    
    RESET_RNIFEG6 : CLKINT
      port map(A => \RESET\, Y => un2_apb3_reset);
    
    \ClkDivider_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \ClkDivider[0]_net_1\, Y => \ClkDivider_i[0]\);
    
    \long_reset_cntr[5]\ : SLE
      port map(D => \long_reset_cntr_3[5]_net_1\, CLK => 
        \BIT_CLK\, EN => VCC_net_1, ALn => bd_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \long_reset_cntr[5]_net_1\);
    
    TRIPLE_DEBOUNCE_INST : TriDebounce
      port map(DEBOUNCE_IN_c(2) => DEBOUNCE_IN_c(2), 
        DEBOUNCE_IN_c(1) => DEBOUNCE_IN_c(1), DEBOUNCE_IN_c(0)
         => DEBOUNCE_IN_c(0), DEBOUNCE_OUT_net_0_0 => 
        DEBOUNCE_OUT_net_0_0, DEBOUNCE_OUT_2_c => 
        DEBOUNCE_OUT_2_c, DEBOUNCE_OUT_1_c => DEBOUNCE_OUT_1_c, 
        BIT_CLK => \BIT_CLK\, un2_apb3_reset_set => 
        un2_apb3_reset_set, un2_apb3_reset => un2_apb3_reset);
    
    un4_long_reset_cntr_cry_3 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \long_reset_cntr[3]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un4_long_reset_cntr_cry_2\, S => 
        un4_long_reset_cntr_cry_3_S, Y => OPEN, FCO => 
        \un4_long_reset_cntr_cry_3\);
    
    MANCHESTER_ENCODER_INST : ManchesEncoder
      port map(manches_in_dly(1) => \manches_in_dly[1]\, 
        manches_in_dly(0) => \manches_in_dly[0]\, start_tx_FIFO
         => start_tx_FIFO, un1_tx_packet_length_0_sqmuxa_o => 
        un1_tx_packet_length_0_sqmuxa_o, TX_DataEn_1_o => 
        TX_DataEn_1_o, TX_FIFO_Empty => TX_FIFO_Empty, idle_line5
         => idle_line5, tx_col_detect_en => tx_col_detect_en, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, DRVR_EN_c => 
        \DRVR_EN_c\, internal_loopback => internal_loopback, 
        external_loopback => external_loopback, tx_packet_complt
         => tx_packet_complt, un2_apb3_reset => un2_apb3_reset, 
        N_706 => N_706, N_704 => N_704, N_709 => N_709, N_708 => 
        N_708, N_707 => N_707, N_710 => N_710, N_711 => N_711, 
        N_705 => N_705, TX_PreAmble => TX_PreAmble, 
        CommsFPGA_CCC_0_GL1 => CommsFPGA_CCC_0_GL1, byte_clk_en
         => \byte_clk_en\, BIT_CLK => \BIT_CLK\, un2_apb3_reset_i
         => un2_apb3_reset_i, MANCH_OUT_P_c_i => MANCH_OUT_P_c_i, 
        MANCH_OUT_P_c => \MANCH_OUT_P_c\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \SAMPLE_5MHZ_EN_PROC.byte_clk_en_1\ : CFG3
      generic map(INIT => x"08")

      port map(A => \ClkDivider[2]_net_1\, B => 
        \ClkDivider[1]_net_1\, C => \ClkDivider[0]_net_1\, Y => 
        byte_clk_en_1);
    
    \long_reset_cntr[7]\ : SLE
      port map(D => un4_long_reset_cntr_s_7_S, CLK => \BIT_CLK\, 
        EN => VCC_net_1, ALn => bd_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \long_reset_cntr[7]_net_1\);
    
    long_reset : SLE
      port map(D => un2_long_reset_cntr_i, CLK => \BIT_CLK\, EN
         => VCC_net_1, ALn => bd_reset_i, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        long_reset_0);
    
    TX_FIFO_OVERFLOW_set : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => un19_int_reg_clr, ALn => TX_FIFO_OVERFLOW_i, ADn
         => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \TX_FIFO_OVERFLOW_set\);
    
    RX_FIFO_OVERFLOW_set : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => un27_int_reg_clr, ALn => RX_FIFO_OVERFLOW_i, ADn
         => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_OVERFLOW_set\);
    
    un4_long_reset_cntr_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \long_reset_cntr[4]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un4_long_reset_cntr_cry_3\, S => 
        un4_long_reset_cntr_cry_4_S, Y => OPEN, FCO => 
        \un4_long_reset_cntr_cry_4\);
    
    long_reset_RNO : CFG2
      generic map(INIT => x"7")

      port map(A => un2_long_reset_cntr_5, B => 
        un2_long_reset_cntr_4, Y => un2_long_reset_cntr_i);
    
    BIT_CLK : SLE
      port map(D => BIT_CLK_i_i, CLK => CommsFPGA_CCC_0_GL1, EN
         => VCC_net_1, ALn => bd_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        BIT_CLK_0);
    
    MANCHESTER_DECODER_INST : ManchesDecoder
      port map(RX_FIFO_DIN_pipe(8) => \RX_FIFO_DIN_pipe[8]\, 
        RX_FIFO_DIN_pipe(7) => \RX_FIFO_DIN_pipe[7]\, 
        RX_FIFO_DIN_pipe(6) => \RX_FIFO_DIN_pipe[6]\, 
        RX_FIFO_DIN_pipe(5) => \RX_FIFO_DIN_pipe[5]\, 
        RX_FIFO_DIN_pipe(4) => \RX_FIFO_DIN_pipe[4]\, 
        RX_FIFO_DIN_pipe(3) => \RX_FIFO_DIN_pipe[3]\, 
        RX_FIFO_DIN_pipe(2) => \RX_FIFO_DIN_pipe[2]\, 
        RX_FIFO_DIN_pipe(1) => \RX_FIFO_DIN_pipe[1]\, 
        RX_FIFO_DIN_pipe(0) => \RX_FIFO_DIN_pipe[0]\, 
        rx_crc_data_calc(11) => \rx_crc_data_calc[11]\, 
        rx_crc_data_calc(10) => \rx_crc_data_calc[10]\, 
        consumer_type1_reg(9) => \consumer_type1_reg[9]\, 
        consumer_type1_reg(8) => \consumer_type1_reg[8]\, 
        consumer_type1_reg(7) => \consumer_type1_reg[7]\, 
        consumer_type1_reg(6) => \consumer_type1_reg[6]\, 
        consumer_type1_reg(5) => \consumer_type1_reg[5]\, 
        consumer_type1_reg(4) => \consumer_type1_reg[4]\, 
        consumer_type1_reg(3) => \consumer_type1_reg[3]\, 
        consumer_type1_reg(2) => \consumer_type1_reg[2]\, 
        consumer_type1_reg(1) => \consumer_type1_reg[1]\, 
        consumer_type1_reg(0) => \consumer_type1_reg[0]\, 
        consumer_type3_reg(9) => \consumer_type3_reg[9]\, 
        consumer_type3_reg(8) => \consumer_type3_reg[8]\, 
        consumer_type3_reg(7) => \consumer_type3_reg[7]\, 
        consumer_type3_reg(6) => \consumer_type3_reg[6]\, 
        consumer_type3_reg(5) => \consumer_type3_reg[5]\, 
        consumer_type3_reg(4) => \consumer_type3_reg[4]\, 
        consumer_type3_reg(3) => \consumer_type3_reg[3]\, 
        consumer_type3_reg(2) => \consumer_type3_reg[2]\, 
        consumer_type3_reg(1) => \consumer_type3_reg[1]\, 
        consumer_type3_reg(0) => \consumer_type3_reg[0]\, 
        consumer_type4_reg(9) => \consumer_type4_reg[9]\, 
        consumer_type4_reg(8) => \consumer_type4_reg[8]\, 
        consumer_type4_reg(7) => \consumer_type4_reg[7]\, 
        consumer_type4_reg(6) => \consumer_type4_reg[6]\, 
        consumer_type4_reg(5) => \consumer_type4_reg[5]\, 
        consumer_type4_reg(4) => \consumer_type4_reg[4]\, 
        consumer_type4_reg(3) => \consumer_type4_reg[3]\, 
        consumer_type4_reg(2) => \consumer_type4_reg[2]\, 
        consumer_type4_reg(1) => \consumer_type4_reg[1]\, 
        consumer_type4_reg(0) => \consumer_type4_reg[0]\, 
        consumer_type2_reg(9) => \consumer_type2_reg[9]\, 
        consumer_type2_reg(8) => \consumer_type2_reg[8]\, 
        consumer_type2_reg(7) => \consumer_type2_reg[7]\, 
        consumer_type2_reg(6) => \consumer_type2_reg[6]\, 
        consumer_type2_reg(5) => \consumer_type2_reg[5]\, 
        consumer_type2_reg(4) => \consumer_type2_reg[4]\, 
        consumer_type2_reg(3) => \consumer_type2_reg[3]\, 
        consumer_type2_reg(2) => \consumer_type2_reg[2]\, 
        consumer_type2_reg(1) => \consumer_type2_reg[1]\, 
        consumer_type2_reg(0) => \consumer_type2_reg[0]\, 
        manches_in_dly(1) => \manches_in_dly[1]\, 
        manches_in_dly(0) => \manches_in_dly[0]\, RX_FIFO_DIN(3)
         => \RX_FIFO_DIN[3]\, RX_FIFO_DIN(2) => \RX_FIFO_DIN[2]\, 
        lfsr_c_i_i_0 => \lfsr_c_i_i[4]\, rx_CRC_error => 
        rx_CRC_error, rx_CRC_error_i => rx_CRC_error_i, N_993_i
         => N_993_i, N_41_i => N_41_i, iRX_FIFO_wr_en => 
        iRX_FIFO_wr_en, rx_crc_HighByte_en => rx_crc_HighByte_en, 
        SM_advance_i => SM_advance_i, N_535 => N_535, 
        rx_packet_complt => rx_packet_complt, RX_InProcess_d1 => 
        RX_InProcess_d1, tx_col_detect_en => tx_col_detect_en, 
        DRVR_EN_c => \DRVR_EN_c\, RX_EarlyTerm => RX_EarlyTerm, 
        un2_apb3_reset_i => un2_apb3_reset_i, CommsFPGA_CCC_0_GL0
         => CommsFPGA_CCC_0_GL0, sampler_clk1x_en => 
        sampler_clk1x_en, MANCH_OUT_P_c => \MANCH_OUT_P_c\, 
        MANCHESTER_IN_c => MANCHESTER_IN_c, internal_loopback => 
        internal_loopback, un2_apb3_reset => un2_apb3_reset, 
        idle_line5 => idle_line5);
    
    RESET : CFG2
      generic map(INIT => x"D")

      port map(A => CommsFPGA_CCC_0_LOCK, B => \long_reset\, Y
         => \RESET\);
    
    \long_reset_cntr_3[2]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => un2_long_reset_cntr_4, B => 
        un2_long_reset_cntr_5, C => un4_long_reset_cntr_cry_2_S, 
        Y => \long_reset_cntr_3[2]_net_1\);
    
    \long_reset_cntr_3[1]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => un2_long_reset_cntr_4, B => 
        un2_long_reset_cntr_5, C => un4_long_reset_cntr_cry_1_S, 
        Y => \long_reset_cntr_3[1]_net_1\);
    
    un4_long_reset_cntr_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \long_reset_cntr[5]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un4_long_reset_cntr_cry_4\, S => 
        un4_long_reset_cntr_cry_5_S, Y => OPEN, FCO => 
        \un4_long_reset_cntr_cry_5\);
    
    un4_long_reset_cntr_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \long_reset_cntr[6]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un4_long_reset_cntr_cry_5\, S => 
        un4_long_reset_cntr_cry_6_S, Y => OPEN, FCO => 
        \un4_long_reset_cntr_cry_6\);
    
    rx_CRC_error_set : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => un31_int_reg_clr, ALn => rx_CRC_error_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_CRC_error_set\);
    
    BIT_CLK_RNO : CFG1
      generic map(INIT => "01")

      port map(A => BIT_CLK_0, Y => BIT_CLK_i_i);
    
    un4_long_reset_cntr_s_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \long_reset_cntr[7]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un4_long_reset_cntr_cry_6\, S => 
        un4_long_reset_cntr_s_7_S, Y => OPEN, FCO => OPEN);
    
    long_reset_RNIUA27 : CLKINT
      port map(A => long_reset_0, Y => \long_reset\);
    
    \ClkDivider[2]\ : SLE
      port map(D => \ClkDivider_RNO[2]_net_1\, CLK => \BIT_CLK\, 
        EN => VCC_net_1, ALn => bd_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ClkDivider[2]_net_1\);
    
    un4_long_reset_cntr_cry_1 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \long_reset_cntr[1]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        un4_long_reset_cntr_s_1_396_FCO, S => 
        un4_long_reset_cntr_cry_1_S, Y => OPEN, FCO => 
        \un4_long_reset_cntr_cry_1\);
    
    \long_reset_cntr_3[5]\ : CFG3
      generic map(INIT => x"70")

      port map(A => un2_long_reset_cntr_4, B => 
        un2_long_reset_cntr_5, C => un4_long_reset_cntr_cry_5_S, 
        Y => \long_reset_cntr_3[5]_net_1\);
    
    un4_long_reset_cntr_s_1_396 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \long_reset_cntr[0]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => 
        OPEN, Y => OPEN, FCO => un4_long_reset_cntr_s_1_396_FCO);
    
    RX_FIFO_RST : SLE
      port map(D => RX_FIFO_RST_1, CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => bd_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RX_FIFO_RST\);
    
    \ClkDivider[0]\ : SLE
      port map(D => \ClkDivider_i[0]\, CLK => \BIT_CLK\, EN => 
        VCC_net_1, ALn => bd_reset_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ClkDivider[0]_net_1\);
    
    long_reset_RNIUA27_0 : CFG1
      generic map(INIT => "01")

      port map(A => \long_reset\, Y => long_reset_i);
    
    \long_reset_cntr[2]\ : SLE
      port map(D => \long_reset_cntr_3[2]_net_1\, CLK => 
        \BIT_CLK\, EN => VCC_net_1, ALn => bd_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \long_reset_cntr[2]_net_1\);
    
    \long_reset_cntr[1]\ : SLE
      port map(D => \long_reset_cntr_3[1]_net_1\, CLK => 
        \BIT_CLK\, EN => VCC_net_1, ALn => bd_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \long_reset_cntr[1]_net_1\);
    
    \long_reset_cntr_3[0]\ : CFG3
      generic map(INIT => x"B3")

      port map(A => un2_long_reset_cntr_5, B => 
        \long_reset_cntr[0]_net_1\, C => un2_long_reset_cntr_4, Y
         => \long_reset_cntr_3[0]_net_1\);
    
    \long_reset_cntr[0]\ : SLE
      port map(D => \long_reset_cntr_3[0]_net_1\, CLK => 
        \BIT_CLK\, EN => VCC_net_1, ALn => bd_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \long_reset_cntr[0]_net_1\);
    
    TX_FIFO_UNDERRUN_set : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => un15_int_reg_clr, ALn => TX_FIFO_UNDERRUN_i, ADn
         => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \TX_FIFO_UNDERRUN_set\);
    
    \long_reset_cntr_3[4]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => un2_long_reset_cntr_4, B => 
        un2_long_reset_cntr_5, C => un4_long_reset_cntr_cry_4_S, 
        Y => \long_reset_cntr_3[4]_net_1\);
    
    FIFOS_INST : FIFOs
      port map(iRX_FIFO_Full(3) => \iRX_FIFO_Full[3]\, 
        iRX_FIFO_Full(2) => \iRX_FIFO_Full[2]\, iRX_FIFO_Full(1)
         => \iRX_FIFO_Full[1]\, iRX_FIFO_Full(0) => 
        \iRX_FIFO_Full[0]\, RX_FIFO_DIN_pipe(8) => 
        \RX_FIFO_DIN_pipe[8]\, RX_FIFO_DIN_pipe(7) => 
        \RX_FIFO_DIN_pipe[7]\, RX_FIFO_DIN_pipe(6) => 
        \RX_FIFO_DIN_pipe[6]\, RX_FIFO_DIN_pipe(5) => 
        \RX_FIFO_DIN_pipe[5]\, RX_FIFO_DIN_pipe(4) => 
        \RX_FIFO_DIN_pipe[4]\, RX_FIFO_DIN_pipe(3) => 
        \RX_FIFO_DIN_pipe[3]\, RX_FIFO_DIN_pipe(2) => 
        \RX_FIFO_DIN_pipe[2]\, RX_FIFO_DIN_pipe(1) => 
        \RX_FIFO_DIN_pipe[1]\, RX_FIFO_DIN_pipe(0) => 
        \RX_FIFO_DIN_pipe[0]\, CoreAPB3_0_APBmslave0_PWDATA(7)
         => CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), up_EOP_sync(2) => 
        \up_EOP_sync[2]\, up_EOP_sync(1) => \up_EOP_sync[1]\, 
        RX_FIFO_DOUT(7) => \RX_FIFO_DOUT[7]\, RX_FIFO_DOUT(6) => 
        \RX_FIFO_DOUT[6]\, RX_FIFO_DOUT(5) => \RX_FIFO_DOUT[5]\, 
        ReadFIFO_Read_Ptr(1) => \ReadFIFO_Read_Ptr[1]\, 
        ReadFIFO_Read_Ptr(0) => \ReadFIFO_Read_Ptr[0]\, 
        RX_FIFO_DOUT_3_0 => \RX_FIFO_DOUT_3[1]\, RX_FIFO_DOUT_2_0
         => \RX_FIFO_DOUT_2[1]\, RX_FIFO_DOUT_1_0 => 
        \RX_FIFO_DOUT_1[1]\, RX_FIFO_DOUT_0_0 => 
        \RX_FIFO_DOUT_0[1]\, N_674 => N_674, N_673 => N_673, 
        N_672 => N_672, N_667 => N_667, N_666 => N_666, N_665 => 
        N_665, N_660 => N_660, N_659 => N_659, N_658 => N_658, 
        iRX_FIFO_wr_en => iRX_FIFO_wr_en, sampler_clk1x_en => 
        sampler_clk1x_en, RX_InProcess_d1 => RX_InProcess_d1, 
        tx_col_detect_en => tx_col_detect_en, N_653 => N_653, 
        N_652 => N_652, N_651 => N_651, TX_FIFO_UNDERRUN => 
        TX_FIFO_UNDERRUN, TX_FIFO_UNDERRUN_i => 
        TX_FIFO_UNDERRUN_i, TX_FIFO_OVERFLOW => TX_FIFO_OVERFLOW, 
        TX_FIFO_OVERFLOW_i => TX_FIFO_OVERFLOW_i, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz, 
        TX_FIFO_Full => TX_FIFO_Full, TX_FIFO_wr_en => 
        TX_FIFO_wr_en, un1_tx_packet_length_0_sqmuxa_o => 
        un1_tx_packet_length_0_sqmuxa_o, TX_DataEn_1_o => 
        TX_DataEn_1_o, TX_PreAmble => TX_PreAmble, N_704 => N_704, 
        N_705 => N_705, N_706 => N_706, N_707 => N_707, N_708 => 
        N_708, N_709 => N_709, N_710 => N_710, N_711 => N_711, 
        byte_clk_en => \byte_clk_en\, TX_FIFO_Empty => 
        TX_FIFO_Empty, BIT_CLK => \BIT_CLK\, RX_FIFO_RST => 
        \RX_FIFO_RST\, RX_FIFO_rd_en => RX_FIFO_rd_en, 
        TX_FIFO_RST => TX_FIFO_RST, un2_apb3_reset => 
        un2_apb3_reset, rx_packet_complt => rx_packet_complt, 
        N_678 => N_678, N_712 => N_712, N_693 => N_693, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, 
        RX_FIFO_OVERFLOW_i => RX_FIFO_OVERFLOW_i, 
        RX_FIFO_OVERFLOW => RX_FIFO_OVERFLOW, RX_FIFO_UNDERRUN_i
         => RX_FIFO_UNDERRUN_i, RX_FIFO_UNDERRUN => 
        RX_FIFO_UNDERRUN);
    
    PROCESSOR_INTERFACE_INST : uP_if
      port map(RX_FIFO_DIN(3) => \RX_FIFO_DIN[3]\, RX_FIFO_DIN(2)
         => \RX_FIFO_DIN[2]\, rx_crc_data_calc(11) => 
        \rx_crc_data_calc[11]\, rx_crc_data_calc(10) => 
        \rx_crc_data_calc[10]\, CoreAPB3_0_APBmslave0_PADDR(7)
         => CoreAPB3_0_APBmslave0_PADDR(7), 
        CoreAPB3_0_APBmslave0_PADDR(6) => 
        CoreAPB3_0_APBmslave0_PADDR(6), 
        CoreAPB3_0_APBmslave0_PADDR(5) => 
        CoreAPB3_0_APBmslave0_PADDR(5), 
        CoreAPB3_0_APBmslave0_PADDR(4) => 
        CoreAPB3_0_APBmslave0_PADDR(4), 
        CoreAPB3_0_APBmslave0_PADDR(3) => 
        CoreAPB3_0_APBmslave0_PADDR(3), 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        CoreAPB3_0_APBmslave0_PADDR(2), 
        CoreAPB3_0_APBmslave0_PADDR(1) => 
        CoreAPB3_0_APBmslave0_PADDR(1), 
        CoreAPB3_0_APBmslave0_PADDR(0) => 
        CoreAPB3_0_APBmslave0_PADDR(0), 
        CoreAPB3_0_APBmslave0_PRDATA_m(7) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(7), 
        CoreAPB3_0_APBmslave0_PRDATA_m(6) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(6), 
        CoreAPB3_0_APBmslave0_PRDATA_m(5) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(5), 
        CoreAPB3_0_APBmslave0_PRDATA_m(4) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(4), 
        CoreAPB3_0_APBmslave0_PRDATA_m(3) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(3), 
        CoreAPB3_0_APBmslave0_PRDATA_m(2) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(2), 
        CoreAPB3_0_APBmslave0_PRDATA_m(1) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(1), 
        CoreAPB3_0_APBmslave0_PRDATA_m(0) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(0), RX_FIFO_DOUT(7) => 
        \RX_FIFO_DOUT[7]\, RX_FIFO_DOUT(6) => \RX_FIFO_DOUT[6]\, 
        RX_FIFO_DOUT(5) => \RX_FIFO_DOUT[5]\, iRX_FIFO_Full(3)
         => \iRX_FIFO_Full[3]\, iRX_FIFO_Full(2) => 
        \iRX_FIFO_Full[2]\, iRX_FIFO_Full(1) => 
        \iRX_FIFO_Full[1]\, iRX_FIFO_Full(0) => 
        \iRX_FIFO_Full[0]\, ReadFIFO_Read_Ptr(1) => 
        \ReadFIFO_Read_Ptr[1]\, ReadFIFO_Read_Ptr(0) => 
        \ReadFIFO_Read_Ptr[0]\, consumer_type4_reg(9) => 
        \consumer_type4_reg[9]\, consumer_type4_reg(8) => 
        \consumer_type4_reg[8]\, consumer_type4_reg(7) => 
        \consumer_type4_reg[7]\, consumer_type4_reg(6) => 
        \consumer_type4_reg[6]\, consumer_type4_reg(5) => 
        \consumer_type4_reg[5]\, consumer_type4_reg(4) => 
        \consumer_type4_reg[4]\, consumer_type4_reg(3) => 
        \consumer_type4_reg[3]\, consumer_type4_reg(2) => 
        \consumer_type4_reg[2]\, consumer_type4_reg(1) => 
        \consumer_type4_reg[1]\, consumer_type4_reg(0) => 
        \consumer_type4_reg[0]\, consumer_type3_reg(9) => 
        \consumer_type3_reg[9]\, consumer_type3_reg(8) => 
        \consumer_type3_reg[8]\, consumer_type3_reg(7) => 
        \consumer_type3_reg[7]\, consumer_type3_reg(6) => 
        \consumer_type3_reg[6]\, consumer_type3_reg(5) => 
        \consumer_type3_reg[5]\, consumer_type3_reg(4) => 
        \consumer_type3_reg[4]\, consumer_type3_reg(3) => 
        \consumer_type3_reg[3]\, consumer_type3_reg(2) => 
        \consumer_type3_reg[2]\, consumer_type3_reg(1) => 
        \consumer_type3_reg[1]\, consumer_type3_reg(0) => 
        \consumer_type3_reg[0]\, consumer_type2_reg(9) => 
        \consumer_type2_reg[9]\, consumer_type2_reg(8) => 
        \consumer_type2_reg[8]\, consumer_type2_reg(7) => 
        \consumer_type2_reg[7]\, consumer_type2_reg(6) => 
        \consumer_type2_reg[6]\, consumer_type2_reg(5) => 
        \consumer_type2_reg[5]\, consumer_type2_reg(4) => 
        \consumer_type2_reg[4]\, consumer_type2_reg(3) => 
        \consumer_type2_reg[3]\, consumer_type2_reg(2) => 
        \consumer_type2_reg[2]\, consumer_type2_reg(1) => 
        \consumer_type2_reg[1]\, consumer_type2_reg(0) => 
        \consumer_type2_reg[0]\, consumer_type1_reg(9) => 
        \consumer_type1_reg[9]\, consumer_type1_reg(8) => 
        \consumer_type1_reg[8]\, consumer_type1_reg(7) => 
        \consumer_type1_reg[7]\, consumer_type1_reg(6) => 
        \consumer_type1_reg[6]\, consumer_type1_reg(5) => 
        \consumer_type1_reg[5]\, consumer_type1_reg(4) => 
        \consumer_type1_reg[4]\, consumer_type1_reg(3) => 
        \consumer_type1_reg[3]\, consumer_type1_reg(2) => 
        \consumer_type1_reg[2]\, consumer_type1_reg(1) => 
        \consumer_type1_reg[1]\, consumer_type1_reg(0) => 
        \consumer_type1_reg[0]\, CoreAPB3_0_APBmslave0_PWDATA(7)
         => CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), up_EOP_sync(2) => 
        \up_EOP_sync[2]\, up_EOP_sync(1) => \up_EOP_sync[1]\, 
        lfsr_c_i_i_0 => \lfsr_c_i_i[4]\, RX_FIFO_DIN_pipe_0 => 
        \RX_FIFO_DIN_pipe[8]\, RX_FIFO_DOUT_1_0 => 
        \RX_FIFO_DOUT_1[1]\, RX_FIFO_DOUT_0_0 => 
        \RX_FIFO_DOUT_0[1]\, RX_FIFO_DOUT_3_0 => 
        \RX_FIFO_DOUT_3[1]\, RX_FIFO_DOUT_2_0 => 
        \RX_FIFO_DOUT_2[1]\, un2_apb3_reset_set => 
        un2_apb3_reset_set, un2_apb3_reset_i => un2_apb3_reset_i, 
        BIT_CLK => \BIT_CLK\, tx_packet_complt => 
        tx_packet_complt, rx_CRC_error_set => \rx_CRC_error_set\, 
        un31_int_reg_clr => un31_int_reg_clr, rx_CRC_error => 
        rx_CRC_error, RX_FIFO_OVERFLOW_set => 
        \RX_FIFO_OVERFLOW_set\, un27_int_reg_clr => 
        un27_int_reg_clr, RX_FIFO_OVERFLOW => RX_FIFO_OVERFLOW, 
        RX_FIFO_UNDERRUN_set => \RX_FIFO_UNDERRUN_set\, 
        un23_int_reg_clr => un23_int_reg_clr, RX_FIFO_UNDERRUN
         => RX_FIFO_UNDERRUN, TX_FIFO_OVERFLOW_set => 
        \TX_FIFO_OVERFLOW_set\, un19_int_reg_clr => 
        un19_int_reg_clr, TX_FIFO_OVERFLOW => TX_FIFO_OVERFLOW, 
        TX_FIFO_UNDERRUN_set => \TX_FIFO_UNDERRUN_set\, 
        un15_int_reg_clr => un15_int_reg_clr, TX_FIFO_UNDERRUN
         => TX_FIFO_UNDERRUN, un2_apb3_reset => un2_apb3_reset, 
        CommsFPGA_top_0_INT => CommsFPGA_top_0_INT, TX_PreAmble
         => TX_PreAmble, N_712 => N_712, N_855_i => N_855_i, 
        CoreAPB3_0_APBmslave0_PWRITE => 
        CoreAPB3_0_APBmslave0_PWRITE, N_993_i => N_993_i, 
        sampler_clk1x_en => sampler_clk1x_en, SM_advance_i => 
        SM_advance_i, N_41_i => N_41_i, rx_crc_HighByte_en => 
        rx_crc_HighByte_en, N_535 => N_535, 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i => 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i, 
        CoreAPB3_0_APBmslave0_PENABLE => 
        CoreAPB3_0_APBmslave0_PENABLE, RX_FIFO_RST_1 => 
        RX_FIFO_RST_1, RX_EarlyTerm => RX_EarlyTerm, 
        CoreAPB3_0_APBmslave0_PSELx => 
        CoreAPB3_0_APBmslave0_PSELx, TX_FIFO_Empty => 
        TX_FIFO_Empty, TX_FIFO_Full => TX_FIFO_Full, N_693 => 
        N_693, N_678 => N_678, N_658 => N_658, N_651 => N_651, 
        N_672 => N_672, N_665 => N_665, N_659 => N_659, N_652 => 
        N_652, N_673 => N_673, N_666 => N_666, N_660 => N_660, 
        N_653 => N_653, N_674 => N_674, N_667 => N_667, 
        rx_packet_complt => rx_packet_complt, RX_FIFO_rd_en => 
        RX_FIFO_rd_en, TX_FIFO_wr_en => TX_FIFO_wr_en, N_855_i_i
         => N_855_i_i, TX_FIFO_RST => TX_FIFO_RST, start_tx_FIFO
         => start_tx_FIFO, internal_loopback => internal_loopback, 
        external_loopback => external_loopback, long_reset => 
        \long_reset\, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, long_reset_set => 
        \long_reset_set\, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, long_reset_i => long_reset_i);
    
    bd_reset_RNIK1J6 : CLKINT
      port map(A => \bd_reset\, Y => bd_reset_i);
    
    RX_FIFO_UNDERRUN_set : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => un23_int_reg_clr, ALn => RX_FIFO_UNDERRUN_i, ADn
         => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_UNDERRUN_set\);
    
    \long_reset_cntr[4]\ : SLE
      port map(D => \long_reset_cntr_3[4]_net_1\, CLK => 
        \BIT_CLK\, EN => VCC_net_1, ALn => bd_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \long_reset_cntr[4]_net_1\);
    
    RESET_RNIFEG6_0 : CFG1
      generic map(INIT => "01")

      port map(A => un2_apb3_reset, Y => un2_apb3_reset_i);
    
    \ClkDivider[1]\ : SLE
      port map(D => \ClkDivider_RNO[1]_net_1\, CLK => \BIT_CLK\, 
        EN => VCC_net_1, ALn => bd_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ClkDivider[1]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som is

    port( DEBOUNCE_IN           : in    std_logic_vector(2 downto 0);
          ID_RES                : in    std_logic_vector(3 downto 0);
          MAC_MII_RXD           : in    std_logic_vector(3 downto 0);
          MAC_MII_TXD           : out   std_logic_vector(3 downto 0);
          MDDR_ADDR             : out   std_logic_vector(15 downto 0);
          MDDR_BA               : out   std_logic_vector(2 downto 0);
          GPIO_1_BI             : inout std_logic_vector(0 to 0) := (others => 'Z');
          GPIO_1_BIDI           : in    std_logic_vector(0 to 0);
          GPIO_6_PAD            : inout std_logic_vector(0 to 0) := (others => 'Z');
          GPIO_7_PADI           : inout std_logic_vector(0 to 0) := (others => 'Z');
          MDDR_DM_RDQS          : inout std_logic_vector(1 downto 0) := (others => 'Z');
          MDDR_DQ               : inout std_logic_vector(15 downto 0) := (others => 'Z');
          MDDR_DQS              : inout std_logic_vector(1 downto 0) := (others => 'Z');
          SPI_1_CLK             : inout std_logic_vector(0 to 0) := (others => 'Z');
          SPI_1_SS0_CAM         : inout std_logic_vector(0 to 0) := (others => 'Z');
          SPI_1_SS0_OTH         : inout std_logic_vector(0 to 0) := (others => 'Z');
          DEVRST_N              : in    std_logic;
          MAC_MII_COL           : in    std_logic;
          MAC_MII_CRS           : in    std_logic;
          MAC_MII_RX_CLK        : in    std_logic;
          MAC_MII_RX_DV         : in    std_logic;
          MAC_MII_RX_ER         : in    std_logic;
          MAC_MII_TX_CLK        : in    std_logic;
          MANCHESTER_IN         : in    std_logic;
          MDDR_DQS_TMATCH_0_IN  : in    std_logic;
          MMUART_0_RXD_F2M      : in    std_logic;
          MMUART_1_RXD          : in    std_logic;
          PULLDOWN_R9           : in    std_logic;
          SPI_0_DI              : in    std_logic;
          SPI_1_DI_CAM          : in    std_logic;
          SPI_1_DI_OTH          : in    std_logic;
          XTL                   : in    std_logic;
          DEBOUNCE_OUT_1        : out   std_logic;
          DEBOUNCE_OUT_2        : out   std_logic;
          DRVR_EN               : out   std_logic;
          Data_FAIL             : out   std_logic;
          GPIO_11_M2F           : out   std_logic;
          GPIO_20_OUT           : out   std_logic;
          GPIO_21_M2F           : out   std_logic;
          GPIO_22_M2F           : out   std_logic;
          GPIO_24_M2F           : out   std_logic;
          GPIO_5_M2F            : out   std_logic;
          GPIO_8_M2F            : out   std_logic;
          MAC_MII_MDC           : out   std_logic;
          MAC_MII_TX_EN         : out   std_logic;
          MANCH_OUT_N           : out   std_logic;
          MANCH_OUT_P           : out   std_logic;
          MDDR_CAS_N            : out   std_logic;
          MDDR_CKE              : out   std_logic;
          MDDR_CLK              : out   std_logic;
          MDDR_CLK_N            : out   std_logic;
          MDDR_CS_N             : out   std_logic;
          MDDR_DQS_TMATCH_0_OUT : out   std_logic;
          MDDR_ODT              : out   std_logic;
          MDDR_RAS_N            : out   std_logic;
          MDDR_RESET_N          : out   std_logic;
          MDDR_WE_N             : out   std_logic;
          MMUART_0_TXD_M2F      : out   std_logic;
          MMUART_1_TXD          : out   std_logic;
          RCVR_EN               : out   std_logic;
          SPI_0_DO              : out   std_logic;
          SPI_0_SS1             : out   std_logic;
          SPI_1_DO_CAM          : out   std_logic;
          SPI_1_DO_OTH          : out   std_logic;
          GPIO_0_BI             : inout std_logic := 'Z';
          GPIO_12_BI            : inout std_logic := 'Z';
          GPIO_14_BI            : inout std_logic := 'Z';
          GPIO_15_BI            : inout std_logic := 'Z';
          GPIO_16_BI            : inout std_logic := 'Z';
          GPIO_17_BI            : inout std_logic := 'Z';
          GPIO_18_BI            : inout std_logic := 'Z';
          GPIO_25_BI            : inout std_logic := 'Z';
          GPIO_26_BI            : inout std_logic := 'Z';
          GPIO_31_BI            : inout std_logic := 'Z';
          GPIO_3_BI             : inout std_logic := 'Z';
          GPIO_4_BI             : inout std_logic := 'Z';
          I2C_1_SCL             : inout std_logic := 'Z';
          I2C_1_SDA             : inout std_logic := 'Z';
          MAC_MII_MDIO          : inout std_logic := 'Z';
          SPI_0_CLK             : inout std_logic := 'Z';
          SPI_0_SS0             : inout std_logic := 'Z'
        );

end m2s010_som;

architecture DEF_ARCH of m2s010_som is 

  component OUTBUF
    generic (IOSTD:string := "");

    port( D   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component INBUF
    generic (IOSTD:string := "");

    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component CoreAPB3
    port( m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR : in    std_logic_vector(15 downto 12) := (others => 'U');
          CoreAPB3_0_APBmslave0_PSELx            : out   std_logic;
          m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component m2s010_som_CommsFPGA_CCC_0_FCCC
    port( m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC : in    std_logic := 'U';
          CommsFPGA_CCC_0_LOCK                      : out   std_logic;
          CommsFPGA_CCC_0_GL1                       : out   std_logic;
          CommsFPGA_CCC_0_GL0                       : out   std_logic
        );
  end component;

  component m2s010_som_ID_RES_0_IO
    port( ID_RES  : in    std_logic_vector(3 downto 0) := (others => 'U');
          Y_net_0 : out   std_logic_vector(3 downto 0)
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component m2s010_som_sb
    port( MDDR_DQS                                  : inout   std_logic_vector(1 downto 0);
          MDDR_DQ                                   : inout   std_logic_vector(15 downto 0);
          MDDR_DM_RDQS                              : inout   std_logic_vector(1 downto 0);
          MDDR_BA                                   : out   std_logic_vector(2 downto 0);
          MDDR_ADDR                                 : out   std_logic_vector(15 downto 0);
          CoreAPB3_0_APBmslave0_PADDR               : out   std_logic_vector(7 downto 0);
          m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR    : out   std_logic_vector(15 downto 12);
          CoreAPB3_0_APBmslave0_PWDATA              : out   std_logic_vector(7 downto 0);
          MAC_MII_TXD_c                             : out   std_logic_vector(3 downto 0);
          CoreAPB3_0_APBmslave0_PRDATA_m            : in    std_logic_vector(7 downto 0) := (others => 'U');
          Y_net_0                                   : in    std_logic_vector(3 downto 0) := (others => 'U');
          MAC_MII_RXD_c                             : in    std_logic_vector(3 downto 0) := (others => 'U');
          SPI_1_SS0_OTH_0                           : inout   std_logic;
          DEBOUNCE_OUT_net_0_0                      : in    std_logic := 'U';
          GPIO_7_PADI_0                             : inout   std_logic;
          GPIO_6_PAD_0                              : inout   std_logic;
          GPIO_1_BI_0                               : inout   std_logic;
          SPI_1_SS0_CAM_0                           : inout   std_logic;
          SPI_1_CLK_0                               : inout   std_logic;
          SPI_0_SS1                                 : out   std_logic;
          SPI_0_SS0                                 : inout   std_logic;
          SPI_0_DO                                  : out   std_logic;
          SPI_0_DI                                  : in    std_logic := 'U';
          SPI_0_CLK                                 : inout   std_logic;
          MMUART_1_TXD                              : out   std_logic;
          MMUART_1_RXD                              : in    std_logic := 'U';
          MDDR_WE_N                                 : out   std_logic;
          MDDR_RESET_N                              : out   std_logic;
          MDDR_RAS_N                                : out   std_logic;
          MDDR_ODT                                  : out   std_logic;
          MDDR_DQS_TMATCH_0_OUT                     : out   std_logic;
          MDDR_DQS_TMATCH_0_IN                      : in    std_logic := 'U';
          MDDR_CS_N                                 : out   std_logic;
          MDDR_CKE                                  : out   std_logic;
          MDDR_CAS_N                                : out   std_logic;
          I2C_1_SDA                                 : inout   std_logic;
          I2C_1_SCL                                 : inout   std_logic;
          GPIO_31_BI                                : inout   std_logic;
          GPIO_26_BI                                : inout   std_logic;
          GPIO_25_BI                                : inout   std_logic;
          GPIO_20_OUT                               : out   std_logic;
          GPIO_18_BI                                : inout   std_logic;
          GPIO_17_BI                                : inout   std_logic;
          GPIO_16_BI                                : inout   std_logic;
          GPIO_15_BI                                : inout   std_logic;
          GPIO_14_BI                                : inout   std_logic;
          GPIO_12_BI                                : inout   std_logic;
          GPIO_4_BI                                 : inout   std_logic;
          GPIO_3_BI                                 : inout   std_logic;
          GPIO_0_BI                                 : inout   std_logic;
          CoreAPB3_0_APBmslave0_PENABLE             : out   std_logic;
          m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx    : out   std_logic;
          CoreAPB3_0_APBmslave0_PWRITE              : out   std_logic;
          MAC_MII_MDC_c                             : out   std_logic;
          GPIO_22_M2F_c                             : out   std_logic;
          GPIO_21_M2F_c                             : out   std_logic;
          m2s010_som_sb_0_GPIO_28_SW_RESET          : out   std_logic;
          MMUART_0_TXD_M2F_c                        : out   std_logic;
          GPIO_24_M2F_c                             : out   std_logic;
          GPIO_5_M2F_c                              : out   std_logic;
          GPIO_8_M2F_c                              : out   std_logic;
          GPIO_11_M2F_c                             : out   std_logic;
          MAC_MII_TX_EN_c                           : out   std_logic;
          MAC_MII_COL_c                             : in    std_logic := 'U';
          MAC_MII_CRS_c                             : in    std_logic := 'U';
          CommsFPGA_top_0_INT                       : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PREADY_i_m_i        : in    std_logic := 'U';
          DEBOUNCE_OUT_1_c                          : in    std_logic := 'U';
          DEBOUNCE_OUT_2_c                          : in    std_logic := 'U';
          MMUART_0_RXD_F2M_c                        : in    std_logic := 'U';
          MAC_MII_RX_CLK_c                          : in    std_logic := 'U';
          MAC_MII_RX_DV_c                           : in    std_logic := 'U';
          MAC_MII_RX_ER_c                           : in    std_logic := 'U';
          MAC_MII_TX_CLK_c                          : in    std_logic := 'U';
          MDDR_CLK_N                                : out   std_logic;
          MDDR_CLK                                  : out   std_logic;
          XTL                                       : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz                 : out   std_logic;
          m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC : inout   std_logic;
          SPI_1_DI_CAM_c                            : in    std_logic := 'U';
          SPI_1_DI_OTH_c                            : in    std_logic := 'U';
          CommsFPGA_top_0_CAMERA_NODE               : in    std_logic := 'U';
          DEVRST_N                                  : in    std_logic := 'U';
          m2s010_som_sb_0_POWER_ON_RESET_N          : out   std_logic;
          MAC_MII_MDIO                              : inout   std_logic;
          SPI_1_DO_CAM_c                            : inout   std_logic;
          SPI_1_DO_OTH                              : out   std_logic
        );
  end component;

  component CommsFPGA_top
    port( CoreAPB3_0_APBmslave0_PWDATA       : in    std_logic_vector(7 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PRDATA_m     : out   std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PADDR        : in    std_logic_vector(7 downto 0) := (others => 'U');
          DEBOUNCE_IN_c                      : in    std_logic_vector(2 downto 0) := (others => 'U');
          Y_net_0                            : in    std_logic_vector(3 downto 1) := (others => 'U');
          DEBOUNCE_OUT_net_0_0               : out   std_logic;
          MANCHESTER_IN_c                    : in    std_logic := 'U';
          MANCH_OUT_P_c                      : out   std_logic;
          MANCH_OUT_P_c_i                    : out   std_logic;
          DRVR_EN_c                          : out   std_logic;
          N_855_i_i                          : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PSELx        : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PENABLE      : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PREADY_i_m_i : out   std_logic;
          CoreAPB3_0_APBmslave0_PWRITE       : in    std_logic := 'U';
          N_855_i                            : out   std_logic;
          CommsFPGA_top_0_INT                : out   std_logic;
          DEBOUNCE_OUT_1_c                   : out   std_logic;
          DEBOUNCE_OUT_2_c                   : out   std_logic;
          CommsFPGA_top_0_CAMERA_NODE        : out   std_logic;
          m2s010_som_sb_0_POWER_ON_RESET_N   : in    std_logic := 'U';
          m2s010_som_sb_0_GPIO_28_SW_RESET   : in    std_logic := 'U';
          CommsFPGA_CCC_0_LOCK               : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL1                : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0                : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz          : in    std_logic := 'U'
        );
  end component;

    signal m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC, 
        CommsFPGA_CCC_0_LOCK, CommsFPGA_CCC_0_GL0, 
        CommsFPGA_CCC_0_GL1, m2s010_som_sb_0_GPIO_28_SW_RESET, 
        m2s010_som_sb_0_POWER_ON_RESET_N, 
        m2s010_som_sb_0_CCC_71MHz, \Y_net_0[0]\, \Y_net_0[1]\, 
        \Y_net_0[2]\, \Y_net_0[3]\, CommsFPGA_top_0_CAMERA_NODE, 
        CommsFPGA_top_0_INT, \DEBOUNCE_OUT_net_0[0]\, GND_net_1, 
        \CoreAPB3_0_APBmslave0_PADDR[0]\, 
        \CoreAPB3_0_APBmslave0_PADDR[1]\, 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, 
        \CoreAPB3_0_APBmslave0_PADDR[4]\, 
        \CoreAPB3_0_APBmslave0_PADDR[5]\, 
        \CoreAPB3_0_APBmslave0_PADDR[6]\, 
        \CoreAPB3_0_APBmslave0_PADDR[7]\, 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[12]\, 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[13]\, 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[14]\, 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[15]\, 
        CoreAPB3_0_APBmslave0_PWRITE, 
        CoreAPB3_0_APBmslave0_PENABLE, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx, 
        \CoreAPB3_0_APBmslave0_PWDATA[0]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[1]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[2]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[3]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[4]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[5]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[6]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[7]\, VCC_net_1, 
        \CoreAPB3_0_APBmslave0_PRDATA_m[0]\, 
        \CoreAPB3_0_APBmslave0_PRDATA_m[1]\, 
        \CoreAPB3_0_APBmslave0_PRDATA_m[2]\, 
        \CoreAPB3_0_APBmslave0_PRDATA_m[3]\, 
        \CoreAPB3_0_APBmslave0_PRDATA_m[4]\, 
        \CoreAPB3_0_APBmslave0_PRDATA_m[5]\, 
        \CoreAPB3_0_APBmslave0_PRDATA_m[6]\, 
        \CoreAPB3_0_APBmslave0_PRDATA_m[7]\, 
        CoreAPB3_0_APBmslave0_PSELx, \DEBOUNCE_IN_c[0]\, 
        \DEBOUNCE_IN_c[1]\, \DEBOUNCE_IN_c[2]\, MAC_MII_COL_c, 
        MAC_MII_CRS_c, \MAC_MII_RXD_c[0]\, \MAC_MII_RXD_c[1]\, 
        \MAC_MII_RXD_c[2]\, \MAC_MII_RXD_c[3]\, MAC_MII_RX_CLK_c, 
        MAC_MII_RX_DV_c, MAC_MII_RX_ER_c, MAC_MII_TX_CLK_c, 
        MANCHESTER_IN_c, MMUART_0_RXD_F2M_c, Data_FAIL_c, 
        SPI_1_DI_CAM_c, SPI_1_DI_OTH_c, DEBOUNCE_OUT_1_c, 
        DEBOUNCE_OUT_2_c, DRVR_EN_c, GPIO_11_M2F_c, GPIO_21_M2F_c, 
        GPIO_22_M2F_c, GPIO_24_M2F_c, GPIO_5_M2F_c, GPIO_8_M2F_c, 
        MAC_MII_MDC_c, \MAC_MII_TXD_c[0]\, \MAC_MII_TXD_c[1]\, 
        \MAC_MII_TXD_c[2]\, \MAC_MII_TXD_c[3]\, MAC_MII_TX_EN_c, 
        MANCH_OUT_P_c, MMUART_0_TXD_M2F_c, SPI_1_DO_CAM_c, 
        MANCH_OUT_P_c_i, CoreAPB3_0_APBmslave0_PREADY_i_m_i, 
        \CommsFPGA_top_0.N_855_i_i\, N_855_i : std_logic;

    for all : CoreAPB3
	Use entity work.CoreAPB3(DEF_ARCH);
    for all : m2s010_som_CommsFPGA_CCC_0_FCCC
	Use entity work.m2s010_som_CommsFPGA_CCC_0_FCCC(DEF_ARCH);
    for all : m2s010_som_ID_RES_0_IO
	Use entity work.m2s010_som_ID_RES_0_IO(DEF_ARCH);
    for all : m2s010_som_sb
	Use entity work.m2s010_som_sb(DEF_ARCH);
    for all : CommsFPGA_top
	Use entity work.CommsFPGA_top(DEF_ARCH);
begin 


    RCVR_EN_obuf : OUTBUF
      port map(D => VCC_net_1, PAD => RCVR_EN);
    
    MANCH_OUT_N_obuf : OUTBUF
      port map(D => MANCH_OUT_P_c_i, PAD => MANCH_OUT_N);
    
    \MAC_MII_RXD_ibuf[1]\ : INBUF
      port map(PAD => MAC_MII_RXD(1), Y => \MAC_MII_RXD_c[1]\);
    
    MMUART_0_RXD_F2M_ibuf : INBUF
      port map(PAD => MMUART_0_RXD_F2M, Y => MMUART_0_RXD_F2M_c);
    
    MAC_MII_RX_CLK_ibuf : INBUF
      port map(PAD => MAC_MII_RX_CLK, Y => MAC_MII_RX_CLK_c);
    
    MAC_MII_CRS_ibuf : INBUF
      port map(PAD => MAC_MII_CRS, Y => MAC_MII_CRS_c);
    
    CoreAPB3_0 : CoreAPB3
      port map(m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(15) => 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[15]\, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(14) => 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[14]\, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(13) => 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[13]\, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(12) => 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[12]\, 
        CoreAPB3_0_APBmslave0_PSELx => 
        CoreAPB3_0_APBmslave0_PSELx, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    CommsFPGA_CCC_0 : m2s010_som_CommsFPGA_CCC_0_FCCC
      port map(m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC => 
        m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC, 
        CommsFPGA_CCC_0_LOCK => CommsFPGA_CCC_0_LOCK, 
        CommsFPGA_CCC_0_GL1 => CommsFPGA_CCC_0_GL1, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0);
    
    MAC_MII_TX_EN_obuf : OUTBUF
      port map(D => MAC_MII_TX_EN_c, PAD => MAC_MII_TX_EN);
    
    MAC_MII_TX_CLK_ibuf : INBUF
      port map(PAD => MAC_MII_TX_CLK, Y => MAC_MII_TX_CLK_c);
    
    \MAC_MII_TXD_obuf[1]\ : OUTBUF
      port map(D => \MAC_MII_TXD_c[1]\, PAD => MAC_MII_TXD(1));
    
    DEBOUNCE_OUT_2_obuf : OUTBUF
      port map(D => DEBOUNCE_OUT_2_c, PAD => DEBOUNCE_OUT_2);
    
    ID_RES_0 : m2s010_som_ID_RES_0_IO
      port map(ID_RES(3) => ID_RES(3), ID_RES(2) => ID_RES(2), 
        ID_RES(1) => ID_RES(1), ID_RES(0) => ID_RES(0), 
        Y_net_0(3) => \Y_net_0[3]\, Y_net_0(2) => \Y_net_0[2]\, 
        Y_net_0(1) => \Y_net_0[1]\, Y_net_0(0) => \Y_net_0[0]\);
    
    \MAC_MII_RXD_ibuf[0]\ : INBUF
      port map(PAD => MAC_MII_RXD(0), Y => \MAC_MII_RXD_c[0]\);
    
    MMUART_0_TXD_M2F_obuf : OUTBUF
      port map(D => MMUART_0_TXD_M2F_c, PAD => MMUART_0_TXD_M2F);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \MAC_MII_RXD_ibuf[3]\ : INBUF
      port map(PAD => MAC_MII_RXD(3), Y => \MAC_MII_RXD_c[3]\);
    
    SPI_1_DI_CAM_ibuf : INBUF
      port map(PAD => SPI_1_DI_CAM, Y => SPI_1_DI_CAM_c);
    
    \MAC_MII_TXD_obuf[0]\ : OUTBUF
      port map(D => \MAC_MII_TXD_c[0]\, PAD => MAC_MII_TXD(0));
    
    Data_FAIL_obuf : OUTBUF
      port map(D => Data_FAIL_c, PAD => Data_FAIL);
    
    MAC_MII_COL_ibuf : INBUF
      port map(PAD => MAC_MII_COL, Y => MAC_MII_COL_c);
    
    MANCH_OUT_P_obuf : OUTBUF
      port map(D => MANCH_OUT_P_c, PAD => MANCH_OUT_P);
    
    MAC_MII_MDC_obuf : OUTBUF
      port map(D => MAC_MII_MDC_c, PAD => MAC_MII_MDC);
    
    MANCHESTER_IN_ibuf : INBUF
      port map(PAD => MANCHESTER_IN, Y => MANCHESTER_IN_c);
    
    I_404 : CLKINT
      port map(A => N_855_i, Y => \CommsFPGA_top_0.N_855_i_i\);
    
    GPIO_22_M2F_obuf : OUTBUF
      port map(D => GPIO_22_M2F_c, PAD => GPIO_22_M2F);
    
    GPIO_21_M2F_obuf : OUTBUF
      port map(D => GPIO_21_M2F_c, PAD => GPIO_21_M2F);
    
    SPI_1_DO_CAM_obuf : OUTBUF
      port map(D => SPI_1_DO_CAM_c, PAD => SPI_1_DO_CAM);
    
    \MAC_MII_TXD_obuf[3]\ : OUTBUF
      port map(D => \MAC_MII_TXD_c[3]\, PAD => MAC_MII_TXD(3));
    
    \DEBOUNCE_IN_ibuf[1]\ : INBUF
      port map(PAD => DEBOUNCE_IN(1), Y => \DEBOUNCE_IN_c[1]\);
    
    MAC_MII_RX_DV_ibuf : INBUF
      port map(PAD => MAC_MII_RX_DV, Y => MAC_MII_RX_DV_c);
    
    DRVR_EN_obuf : OUTBUF
      port map(D => DRVR_EN_c, PAD => DRVR_EN);
    
    DEBOUNCE_OUT_1_obuf : OUTBUF
      port map(D => DEBOUNCE_OUT_1_c, PAD => DEBOUNCE_OUT_1);
    
    SPI_1_DI_OTH_ibuf : INBUF
      port map(PAD => SPI_1_DI_OTH, Y => SPI_1_DI_OTH_c);
    
    m2s010_som_sb_0 : m2s010_som_sb
      port map(MDDR_DQS(1) => MDDR_DQS(1), MDDR_DQS(0) => 
        MDDR_DQS(0), MDDR_DQ(15) => MDDR_DQ(15), MDDR_DQ(14) => 
        MDDR_DQ(14), MDDR_DQ(13) => MDDR_DQ(13), MDDR_DQ(12) => 
        MDDR_DQ(12), MDDR_DQ(11) => MDDR_DQ(11), MDDR_DQ(10) => 
        MDDR_DQ(10), MDDR_DQ(9) => MDDR_DQ(9), MDDR_DQ(8) => 
        MDDR_DQ(8), MDDR_DQ(7) => MDDR_DQ(7), MDDR_DQ(6) => 
        MDDR_DQ(6), MDDR_DQ(5) => MDDR_DQ(5), MDDR_DQ(4) => 
        MDDR_DQ(4), MDDR_DQ(3) => MDDR_DQ(3), MDDR_DQ(2) => 
        MDDR_DQ(2), MDDR_DQ(1) => MDDR_DQ(1), MDDR_DQ(0) => 
        MDDR_DQ(0), MDDR_DM_RDQS(1) => MDDR_DM_RDQS(1), 
        MDDR_DM_RDQS(0) => MDDR_DM_RDQS(0), MDDR_BA(2) => 
        MDDR_BA(2), MDDR_BA(1) => MDDR_BA(1), MDDR_BA(0) => 
        MDDR_BA(0), MDDR_ADDR(15) => MDDR_ADDR(15), MDDR_ADDR(14)
         => MDDR_ADDR(14), MDDR_ADDR(13) => MDDR_ADDR(13), 
        MDDR_ADDR(12) => MDDR_ADDR(12), MDDR_ADDR(11) => 
        MDDR_ADDR(11), MDDR_ADDR(10) => MDDR_ADDR(10), 
        MDDR_ADDR(9) => MDDR_ADDR(9), MDDR_ADDR(8) => 
        MDDR_ADDR(8), MDDR_ADDR(7) => MDDR_ADDR(7), MDDR_ADDR(6)
         => MDDR_ADDR(6), MDDR_ADDR(5) => MDDR_ADDR(5), 
        MDDR_ADDR(4) => MDDR_ADDR(4), MDDR_ADDR(3) => 
        MDDR_ADDR(3), MDDR_ADDR(2) => MDDR_ADDR(2), MDDR_ADDR(1)
         => MDDR_ADDR(1), MDDR_ADDR(0) => MDDR_ADDR(0), 
        CoreAPB3_0_APBmslave0_PADDR(7) => 
        \CoreAPB3_0_APBmslave0_PADDR[7]\, 
        CoreAPB3_0_APBmslave0_PADDR(6) => 
        \CoreAPB3_0_APBmslave0_PADDR[6]\, 
        CoreAPB3_0_APBmslave0_PADDR(5) => 
        \CoreAPB3_0_APBmslave0_PADDR[5]\, 
        CoreAPB3_0_APBmslave0_PADDR(4) => 
        \CoreAPB3_0_APBmslave0_PADDR[4]\, 
        CoreAPB3_0_APBmslave0_PADDR(3) => 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, 
        CoreAPB3_0_APBmslave0_PADDR(1) => 
        \CoreAPB3_0_APBmslave0_PADDR[1]\, 
        CoreAPB3_0_APBmslave0_PADDR(0) => 
        \CoreAPB3_0_APBmslave0_PADDR[0]\, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(15) => 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[15]\, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(14) => 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[14]\, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(13) => 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[13]\, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(12) => 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[12]\, 
        CoreAPB3_0_APBmslave0_PWDATA(7) => 
        \CoreAPB3_0_APBmslave0_PWDATA[7]\, 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        \CoreAPB3_0_APBmslave0_PWDATA[6]\, 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        \CoreAPB3_0_APBmslave0_PWDATA[5]\, 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        \CoreAPB3_0_APBmslave0_PWDATA[4]\, 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        \CoreAPB3_0_APBmslave0_PWDATA[3]\, 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        \CoreAPB3_0_APBmslave0_PWDATA[2]\, 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        \CoreAPB3_0_APBmslave0_PWDATA[1]\, 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        \CoreAPB3_0_APBmslave0_PWDATA[0]\, MAC_MII_TXD_c(3) => 
        \MAC_MII_TXD_c[3]\, MAC_MII_TXD_c(2) => 
        \MAC_MII_TXD_c[2]\, MAC_MII_TXD_c(1) => 
        \MAC_MII_TXD_c[1]\, MAC_MII_TXD_c(0) => 
        \MAC_MII_TXD_c[0]\, CoreAPB3_0_APBmslave0_PRDATA_m(7) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[7]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(6) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[6]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(5) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[5]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(4) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[4]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(3) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[3]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(2) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[2]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(1) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[1]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(0) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[0]\, Y_net_0(3) => 
        \Y_net_0[3]\, Y_net_0(2) => \Y_net_0[2]\, Y_net_0(1) => 
        \Y_net_0[1]\, Y_net_0(0) => \Y_net_0[0]\, 
        MAC_MII_RXD_c(3) => \MAC_MII_RXD_c[3]\, MAC_MII_RXD_c(2)
         => \MAC_MII_RXD_c[2]\, MAC_MII_RXD_c(1) => 
        \MAC_MII_RXD_c[1]\, MAC_MII_RXD_c(0) => 
        \MAC_MII_RXD_c[0]\, SPI_1_SS0_OTH_0 => SPI_1_SS0_OTH(0), 
        DEBOUNCE_OUT_net_0_0 => \DEBOUNCE_OUT_net_0[0]\, 
        GPIO_7_PADI_0 => GPIO_7_PADI(0), GPIO_6_PAD_0 => 
        GPIO_6_PAD(0), GPIO_1_BI_0 => GPIO_1_BI(0), 
        SPI_1_SS0_CAM_0 => SPI_1_SS0_CAM(0), SPI_1_CLK_0 => 
        SPI_1_CLK(0), SPI_0_SS1 => SPI_0_SS1, SPI_0_SS0 => 
        SPI_0_SS0, SPI_0_DO => SPI_0_DO, SPI_0_DI => SPI_0_DI, 
        SPI_0_CLK => SPI_0_CLK, MMUART_1_TXD => MMUART_1_TXD, 
        MMUART_1_RXD => MMUART_1_RXD, MDDR_WE_N => MDDR_WE_N, 
        MDDR_RESET_N => MDDR_RESET_N, MDDR_RAS_N => MDDR_RAS_N, 
        MDDR_ODT => MDDR_ODT, MDDR_DQS_TMATCH_0_OUT => 
        MDDR_DQS_TMATCH_0_OUT, MDDR_DQS_TMATCH_0_IN => 
        MDDR_DQS_TMATCH_0_IN, MDDR_CS_N => MDDR_CS_N, MDDR_CKE
         => MDDR_CKE, MDDR_CAS_N => MDDR_CAS_N, I2C_1_SDA => 
        I2C_1_SDA, I2C_1_SCL => I2C_1_SCL, GPIO_31_BI => 
        GPIO_31_BI, GPIO_26_BI => GPIO_26_BI, GPIO_25_BI => 
        GPIO_25_BI, GPIO_20_OUT => GPIO_20_OUT, GPIO_18_BI => 
        GPIO_18_BI, GPIO_17_BI => GPIO_17_BI, GPIO_16_BI => 
        GPIO_16_BI, GPIO_15_BI => GPIO_15_BI, GPIO_14_BI => 
        GPIO_14_BI, GPIO_12_BI => GPIO_12_BI, GPIO_4_BI => 
        GPIO_4_BI, GPIO_3_BI => GPIO_3_BI, GPIO_0_BI => GPIO_0_BI, 
        CoreAPB3_0_APBmslave0_PENABLE => 
        CoreAPB3_0_APBmslave0_PENABLE, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx, 
        CoreAPB3_0_APBmslave0_PWRITE => 
        CoreAPB3_0_APBmslave0_PWRITE, MAC_MII_MDC_c => 
        MAC_MII_MDC_c, GPIO_22_M2F_c => GPIO_22_M2F_c, 
        GPIO_21_M2F_c => GPIO_21_M2F_c, 
        m2s010_som_sb_0_GPIO_28_SW_RESET => 
        m2s010_som_sb_0_GPIO_28_SW_RESET, MMUART_0_TXD_M2F_c => 
        MMUART_0_TXD_M2F_c, GPIO_24_M2F_c => GPIO_24_M2F_c, 
        GPIO_5_M2F_c => GPIO_5_M2F_c, GPIO_8_M2F_c => 
        GPIO_8_M2F_c, GPIO_11_M2F_c => GPIO_11_M2F_c, 
        MAC_MII_TX_EN_c => MAC_MII_TX_EN_c, MAC_MII_COL_c => 
        MAC_MII_COL_c, MAC_MII_CRS_c => MAC_MII_CRS_c, 
        CommsFPGA_top_0_INT => CommsFPGA_top_0_INT, 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i => 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i, DEBOUNCE_OUT_1_c => 
        DEBOUNCE_OUT_1_c, DEBOUNCE_OUT_2_c => DEBOUNCE_OUT_2_c, 
        MMUART_0_RXD_F2M_c => MMUART_0_RXD_F2M_c, 
        MAC_MII_RX_CLK_c => MAC_MII_RX_CLK_c, MAC_MII_RX_DV_c => 
        MAC_MII_RX_DV_c, MAC_MII_RX_ER_c => MAC_MII_RX_ER_c, 
        MAC_MII_TX_CLK_c => MAC_MII_TX_CLK_c, MDDR_CLK_N => 
        MDDR_CLK_N, MDDR_CLK => MDDR_CLK, XTL => XTL, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz, 
        m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC => 
        m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC, SPI_1_DI_CAM_c
         => SPI_1_DI_CAM_c, SPI_1_DI_OTH_c => SPI_1_DI_OTH_c, 
        CommsFPGA_top_0_CAMERA_NODE => 
        CommsFPGA_top_0_CAMERA_NODE, DEVRST_N => DEVRST_N, 
        m2s010_som_sb_0_POWER_ON_RESET_N => 
        m2s010_som_sb_0_POWER_ON_RESET_N, MAC_MII_MDIO => 
        MAC_MII_MDIO, SPI_1_DO_CAM_c => SPI_1_DO_CAM_c, 
        SPI_1_DO_OTH => SPI_1_DO_OTH);
    
    GPIO_24_M2F_obuf : OUTBUF
      port map(D => GPIO_24_M2F_c, PAD => GPIO_24_M2F);
    
    \DEBOUNCE_IN_ibuf[2]\ : INBUF
      port map(PAD => DEBOUNCE_IN(2), Y => \DEBOUNCE_IN_c[2]\);
    
    \MAC_MII_RXD_ibuf[2]\ : INBUF
      port map(PAD => MAC_MII_RXD(2), Y => \MAC_MII_RXD_c[2]\);
    
    PULLDOWN_R9_ibuf : INBUF
      port map(PAD => PULLDOWN_R9, Y => Data_FAIL_c);
    
    GPIO_11_M2F_obuf : OUTBUF
      port map(D => GPIO_11_M2F_c, PAD => GPIO_11_M2F);
    
    GPIO_8_M2F_obuf : OUTBUF
      port map(D => GPIO_8_M2F_c, PAD => GPIO_8_M2F);
    
    \MAC_MII_TXD_obuf[2]\ : OUTBUF
      port map(D => \MAC_MII_TXD_c[2]\, PAD => MAC_MII_TXD(2));
    
    MAC_MII_RX_ER_ibuf : INBUF
      port map(PAD => MAC_MII_RX_ER, Y => MAC_MII_RX_ER_c);
    
    \DEBOUNCE_IN_ibuf[0]\ : INBUF
      port map(PAD => DEBOUNCE_IN(0), Y => \DEBOUNCE_IN_c[0]\);
    
    GPIO_5_M2F_obuf : OUTBUF
      port map(D => GPIO_5_M2F_c, PAD => GPIO_5_M2F);
    
    CommsFPGA_top_0 : CommsFPGA_top
      port map(CoreAPB3_0_APBmslave0_PWDATA(7) => 
        \CoreAPB3_0_APBmslave0_PWDATA[7]\, 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        \CoreAPB3_0_APBmslave0_PWDATA[6]\, 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        \CoreAPB3_0_APBmslave0_PWDATA[5]\, 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        \CoreAPB3_0_APBmslave0_PWDATA[4]\, 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        \CoreAPB3_0_APBmslave0_PWDATA[3]\, 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        \CoreAPB3_0_APBmslave0_PWDATA[2]\, 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        \CoreAPB3_0_APBmslave0_PWDATA[1]\, 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        \CoreAPB3_0_APBmslave0_PWDATA[0]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(7) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[7]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(6) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[6]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(5) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[5]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(4) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[4]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(3) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[3]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(2) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[2]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(1) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[1]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(0) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[0]\, 
        CoreAPB3_0_APBmslave0_PADDR(7) => 
        \CoreAPB3_0_APBmslave0_PADDR[7]\, 
        CoreAPB3_0_APBmslave0_PADDR(6) => 
        \CoreAPB3_0_APBmslave0_PADDR[6]\, 
        CoreAPB3_0_APBmslave0_PADDR(5) => 
        \CoreAPB3_0_APBmslave0_PADDR[5]\, 
        CoreAPB3_0_APBmslave0_PADDR(4) => 
        \CoreAPB3_0_APBmslave0_PADDR[4]\, 
        CoreAPB3_0_APBmslave0_PADDR(3) => 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, 
        CoreAPB3_0_APBmslave0_PADDR(1) => 
        \CoreAPB3_0_APBmslave0_PADDR[1]\, 
        CoreAPB3_0_APBmslave0_PADDR(0) => 
        \CoreAPB3_0_APBmslave0_PADDR[0]\, DEBOUNCE_IN_c(2) => 
        \DEBOUNCE_IN_c[2]\, DEBOUNCE_IN_c(1) => 
        \DEBOUNCE_IN_c[1]\, DEBOUNCE_IN_c(0) => 
        \DEBOUNCE_IN_c[0]\, Y_net_0(3) => \Y_net_0[3]\, 
        Y_net_0(2) => \Y_net_0[2]\, Y_net_0(1) => \Y_net_0[1]\, 
        DEBOUNCE_OUT_net_0_0 => \DEBOUNCE_OUT_net_0[0]\, 
        MANCHESTER_IN_c => MANCHESTER_IN_c, MANCH_OUT_P_c => 
        MANCH_OUT_P_c, MANCH_OUT_P_c_i => MANCH_OUT_P_c_i, 
        DRVR_EN_c => DRVR_EN_c, N_855_i_i => 
        \CommsFPGA_top_0.N_855_i_i\, CoreAPB3_0_APBmslave0_PSELx
         => CoreAPB3_0_APBmslave0_PSELx, 
        CoreAPB3_0_APBmslave0_PENABLE => 
        CoreAPB3_0_APBmslave0_PENABLE, 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i => 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i, 
        CoreAPB3_0_APBmslave0_PWRITE => 
        CoreAPB3_0_APBmslave0_PWRITE, N_855_i => N_855_i, 
        CommsFPGA_top_0_INT => CommsFPGA_top_0_INT, 
        DEBOUNCE_OUT_1_c => DEBOUNCE_OUT_1_c, DEBOUNCE_OUT_2_c
         => DEBOUNCE_OUT_2_c, CommsFPGA_top_0_CAMERA_NODE => 
        CommsFPGA_top_0_CAMERA_NODE, 
        m2s010_som_sb_0_POWER_ON_RESET_N => 
        m2s010_som_sb_0_POWER_ON_RESET_N, 
        m2s010_som_sb_0_GPIO_28_SW_RESET => 
        m2s010_som_sb_0_GPIO_28_SW_RESET, CommsFPGA_CCC_0_LOCK
         => CommsFPGA_CCC_0_LOCK, CommsFPGA_CCC_0_GL1 => 
        CommsFPGA_CCC_0_GL1, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz);
    

end DEF_ARCH; 
