-- Version: v11.8 11.8.0.26

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b19_nczQ_DYg_YFaRM_oUoP_28s_1s_x_0 is

    port( b8_FZFFLXYE      : in    std_logic_vector(11 downto 0);
          b12_PSyi_KyDbLbb : in    std_logic_vector(11 downto 0);
          IICE_comm2iice_5 : in    std_logic;
          IICE_comm2iice_3 : in    std_logic;
          IICE_comm2iice_0 : in    std_logic;
          IICE_comm2iice_4 : in    std_logic;
          b7_yYh03wy5      : in    std_logic;
          b8_jAA_KlCO      : in    std_logic;
          ttdo             : out   std_logic
        );

end b19_nczQ_DYg_YFaRM_oUoP_28s_1s_x_0;

architecture DEF_ARCH of b19_nczQ_DYg_YFaRM_oUoP_28s_1s_x_0 is 

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \b13_PLF_2grFt_FH9[22]\, VCC_net_1, 
        \b13_PLF_2grFt_FH9_10[22]\, N_27, GND_net_1, 
        \b13_PLF_2grFt_FH9[23]\, \b13_PLF_2grFt_FH9_10[23]\, 
        \b13_PLF_2grFt_FH9[24]\, \b13_PLF_2grFt_FH9_10[24]\, 
        \b13_PLF_2grFt_FH9[25]\, \b13_PLF_2grFt_FH9_10[25]\, 
        \b13_PLF_2grFt_FH9[26]\, \b13_PLF_2grFt_FH9_10[26]\, 
        \b13_PLF_2grFt_FH9[27]\, \b13_PLF_2grFt_FH9_10[27]\, 
        \b13_PLF_2grFt_FH9[7]\, \b13_PLF_2grFt_FH9_10[7]\, 
        \b13_PLF_2grFt_FH9[8]\, \b13_PLF_2grFt_FH9_10[8]\, 
        \b13_PLF_2grFt_FH9[9]\, \b13_PLF_2grFt_FH9_10[9]\, 
        \b13_PLF_2grFt_FH9[10]\, \b13_PLF_2grFt_FH9_10[10]\, 
        \b13_PLF_2grFt_FH9[11]\, \b13_PLF_2grFt_FH9_10[11]\, 
        \b13_PLF_2grFt_FH9[12]\, \b13_PLF_2grFt_FH9_10[12]\, 
        \b13_PLF_2grFt_FH9[13]\, \b13_PLF_2grFt_FH9_10[13]\, 
        \b13_PLF_2grFt_FH9[14]\, \b13_PLF_2grFt_FH9_10[14]\, 
        \b13_PLF_2grFt_FH9[15]\, \b13_PLF_2grFt_FH9_10[15]\, 
        \b13_PLF_2grFt_FH9[16]\, \b13_PLF_2grFt_FH9_10[16]\, 
        \b13_PLF_2grFt_FH9[17]\, \b13_PLF_2grFt_FH9_10[17]\, 
        \b13_PLF_2grFt_FH9[18]\, \b13_PLF_2grFt_FH9_10[18]\, 
        \b13_PLF_2grFt_FH9[19]\, \b13_PLF_2grFt_FH9_10[19]\, 
        \b13_PLF_2grFt_FH9[20]\, \b13_PLF_2grFt_FH9_10[20]\, 
        \b13_PLF_2grFt_FH9[21]\, \b13_PLF_2grFt_FH9_10[21]\, 
        \b13_PLF_2grFt_FH9_10[0]\, \b13_PLF_2grFt_FH9[1]\, 
        \b13_PLF_2grFt_FH9_10[1]\, \b13_PLF_2grFt_FH9[2]\, 
        \b13_PLF_2grFt_FH9_10[2]\, \b13_PLF_2grFt_FH9[3]\, 
        \b13_PLF_2grFt_FH9_10[3]\, \b13_PLF_2grFt_FH9[4]\, 
        \b13_PLF_2grFt_FH9_10[4]\, \b13_PLF_2grFt_FH9[5]\, 
        \b13_PLF_2grFt_FH9_10[5]\, \b13_PLF_2grFt_FH9[6]\, 
        \b13_PLF_2grFt_FH9_10[6]\ : std_logic;

begin 


    \genblk1.b13_PLF_2grFt_FH9_10[25]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => b12_PSyi_KyDbLbb(9), B => 
        \b13_PLF_2grFt_FH9[26]\, C => IICE_comm2iice_3, Y => 
        \b13_PLF_2grFt_FH9_10[25]\);
    
    \genblk1.b13_PLF_2grFt_FH9_10[0]\ : CFG2
      generic map(INIT => x"4")

      port map(A => IICE_comm2iice_3, B => \b13_PLF_2grFt_FH9[1]\, 
        Y => \b13_PLF_2grFt_FH9_10[0]\);
    
    \genblk1.b13_PLF_2grFt_FH9_10[19]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => b12_PSyi_KyDbLbb(3), B => 
        \b13_PLF_2grFt_FH9[20]\, C => IICE_comm2iice_3, Y => 
        \b13_PLF_2grFt_FH9_10[19]\);
    
    \genblk1.b13_PLF_2grFt_FH9[2]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_10[2]\, CLK => 
        IICE_comm2iice_5, EN => N_27, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[2]\);
    
    \genblk1.b13_PLF_2grFt_FH9_10[22]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => b12_PSyi_KyDbLbb(6), B => 
        \b13_PLF_2grFt_FH9[23]\, C => IICE_comm2iice_3, Y => 
        \b13_PLF_2grFt_FH9_10[22]\);
    
    \genblk1.b13_PLF_2grFt_FH9_10[15]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => b8_FZFFLXYE(11), B => \b13_PLF_2grFt_FH9[16]\, 
        C => IICE_comm2iice_3, Y => \b13_PLF_2grFt_FH9_10[15]\);
    
    \genblk1.b13_PLF_2grFt_FH9_10[2]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => b8_jAA_KlCO, B => \b13_PLF_2grFt_FH9[3]\, C
         => IICE_comm2iice_3, Y => \b13_PLF_2grFt_FH9_10[2]\);
    
    \genblk1.b13_PLF_2grFt_FH9[5]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_10[5]\, CLK => 
        IICE_comm2iice_5, EN => N_27, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[5]\);
    
    \genblk1.b13_PLF_2grFt_FH9_10[5]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => b8_FZFFLXYE(1), B => \b13_PLF_2grFt_FH9[6]\, 
        C => IICE_comm2iice_3, Y => \b13_PLF_2grFt_FH9_10[5]\);
    
    \genblk1.b13_PLF_2grFt_FH9[16]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_10[16]\, CLK => 
        IICE_comm2iice_5, EN => N_27, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[16]\);
    
    \genblk1.b13_PLF_2grFt_FH9_10[1]\ : CFG2
      generic map(INIT => x"4")

      port map(A => IICE_comm2iice_3, B => \b13_PLF_2grFt_FH9[2]\, 
        Y => \b13_PLF_2grFt_FH9_10[1]\);
    
    \genblk1.b13_PLF_2grFt_FH9_10[3]\ : CFG2
      generic map(INIT => x"4")

      port map(A => IICE_comm2iice_3, B => \b13_PLF_2grFt_FH9[4]\, 
        Y => \b13_PLF_2grFt_FH9_10[3]\);
    
    \genblk1.b13_PLF_2grFt_FH9[10]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_10[10]\, CLK => 
        IICE_comm2iice_5, EN => N_27, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[10]\);
    
    \genblk1.b13_PLF_2grFt_FH9_10[12]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => b8_FZFFLXYE(8), B => \b13_PLF_2grFt_FH9[13]\, 
        C => IICE_comm2iice_3, Y => \b13_PLF_2grFt_FH9_10[12]\);
    
    \genblk1.b13_PLF_2grFt_FH9[23]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_10[23]\, CLK => 
        IICE_comm2iice_5, EN => N_27, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[23]\);
    
    \genblk1.b13_PLF_2grFt_FH9[0]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_10[0]\, CLK => 
        IICE_comm2iice_5, EN => N_27, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => ttdo);
    
    \genblk1.b13_PLF_2grFt_FH9_10[6]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => b8_FZFFLXYE(2), B => \b13_PLF_2grFt_FH9[7]\, 
        C => IICE_comm2iice_3, Y => \b13_PLF_2grFt_FH9_10[6]\);
    
    \genblk1.b13_PLF_2grFt_FH9[11]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_10[11]\, CLK => 
        IICE_comm2iice_5, EN => N_27, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[11]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \genblk1.b13_PLF_2grFt_FH9_10[9]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => b8_FZFFLXYE(5), B => \b13_PLF_2grFt_FH9[10]\, 
        C => IICE_comm2iice_3, Y => \b13_PLF_2grFt_FH9_10[9]\);
    
    \genblk1.b13_PLF_2grFt_FH9[12]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_10[12]\, CLK => 
        IICE_comm2iice_5, EN => N_27, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[12]\);
    
    \genblk1.b13_PLF_2grFt_FH9[17]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_10[17]\, CLK => 
        IICE_comm2iice_5, EN => N_27, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[17]\);
    
    \genblk1.b13_PLF_2grFt_FH9[26]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_10[26]\, CLK => 
        IICE_comm2iice_5, EN => N_27, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[26]\);
    
    \genblk1.b13_PLF_2grFt_FH9[20]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_10[20]\, CLK => 
        IICE_comm2iice_5, EN => N_27, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[20]\);
    
    \genblk1.b13_PLF_2grFt_FH9_10[27]\ : CFG2
      generic map(INIT => x"8")

      port map(A => IICE_comm2iice_3, B => b12_PSyi_KyDbLbb(11), 
        Y => \b13_PLF_2grFt_FH9_10[27]\);
    
    \genblk1.b13_PLF_2grFt_FH9[14]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_10[14]\, CLK => 
        IICE_comm2iice_5, EN => N_27, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[14]\);
    
    \genblk1.b13_PLF_2grFt_FH9[6]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_10[6]\, CLK => 
        IICE_comm2iice_5, EN => N_27, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[6]\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \genblk1.b13_PLF_2grFt_FH9[21]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_10[21]\, CLK => 
        IICE_comm2iice_5, EN => N_27, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[21]\);
    
    \genblk1.b13_PLF_2grFt_FH9_10[17]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => b12_PSyi_KyDbLbb(1), B => 
        \b13_PLF_2grFt_FH9[18]\, C => IICE_comm2iice_3, Y => 
        \b13_PLF_2grFt_FH9_10[17]\);
    
    \genblk1.b13_PLF_2grFt_FH9_10[20]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => b12_PSyi_KyDbLbb(4), B => 
        \b13_PLF_2grFt_FH9[21]\, C => IICE_comm2iice_3, Y => 
        \b13_PLF_2grFt_FH9_10[20]\);
    
    \genblk1.b13_PLF_2grFt_FH9[22]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_10[22]\, CLK => 
        IICE_comm2iice_5, EN => N_27, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[22]\);
    
    \genblk1.b13_PLF_2grFt_FH9[18]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_10[18]\, CLK => 
        IICE_comm2iice_5, EN => N_27, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[18]\);
    
    \genblk1.b13_PLF_2grFt_FH9_10[21]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => b12_PSyi_KyDbLbb(5), B => 
        \b13_PLF_2grFt_FH9[22]\, C => IICE_comm2iice_3, Y => 
        \b13_PLF_2grFt_FH9_10[21]\);
    
    \genblk1.b13_PLF_2grFt_FH9_10[23]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => b12_PSyi_KyDbLbb(7), B => 
        \b13_PLF_2grFt_FH9[24]\, C => IICE_comm2iice_3, Y => 
        \b13_PLF_2grFt_FH9_10[23]\);
    
    \genblk1.b13_PLF_2grFt_FH9[9]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_10[9]\, CLK => 
        IICE_comm2iice_5, EN => N_27, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[9]\);
    
    \genblk1.b13_PLF_2grFt_FH9[4]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_10[4]\, CLK => 
        IICE_comm2iice_5, EN => N_27, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[4]\);
    
    un1_b13_PLF_2grFt_FH923_i_a2 : CFG4
      generic map(INIT => x"A080")

      port map(A => IICE_comm2iice_0, B => IICE_comm2iice_3, C
         => b7_yYh03wy5, D => IICE_comm2iice_4, Y => N_27);
    
    \genblk1.b13_PLF_2grFt_FH9[27]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_10[27]\, CLK => 
        IICE_comm2iice_5, EN => N_27, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[27]\);
    
    \genblk1.b13_PLF_2grFt_FH9_10[24]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => b12_PSyi_KyDbLbb(8), B => 
        \b13_PLF_2grFt_FH9[25]\, C => IICE_comm2iice_3, Y => 
        \b13_PLF_2grFt_FH9_10[24]\);
    
    \genblk1.b13_PLF_2grFt_FH9_10[10]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => b8_FZFFLXYE(6), B => \b13_PLF_2grFt_FH9[11]\, 
        C => IICE_comm2iice_3, Y => \b13_PLF_2grFt_FH9_10[10]\);
    
    \genblk1.b13_PLF_2grFt_FH9_10[11]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => b8_FZFFLXYE(7), B => \b13_PLF_2grFt_FH9[12]\, 
        C => IICE_comm2iice_3, Y => \b13_PLF_2grFt_FH9_10[11]\);
    
    \genblk1.b13_PLF_2grFt_FH9_10[18]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => b12_PSyi_KyDbLbb(2), B => 
        \b13_PLF_2grFt_FH9[19]\, C => IICE_comm2iice_3, Y => 
        \b13_PLF_2grFt_FH9_10[18]\);
    
    \genblk1.b13_PLF_2grFt_FH9_10[13]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => b8_FZFFLXYE(9), B => \b13_PLF_2grFt_FH9[14]\, 
        C => IICE_comm2iice_3, Y => \b13_PLF_2grFt_FH9_10[13]\);
    
    \genblk1.b13_PLF_2grFt_FH9[24]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_10[24]\, CLK => 
        IICE_comm2iice_5, EN => N_27, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[24]\);
    
    \genblk1.b13_PLF_2grFt_FH9[15]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_10[15]\, CLK => 
        IICE_comm2iice_5, EN => N_27, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[15]\);
    
    \genblk1.b13_PLF_2grFt_FH9[3]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_10[3]\, CLK => 
        IICE_comm2iice_5, EN => N_27, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[3]\);
    
    \genblk1.b13_PLF_2grFt_FH9_10[8]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => b8_FZFFLXYE(4), B => \b13_PLF_2grFt_FH9[9]\, 
        C => IICE_comm2iice_3, Y => \b13_PLF_2grFt_FH9_10[8]\);
    
    \genblk1.b13_PLF_2grFt_FH9_10[14]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => b8_FZFFLXYE(10), B => \b13_PLF_2grFt_FH9[15]\, 
        C => IICE_comm2iice_3, Y => \b13_PLF_2grFt_FH9_10[14]\);
    
    \genblk1.b13_PLF_2grFt_FH9[1]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_10[1]\, CLK => 
        IICE_comm2iice_5, EN => N_27, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[1]\);
    
    \genblk1.b13_PLF_2grFt_FH9[7]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_10[7]\, CLK => 
        IICE_comm2iice_5, EN => N_27, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[7]\);
    
    \genblk1.b13_PLF_2grFt_FH9[19]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_10[19]\, CLK => 
        IICE_comm2iice_5, EN => N_27, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[19]\);
    
    \genblk1.b13_PLF_2grFt_FH9_10[7]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => b8_FZFFLXYE(3), B => \b13_PLF_2grFt_FH9[8]\, 
        C => IICE_comm2iice_3, Y => \b13_PLF_2grFt_FH9_10[7]\);
    
    \genblk1.b13_PLF_2grFt_FH9[8]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_10[8]\, CLK => 
        IICE_comm2iice_5, EN => N_27, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[8]\);
    
    \genblk1.b13_PLF_2grFt_FH9_10[26]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => b12_PSyi_KyDbLbb(10), B => 
        \b13_PLF_2grFt_FH9[27]\, C => IICE_comm2iice_3, Y => 
        \b13_PLF_2grFt_FH9_10[26]\);
    
    \genblk1.b13_PLF_2grFt_FH9[25]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_10[25]\, CLK => 
        IICE_comm2iice_5, EN => N_27, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[25]\);
    
    \genblk1.b13_PLF_2grFt_FH9_10[16]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => b12_PSyi_KyDbLbb(0), B => 
        \b13_PLF_2grFt_FH9[17]\, C => IICE_comm2iice_3, Y => 
        \b13_PLF_2grFt_FH9_10[16]\);
    
    \genblk1.b13_PLF_2grFt_FH9_10[4]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => b8_FZFFLXYE(0), B => \b13_PLF_2grFt_FH9[5]\, 
        C => IICE_comm2iice_3, Y => \b13_PLF_2grFt_FH9_10[4]\);
    
    \genblk1.b13_PLF_2grFt_FH9[13]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_10[13]\, CLK => 
        IICE_comm2iice_5, EN => N_27, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[13]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b13_vFW_xNywD_EdR_174s_12s_4096s_0s_x_0 is

    port( b11_OFWNT9L_8tZ     : in    std_logic_vector(167 downto 0);
          b7_vFW_PlM          : out   std_logic_vector(167 downto 0);
          b12_2_St6KCa_jHv    : in    std_logic_vector(11 downto 0);
          b9_v_mzCDYXs        : in    std_logic_vector(11 downto 0);
          IICE_comm2iice_0    : in    std_logic;
          b4_2o_z             : in    std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic
        );

end b13_vFW_xNywD_EdR_174s_12s_4096s_0s_x_0;

architecture DEF_ARCH of b13_vFW_xNywD_EdR_174s_12s_4096s_0s_x_0 is 

  component RAM1K18
    generic (MEMORYFILE:string := "");

    port( A_DOUT        : out   std_logic_vector(17 downto 0);
          B_DOUT        : out   std_logic_vector(17 downto 0);
          BUSY          : out   std_logic;
          A_CLK         : in    std_logic := 'U';
          A_DOUT_CLK    : in    std_logic := 'U';
          A_ARST_N      : in    std_logic := 'U';
          A_DOUT_EN     : in    std_logic := 'U';
          A_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_DOUT_ARST_N : in    std_logic := 'U';
          A_DOUT_SRST_N : in    std_logic := 'U';
          A_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          A_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          A_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          B_CLK         : in    std_logic := 'U';
          B_DOUT_CLK    : in    std_logic := 'U';
          B_ARST_N      : in    std_logic := 'U';
          B_DOUT_EN     : in    std_logic := 'U';
          B_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_DOUT_ARST_N : in    std_logic := 'U';
          B_DOUT_SRST_N : in    std_logic := 'U';
          B_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          B_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          B_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          A_EN          : in    std_logic := 'U';
          A_DOUT_LAT    : in    std_logic := 'U';
          A_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_WMODE       : in    std_logic := 'U';
          B_EN          : in    std_logic := 'U';
          B_DOUT_LAT    : in    std_logic := 'U';
          B_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_WMODE       : in    std_logic := 'U';
          SII_LOCK      : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;
    signal nc1168, nc783, nc488, nc74, nc54, nc302, nc406, nc1104, 
        nc312, nc416, nc461, nc860, nc599, nc309, nc1316, nc863, 
        nc1307, nc753, nc458, nc1339, nc845, nc32, nc1195, nc1088, 
        nc745, nc402, nc978, nc319, nc907, nc228, nc325, nc934, 
        nc8, nc1101, nc148, nc327, nc1228, nc1061, nc346, nc412, 
        nc917, nc98, nc771, nc867, nc60, nc737, nc196, nc224, 
        nc649, nc29, nc898, nc601, nc993, nc677, nc769, nc102, 
        nc120, nc61, nc1082, nc611, nc525, nc1084, nc1006, nc95, 
        nc1188, nc328, nc273, nc946, nc374, nc580, nc112, nc792, 
        nc921, nc866, nc1226, nc10, nc42, nc341, nc602, nc79, 
        nc231, nc135, nc59, nc920, nc869, nc1311, nc1249, nc11, 
        nc734, nc444, nc330, nc550, nc612, nc562, nc427, nc1300, 
        nc1238, nc579, nc1081, nc895, nc588, nc795, nc86, nc1193, 
        nc604, nc460, nc1112, nc1172, nc198, nc322, nc426, nc1069, 
        nc441, nc840, nc280, nc1093, nc396, nc103, nc1124, nc614, 
        nc843, nc1015, nc1075, nc1290, nc1146, nc586, nc329, 
        nc699, nc558, nc113, nc1155, nc176, nc33, nc1327, nc27, 
        nc878, nc973, nc238, nc335, nc1291, nc1236, nc383, nc485, 
        nc422, nc927, nc250, nc683, nc1121, nc1010, nc337, nc1149, 
        nc1070, nc703, nc408, nc847, nc567, nc996, nc1295, nc556, 
        nc772, nc234, nc1197, nc713, nc418, nc749, nc884, nc391, 
        nc62, nc1190, nc353, nc455, nc621, nc788, nc130, nc653, 
        nc77, nc57, nc535, nc760, nc122, nc494, nc583, nc846, 
        nc338, nc1242, nc1026, nc931, nc1089, nc854, nc1134, 
        nc1097, nc849, nc90, nc169, nc1343, nc43, nc758, nc1305, 
        nc12, nc930, nc875, nc766, nc775, nc622, nc542, nc1293, 
        nc685, nc553, nc1337, nc491, nc91, nc890, nc178, nc893, 
        nc581, nc376, nc437, nc1131, nc84, nc1297, nc440, nc1320, 
        nc500, nc679, nc1153, nc1105, nc1294, nc655, nc624, nc332, 
        nc436, nc1053, nc510, nc184, nc897, nc551, nc483, nc1250, 
        nc688, nc123, nc976, nc339, nc799, nc1036, nc584, nc964, 
        nc286, nc1251, nc371, nc432, nc287, nc937, nc547, nc154, 
        nc508, nc896, nc453, nc686, nc658, nc474, nc767, nc723, 
        nc428, nc1255, nc1308, nc1162, nc554, nc200, nc1157, 
        nc256, nc518, nc899, nc3, nc1219, nc680, nc489, nc63, 
        nc1279, nc1150, nc631, nc257, nc740, nc1065, nc1330, 
        nc506, nc210, nc592, nc132, nc656, nc1098, nc471, nc870, 
        nc303, nc405, nc516, nc873, nc149, nc603, nc1057, nc650, 
        nc89, nc459, nc490, nc261, nc165, nc746, nc1060, nc313, 
        nc415, nc13, nc881, nc92, nc1103, nc764, nc613, nc360, 
        nc632, nc1325, nc1253, nc804, nc285, nc1116, nc1302, 
        nc1176, nc1003, nc708, nc877, nc1200, nc1092, nc814, 
        nc1257, nc1094, nc503, nc4, nc1198, nc718, nc851, nc779, 
        nc1119, nc1254, nc1179, nc520, nc1182, nc1201, nc255, 
        nc1125, nc513, nc634, nc597, nc282, nc1085, nc876, nc133, 
        nc605, nc1205, nc944, nc36, nc1107, nc365, nc268, nc982, 
        nc501, nc1100, nc879, nc1248, nc790, nc615, nc367, nc1212, 
        nc1272, nc252, nc1091, nc747, nc1080, nc882, nc572, nc511, 
        nc1335, nc528, nc733, nc438, nc1313, nc264, nc199, nc104, 
        nc1328, nc1007, nc952, nc796, nc160, nc220, nc403, nc87, 
        nc608, nc470, nc565, nc114, nc368, nc852, nc504, nc1203, 
        nc206, nc526, nc413, nc1058, nc618, nc1246, nc961, nc1135, 
        nc985, nc207, nc241, nc145, nc514, nc323, nc425, nc216, 
        nc46, nc6, nc1207, nc989, nc606, nc960, nc623, nc744, 
        nc340, nc217, nc181, nc93, nc187, nc1204, nc1123, nc616, 
        nc600, nc409, nc289, nc577, nc467, nc955, nc824, nc1269, 
        nc1322, nc1023, nc728, nc1052, nc994, nc610, nc419, 
        nc1054, nc959, nc1220, nc1158, nc151, nc523, nc1, nc157, 
        nc362, nc466, nc530, nc1338, nc1144, nc1099, nc770, nc259, 
        nc1221, nc797, nc801, nc34, nc369, nc345, nc248, nc205, 
        nc988, nc625, nc179, nc1225, nc811, nc1319, nc1166, nc347, 
        nc1141, nc462, nc1127, nc967, nc776, nc215, nc521, nc1120, 
        nc1051, nc781, nc244, nc1008, nc538, nc1133, nc291, nc195, 
        nc1169, nc958, nc66, nc140, nc687, nc202, nc1332, nc661, 
        nc545, nc794, nc390, nc1289, nc1033, nc230, nc124, nc1027, 
        nc348, nc162, nc423, nc751, nc1230, nc628, nc1046, nc212, 
        nc283, nc941, nc384, nc902, nc536, nc524, nc1223, nc226, 
        nc44, nc657, nc1231, nc940, nc333, nc435, nc1002, nc227, 
        nc1262, nc912, nc802, nc1004, nc974, nc16, nc633, nc1108, 
        nc662, nc1227, nc626, nc253, nc354, nc1235, nc812, nc447, 
        nc1224, nc1186, nc1137, nc834, nc620, nc429, nc1340, 
        nc1130, nc777, nc589, nc39, nc738, nc395, nc298, nc1218, 
        nc1278, nc342, nc446, nc397, nc533, nc905, nc9, nc664, 
        nc1189, nc1059, nc909, nc1037, nc1001, nc349, nc294, 
        nc915, nc559, nc163, nc101, nc107, nc821, nc919, nc186, 
        nc190, nc28, nc888, nc271, nc442, nc1233, nc983, nc175, 
        nc209, nc947, nc635, nc595, nc225, nc111, nc117, nc398, 
        nc774, nc370, nc1216, nc531, nc1276, nc1282, nc991, nc219, 
        nc1237, nc763, nc468, nc49, nc64, nc782, nc156, nc1192, 
        nc641, nc25, nc990, nc858, nc1234, nc1028, nc953, nc142, 
        nc78, nc58, nc222, nc134, nc1095, nc433, nc908, nc638, 
        nc497, nc752, nc534, nc236, nc922, nc1304, nc918, nc14, 
        nc701, nc37, nc237, nc642, nc1114, nc885, nc375, nc75, 
        nc278, nc392, nc496, nc1090, nc55, nc1174, nc96, nc785, 
        nc1022, nc822, nc1024, nc636, nc711, nc377, nc1128, nc188, 
        nc607, nc1009, nc386, nc1317, nc399, nc630, nc439, nc274, 
        nc617, nc203, nc1111, nc304, nc855, nc1171, nc689, nc492, 
        nc755, nc997, nc644, nc1145, nc170, nc560, nc1038, nc158, 
        nc213, nc575, nc314, nc925, nc356, nc378, nc143, nc971, 
        nc986, nc929, nc69, nc1021, nc691, nc659, nc831, nc121, 
        nc47, nc127, nc970, nc381, nc235, nc1016, nc192, nc509, 
        nc1076, nc229, nc743, nc448, nc484, nc1306, nc1032, 
        nc1034, nc956, nc1268, nc519, nc568, nc477, nc1138, 
        nc1152, nc19, nc351, nc260, nc692, nc232, nc372, nc476, 
        nc1055, nc106, nc454, nc20, nc808, nc566, nc1310, nc903, 
        nc481, nc880, nc928, nc883, nc116, nc363, nc465, nc932, 
        nc379, nc21, nc818, nc913, nc94, nc663, nc1266, nc1324, 
        nc1050, nc694, nc1031, nc721, nc1143, nc702, nc472, nc832, 
        nc977, nc451, nc850, nc1342, nc193, nc1043, nc864, nc853, 
        nc887, nc627, nc70, nc712, nc50, nc1299, nc1029, nc768, 
        nc1240, nc1301, nc67, nc540, nc789, nc563, nc71, nc1288, 
        nc671, nc223, nc51, nc324, nc1241, nc172, nc935, nc793, 
        nc498, nc857, nc805, nc705, nc886, nc1164, nc939, nc1245, 
        nc108, nc1102, nc815, nc759, nc665, nc131, nc1147, nc306, 
        nc137, nc715, nc889, nc17, nc1196, nc1140, nc672, nc118, 
        nc561, nc239, nc1334, nc1005, nc529, nc609, nc582, nc548, 
        nc316, nc1286, nc856, nc1161, nc1326, nc240, nc1315, 
        nc1199, nc619, nc859, nc99, nc1047, nc88, nc480, nc1039, 
        nc164, nc906, nc1000, nc463, nc546, nc674, nc668, nc552, 
        nc1243, nc301, nc916, nc564, nc126, nc266, nc343, nc445, 
        nc22, nc938, nc828, nc923, nc173, nc643, nc1066, nc1115, 
        nc267, nc85, nc1175, nc404, nc450, nc311, nc1292, nc1247, 
        nc590, nc731, nc666, nc1184, nc1244, nc844, nc414, nc722, 
        nc587, nc748, nc660, nc469, nc773, nc637, nc478, nc1259, 
        nc72, nc52, nc543, nc401, nc800, nc1181, nc1336, nc233, 
        nc803, nc1321, nc334, nc780, nc557, nc411, nc810, nc598, 
        nc1318, nc813, nc825, nc645, nc861, nc725, nc290, nc189, 
        nc265, nc128, nc807, nc541, nc1156, nc1122, nc786, nc97, 
        nc750, nc326, nc1086, nc596, nc539, nc817, nc709, nc1025, 
        nc393, nc495, nc629, nc1048, nc693, nc159, nc1159, nc144, 
        nc719, nc1113, nc1173, nc756, nc443, nc806, nc648, nc262, 
        nc1312, nc570, nc1013, nc1073, nc926, nc894, nc544, 
        nc1020, nc246, nc1331, nc816, nc809, nc1210, nc798, 
        nc1270, nc136, nc23, nc962, nc838, nc247, nc933, nc321, 
        nc1209, nc593, nc502, nc1042, nc984, nc819, nc646, nc1252, 
        nc1044, nc1211, nc1271, nc1148, nc862, nc424, nc512, 
        nc640, nc449, nc80, nc732, nc1132, nc400, nc1215, nc1275, 
        nc787, nc578, nc1117, nc695, nc1177, nc954, nc73, nc81, 
        nc1110, nc53, nc410, nc1170, nc1035, nc270, nc591, nc421, 
        nc820, nc1106, nc965, nc823, nc576, nc1165, nc757, nc1041, 
        nc969, nc841, nc1017, nc1030, nc835, nc1077, nc245, nc161, 
        nc373, nc475, nc735, nc167, nc281, nc194, nc507, nc185, 
        nc1109, nc673, nc493, nc138, nc698, nc269, nc1213, nc784, 
        nc380, nc1273, nc336, nc827, nc517, nc594, nc296, nc874, 
        nc1298, nc639, nc729, nc297, nc1217, nc778, nc700, nc251, 
        nc1277, nc155, nc242, nc696, nc1214, nc754, nc573, nc350, 
        nc1202, nc1274, nc710, nc826, nc109, nc936, nc690, nc499, 
        nc942, nc1303, nc968, nc706, nc829, nc119, nc331, nc1344, 
        nc38, nc842, nc385, nc288, nc1185, nc675, nc1229, nc1296, 
        nc761, nc716, nc522, nc434, nc387, nc571, nc1049, nc667, 
        nc1163, nc891, nc2, nc82, nc284, nc420, nc35, nc295, 
        nc355, nc258, nc1063, nc263, nc180, nc364, nc357, nc174, 
        nc945, nc585, nc1260, nc431, nc830, nc473, nc678, nc388, 
        nc904, nc833, nc1018, nc949, nc1126, nc1078, nc981, nc254, 
        nc574, nc141, nc276, nc1261, nc147, nc1194, nc914, nc48, 
        nc7, nc5, nc150, nc277, nc292, nc980, nc249, nc707, nc555, 
        nc527, nc1129, nc676, nc1265, nc358, nc837, nc569, nc1239, 
        nc1167, nc951, nc717, nc992, nc487, nc1160, nc1191, 
        nc1258, nc670, nc479, nc1012, nc45, nc1072, nc1014, nc739, 
        nc1074, nc1118, nc950, nc1309, nc1178, nc892, nc720, 
        nc1183, nc382, nc486, nc1222, nc836, nc201, nc948, nc105, 
        nc1067, nc1083, nc457, nc166, nc26, nc868, nc129, nc963, 
        nc704, nc300, nc1280, nc389, nc1323, nc839, nc211, nc1136, 
        nc115, nc1096, nc871, nc726, nc1263, nc741, nc1256, nc275, 
        nc352, nc456, nc714, nc310, nc482, nc532, nc1281, nc995, 
        nc987, nc1011, nc1071, nc762, nc647, nc1267, nc999, 
        nc1139, nc359, nc191, nc1285, nc83, nc197, nc1264, nc430, 
        nc76, nc56, nc243, nc68, nc1187, nc344, nc1341, nc681, 
        nc452, nc299, nc1180, nc957, nc272, nc182, nc30, nc305, 
        nc208, nc924, nc865, nc1232, nc307, nc31, nc1208, nc1154, 
        nc972, nc765, nc65, nc315, nc218, nc1087, nc651, nc1142, 
        nc168, nc18, nc1333, nc317, nc682, nc549, nc366, nc152, 
        nc204, nc872, nc537, nc727, nc1283, nc1045, nc998, nc100, 
        nc1314, nc669, nc214, nc1151, nc505, nc308, nc1287, nc791, 
        nc15, nc110, nc901, nc730, nc652, nc515, nc1068, nc1329, 
        nc1206, nc1040, nc684, nc1284, nc318, nc1019, nc966, nc40, 
        nc1079, nc146, nc975, nc697, nc24, nc848, nc943, nc911, 
        nc900, nc221, nc125, nc183, nc139, nc979, nc361, nc41, 
        nc1056, nc293, nc910, nc736, nc724, nc171, nc320, nc394, 
        nc177, nc407, nc654, nc464, nc742, nc279, nc1062, nc1064, 
        nc417, nc153 : std_logic;

begin 


    b3_SoW_b3_SoW_0_1 : RAM1K18
      port map(A_DOUT(17) => nc1168, A_DOUT(16) => nc783, 
        A_DOUT(15) => nc488, A_DOUT(14) => nc74, A_DOUT(13) => 
        nc54, A_DOUT(12) => nc302, A_DOUT(11) => nc406, 
        A_DOUT(10) => nc1104, A_DOUT(9) => nc312, A_DOUT(8) => 
        nc416, A_DOUT(7) => nc461, A_DOUT(6) => nc860, A_DOUT(5)
         => nc599, A_DOUT(4) => nc309, A_DOUT(3) => b7_vFW_PlM(7), 
        A_DOUT(2) => b7_vFW_PlM(6), A_DOUT(1) => b7_vFW_PlM(5), 
        A_DOUT(0) => b7_vFW_PlM(4), B_DOUT(17) => nc1316, 
        B_DOUT(16) => nc863, B_DOUT(15) => nc1307, B_DOUT(14) => 
        nc753, B_DOUT(13) => nc458, B_DOUT(12) => nc1339, 
        B_DOUT(11) => nc845, B_DOUT(10) => nc32, B_DOUT(9) => 
        nc1195, B_DOUT(8) => nc1088, B_DOUT(7) => nc745, 
        B_DOUT(6) => nc402, B_DOUT(5) => nc978, B_DOUT(4) => 
        nc319, B_DOUT(3) => nc907, B_DOUT(2) => nc228, B_DOUT(1)
         => nc325, B_DOUT(0) => nc934, BUSY => OPEN, A_CLK => 
        IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, A_ARST_N => 
        VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2) => VCC_net_1, 
        A_BLK(1) => VCC_net_1, A_BLK(0) => VCC_net_1, 
        A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => VCC_net_1, 
        A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, A_DIN(15)
         => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13) => 
        GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => GND_net_1, 
        A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, A_DIN(8)
         => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6) => 
        GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => GND_net_1, 
        A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, A_DIN(1)
         => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13) => 
        b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(7), B_DIN(2) => 
        b11_OFWNT9L_8tZ(6), B_DIN(1) => b11_OFWNT9L_8tZ(5), 
        B_DIN(0) => b11_OFWNT9L_8tZ(4), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_27 : RAM1K18
      port map(A_DOUT(17) => nc8, A_DOUT(16) => nc1101, 
        A_DOUT(15) => nc148, A_DOUT(14) => nc327, A_DOUT(13) => 
        nc1228, A_DOUT(12) => nc1061, A_DOUT(11) => nc346, 
        A_DOUT(10) => nc412, A_DOUT(9) => nc917, A_DOUT(8) => 
        nc98, A_DOUT(7) => nc771, A_DOUT(6) => nc867, A_DOUT(5)
         => nc60, A_DOUT(4) => nc737, A_DOUT(3) => 
        b7_vFW_PlM(111), A_DOUT(2) => b7_vFW_PlM(110), A_DOUT(1)
         => b7_vFW_PlM(109), A_DOUT(0) => b7_vFW_PlM(108), 
        B_DOUT(17) => nc196, B_DOUT(16) => nc224, B_DOUT(15) => 
        nc649, B_DOUT(14) => nc29, B_DOUT(13) => nc898, 
        B_DOUT(12) => nc601, B_DOUT(11) => nc993, B_DOUT(10) => 
        nc677, B_DOUT(9) => nc769, B_DOUT(8) => nc102, B_DOUT(7)
         => nc120, B_DOUT(6) => nc61, B_DOUT(5) => nc1082, 
        B_DOUT(4) => nc611, B_DOUT(3) => nc525, B_DOUT(2) => 
        nc1084, B_DOUT(1) => nc1006, B_DOUT(0) => nc95, BUSY => 
        OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(111), B_DIN(2) => 
        b11_OFWNT9L_8tZ(110), B_DIN(1) => b11_OFWNT9L_8tZ(109), 
        B_DIN(0) => b11_OFWNT9L_8tZ(108), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_11 : RAM1K18
      port map(A_DOUT(17) => nc1188, A_DOUT(16) => nc328, 
        A_DOUT(15) => nc273, A_DOUT(14) => nc946, A_DOUT(13) => 
        nc374, A_DOUT(12) => nc580, A_DOUT(11) => nc112, 
        A_DOUT(10) => nc792, A_DOUT(9) => nc921, A_DOUT(8) => 
        nc866, A_DOUT(7) => nc1226, A_DOUT(6) => nc10, A_DOUT(5)
         => nc42, A_DOUT(4) => nc341, A_DOUT(3) => b7_vFW_PlM(47), 
        A_DOUT(2) => b7_vFW_PlM(46), A_DOUT(1) => b7_vFW_PlM(45), 
        A_DOUT(0) => b7_vFW_PlM(44), B_DOUT(17) => nc602, 
        B_DOUT(16) => nc79, B_DOUT(15) => nc231, B_DOUT(14) => 
        nc135, B_DOUT(13) => nc59, B_DOUT(12) => nc920, 
        B_DOUT(11) => nc869, B_DOUT(10) => nc1311, B_DOUT(9) => 
        nc1249, B_DOUT(8) => nc11, B_DOUT(7) => nc734, B_DOUT(6)
         => nc444, B_DOUT(5) => nc330, B_DOUT(4) => nc550, 
        B_DOUT(3) => nc612, B_DOUT(2) => nc562, B_DOUT(1) => 
        nc427, B_DOUT(0) => nc1300, BUSY => OPEN, A_CLK => 
        IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, A_ARST_N => 
        VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2) => VCC_net_1, 
        A_BLK(1) => VCC_net_1, A_BLK(0) => VCC_net_1, 
        A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => VCC_net_1, 
        A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, A_DIN(15)
         => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13) => 
        GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => GND_net_1, 
        A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, A_DIN(8)
         => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6) => 
        GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => GND_net_1, 
        A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, A_DIN(1)
         => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13) => 
        b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(47), B_DIN(2) => 
        b11_OFWNT9L_8tZ(46), B_DIN(1) => b11_OFWNT9L_8tZ(45), 
        B_DIN(0) => b11_OFWNT9L_8tZ(44), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_37 : RAM1K18
      port map(A_DOUT(17) => nc1238, A_DOUT(16) => nc579, 
        A_DOUT(15) => nc1081, A_DOUT(14) => nc895, A_DOUT(13) => 
        nc588, A_DOUT(12) => nc795, A_DOUT(11) => nc86, 
        A_DOUT(10) => nc1193, A_DOUT(9) => nc604, A_DOUT(8) => 
        nc460, A_DOUT(7) => nc1112, A_DOUT(6) => nc1172, 
        A_DOUT(5) => nc198, A_DOUT(4) => nc322, A_DOUT(3) => 
        b7_vFW_PlM(151), A_DOUT(2) => b7_vFW_PlM(150), A_DOUT(1)
         => b7_vFW_PlM(149), A_DOUT(0) => b7_vFW_PlM(148), 
        B_DOUT(17) => nc426, B_DOUT(16) => nc1069, B_DOUT(15) => 
        nc441, B_DOUT(14) => nc840, B_DOUT(13) => nc280, 
        B_DOUT(12) => nc1093, B_DOUT(11) => nc396, B_DOUT(10) => 
        nc103, B_DOUT(9) => nc1124, B_DOUT(8) => nc614, B_DOUT(7)
         => nc843, B_DOUT(6) => nc1015, B_DOUT(5) => nc1075, 
        B_DOUT(4) => nc1290, B_DOUT(3) => nc1146, B_DOUT(2) => 
        nc586, B_DOUT(1) => nc329, B_DOUT(0) => nc699, BUSY => 
        OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(151), B_DIN(2) => 
        b11_OFWNT9L_8tZ(150), B_DIN(1) => b11_OFWNT9L_8tZ(149), 
        B_DIN(0) => b11_OFWNT9L_8tZ(148), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_25 : RAM1K18
      port map(A_DOUT(17) => nc558, A_DOUT(16) => nc113, 
        A_DOUT(15) => nc1155, A_DOUT(14) => nc176, A_DOUT(13) => 
        nc33, A_DOUT(12) => nc1327, A_DOUT(11) => nc27, 
        A_DOUT(10) => nc878, A_DOUT(9) => nc973, A_DOUT(8) => 
        nc238, A_DOUT(7) => nc335, A_DOUT(6) => nc1291, A_DOUT(5)
         => nc1236, A_DOUT(4) => nc383, A_DOUT(3) => 
        b7_vFW_PlM(103), A_DOUT(2) => b7_vFW_PlM(102), A_DOUT(1)
         => b7_vFW_PlM(101), A_DOUT(0) => b7_vFW_PlM(100), 
        B_DOUT(17) => nc485, B_DOUT(16) => nc422, B_DOUT(15) => 
        nc927, B_DOUT(14) => nc250, B_DOUT(13) => nc683, 
        B_DOUT(12) => nc1121, B_DOUT(11) => nc1010, B_DOUT(10)
         => nc337, B_DOUT(9) => nc1149, B_DOUT(8) => nc1070, 
        B_DOUT(7) => nc703, B_DOUT(6) => nc408, B_DOUT(5) => 
        nc847, B_DOUT(4) => nc567, B_DOUT(3) => nc996, B_DOUT(2)
         => nc1295, B_DOUT(1) => nc556, B_DOUT(0) => nc772, BUSY
         => OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => 
        VCC_net_1, A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, 
        A_BLK(2) => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0)
         => VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N
         => VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        GND_net_1, A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, 
        A_DIN(13) => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11)
         => GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => 
        GND_net_1, A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, 
        A_DIN(6) => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4)
         => GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => 
        GND_net_1, A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, 
        A_ADDR(13) => b9_v_mzCDYXs(11), A_ADDR(12) => 
        b9_v_mzCDYXs(10), A_ADDR(11) => b9_v_mzCDYXs(9), 
        A_ADDR(10) => b9_v_mzCDYXs(8), A_ADDR(9) => 
        b9_v_mzCDYXs(7), A_ADDR(8) => b9_v_mzCDYXs(6), A_ADDR(7)
         => b9_v_mzCDYXs(5), A_ADDR(6) => b9_v_mzCDYXs(4), 
        A_ADDR(5) => b9_v_mzCDYXs(3), A_ADDR(4) => 
        b9_v_mzCDYXs(2), A_ADDR(3) => b9_v_mzCDYXs(1), A_ADDR(2)
         => b9_v_mzCDYXs(0), A_ADDR(1) => GND_net_1, A_ADDR(0)
         => GND_net_1, A_WEN(1) => GND_net_1, A_WEN(0) => 
        GND_net_1, B_CLK => CommsFPGA_CCC_0_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => VCC_net_1, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        GND_net_1, B_DIN(15) => GND_net_1, B_DIN(14) => GND_net_1, 
        B_DIN(13) => GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11)
         => GND_net_1, B_DIN(10) => GND_net_1, B_DIN(9) => 
        GND_net_1, B_DIN(8) => GND_net_1, B_DIN(7) => GND_net_1, 
        B_DIN(6) => GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4)
         => GND_net_1, B_DIN(3) => b11_OFWNT9L_8tZ(103), B_DIN(2)
         => b11_OFWNT9L_8tZ(102), B_DIN(1) => 
        b11_OFWNT9L_8tZ(101), B_DIN(0) => b11_OFWNT9L_8tZ(100), 
        B_ADDR(13) => b12_2_St6KCa_jHv(11), B_ADDR(12) => 
        b12_2_St6KCa_jHv(10), B_ADDR(11) => b12_2_St6KCa_jHv(9), 
        B_ADDR(10) => b12_2_St6KCa_jHv(8), B_ADDR(9) => 
        b12_2_St6KCa_jHv(7), B_ADDR(8) => b12_2_St6KCa_jHv(6), 
        B_ADDR(7) => b12_2_St6KCa_jHv(5), B_ADDR(6) => 
        b12_2_St6KCa_jHv(4), B_ADDR(5) => b12_2_St6KCa_jHv(3), 
        B_ADDR(4) => b12_2_St6KCa_jHv(2), B_ADDR(3) => 
        b12_2_St6KCa_jHv(1), B_ADDR(2) => b12_2_St6KCa_jHv(0), 
        B_ADDR(1) => GND_net_1, B_ADDR(0) => GND_net_1, B_WEN(1)
         => GND_net_1, B_WEN(0) => b4_2o_z, A_EN => VCC_net_1, 
        A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => GND_net_1, 
        A_WIDTH(1) => VCC_net_1, A_WIDTH(0) => GND_net_1, A_WMODE
         => VCC_net_1, B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, 
        B_WIDTH(2) => GND_net_1, B_WIDTH(1) => VCC_net_1, 
        B_WIDTH(0) => GND_net_1, B_WMODE => VCC_net_1, SII_LOCK
         => GND_net_1);
    
    b3_SoW_b3_SoW_0_20 : RAM1K18
      port map(A_DOUT(17) => nc234, A_DOUT(16) => nc1197, 
        A_DOUT(15) => nc713, A_DOUT(14) => nc418, A_DOUT(13) => 
        nc749, A_DOUT(12) => nc884, A_DOUT(11) => nc391, 
        A_DOUT(10) => nc62, A_DOUT(9) => nc1190, A_DOUT(8) => 
        nc353, A_DOUT(7) => nc455, A_DOUT(6) => nc621, A_DOUT(5)
         => nc788, A_DOUT(4) => nc130, A_DOUT(3) => 
        b7_vFW_PlM(83), A_DOUT(2) => b7_vFW_PlM(82), A_DOUT(1)
         => b7_vFW_PlM(81), A_DOUT(0) => b7_vFW_PlM(80), 
        B_DOUT(17) => nc653, B_DOUT(16) => nc77, B_DOUT(15) => 
        nc57, B_DOUT(14) => nc535, B_DOUT(13) => nc760, 
        B_DOUT(12) => nc122, B_DOUT(11) => nc494, B_DOUT(10) => 
        nc583, B_DOUT(9) => nc846, B_DOUT(8) => nc338, B_DOUT(7)
         => nc1242, B_DOUT(6) => nc1026, B_DOUT(5) => nc931, 
        B_DOUT(4) => nc1089, B_DOUT(3) => nc854, B_DOUT(2) => 
        nc1134, B_DOUT(1) => nc1097, B_DOUT(0) => nc849, BUSY => 
        OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(83), B_DIN(2) => 
        b11_OFWNT9L_8tZ(82), B_DIN(1) => b11_OFWNT9L_8tZ(81), 
        B_DIN(0) => b11_OFWNT9L_8tZ(80), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_SoW_b3_SoW_0_35 : RAM1K18
      port map(A_DOUT(17) => nc90, A_DOUT(16) => nc169, 
        A_DOUT(15) => nc1343, A_DOUT(14) => nc43, A_DOUT(13) => 
        nc758, A_DOUT(12) => nc1305, A_DOUT(11) => nc12, 
        A_DOUT(10) => nc930, A_DOUT(9) => nc875, A_DOUT(8) => 
        nc766, A_DOUT(7) => nc775, A_DOUT(6) => nc622, A_DOUT(5)
         => nc542, A_DOUT(4) => nc1293, A_DOUT(3) => 
        b7_vFW_PlM(143), A_DOUT(2) => b7_vFW_PlM(142), A_DOUT(1)
         => b7_vFW_PlM(141), A_DOUT(0) => b7_vFW_PlM(140), 
        B_DOUT(17) => nc685, B_DOUT(16) => nc553, B_DOUT(15) => 
        nc1337, B_DOUT(14) => nc491, B_DOUT(13) => nc91, 
        B_DOUT(12) => nc890, B_DOUT(11) => nc178, B_DOUT(10) => 
        nc893, B_DOUT(9) => nc581, B_DOUT(8) => nc376, B_DOUT(7)
         => nc437, B_DOUT(6) => nc1131, B_DOUT(5) => nc84, 
        B_DOUT(4) => nc1297, B_DOUT(3) => nc440, B_DOUT(2) => 
        nc1320, B_DOUT(1) => nc500, B_DOUT(0) => nc679, BUSY => 
        OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(143), B_DIN(2) => 
        b11_OFWNT9L_8tZ(142), B_DIN(1) => b11_OFWNT9L_8tZ(141), 
        B_DIN(0) => b11_OFWNT9L_8tZ(140), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_30 : RAM1K18
      port map(A_DOUT(17) => nc1153, A_DOUT(16) => nc1105, 
        A_DOUT(15) => nc1294, A_DOUT(14) => nc655, A_DOUT(13) => 
        nc624, A_DOUT(12) => nc332, A_DOUT(11) => nc436, 
        A_DOUT(10) => nc1053, A_DOUT(9) => nc510, A_DOUT(8) => 
        nc184, A_DOUT(7) => nc897, A_DOUT(6) => nc551, A_DOUT(5)
         => nc483, A_DOUT(4) => nc1250, A_DOUT(3) => 
        b7_vFW_PlM(123), A_DOUT(2) => b7_vFW_PlM(122), A_DOUT(1)
         => b7_vFW_PlM(121), A_DOUT(0) => b7_vFW_PlM(120), 
        B_DOUT(17) => nc688, B_DOUT(16) => nc123, B_DOUT(15) => 
        nc976, B_DOUT(14) => nc339, B_DOUT(13) => nc799, 
        B_DOUT(12) => nc1036, B_DOUT(11) => nc584, B_DOUT(10) => 
        nc964, B_DOUT(9) => nc286, B_DOUT(8) => nc1251, B_DOUT(7)
         => nc371, B_DOUT(6) => nc432, B_DOUT(5) => nc287, 
        B_DOUT(4) => nc937, B_DOUT(3) => nc547, B_DOUT(2) => 
        nc154, B_DOUT(1) => nc508, B_DOUT(0) => nc896, BUSY => 
        OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(123), B_DIN(2) => 
        b11_OFWNT9L_8tZ(122), B_DIN(1) => b11_OFWNT9L_8tZ(121), 
        B_DIN(0) => b11_OFWNT9L_8tZ(120), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_5 : RAM1K18
      port map(A_DOUT(17) => nc453, A_DOUT(16) => nc686, 
        A_DOUT(15) => nc658, A_DOUT(14) => nc474, A_DOUT(13) => 
        nc767, A_DOUT(12) => nc723, A_DOUT(11) => nc428, 
        A_DOUT(10) => nc1255, A_DOUT(9) => nc1308, A_DOUT(8) => 
        nc1162, A_DOUT(7) => nc554, A_DOUT(6) => nc200, A_DOUT(5)
         => nc1157, A_DOUT(4) => nc256, A_DOUT(3) => 
        b7_vFW_PlM(23), A_DOUT(2) => b7_vFW_PlM(22), A_DOUT(1)
         => b7_vFW_PlM(21), A_DOUT(0) => b7_vFW_PlM(20), 
        B_DOUT(17) => nc518, B_DOUT(16) => nc899, B_DOUT(15) => 
        nc3, B_DOUT(14) => nc1219, B_DOUT(13) => nc680, 
        B_DOUT(12) => nc489, B_DOUT(11) => nc63, B_DOUT(10) => 
        nc1279, B_DOUT(9) => nc1150, B_DOUT(8) => nc631, 
        B_DOUT(7) => nc257, B_DOUT(6) => nc740, B_DOUT(5) => 
        nc1065, B_DOUT(4) => nc1330, B_DOUT(3) => nc506, 
        B_DOUT(2) => nc210, B_DOUT(1) => nc592, B_DOUT(0) => 
        nc132, BUSY => OPEN, A_CLK => IICE_comm2iice_0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => VCC_net_1, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => VCC_net_1, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => GND_net_1, A_DIN(15) => GND_net_1, 
        A_DIN(14) => GND_net_1, A_DIN(13) => GND_net_1, A_DIN(12)
         => GND_net_1, A_DIN(11) => GND_net_1, A_DIN(10) => 
        GND_net_1, A_DIN(9) => GND_net_1, A_DIN(8) => GND_net_1, 
        A_DIN(7) => GND_net_1, A_DIN(6) => GND_net_1, A_DIN(5)
         => GND_net_1, A_DIN(4) => GND_net_1, A_DIN(3) => 
        GND_net_1, A_DIN(2) => GND_net_1, A_DIN(1) => GND_net_1, 
        A_DIN(0) => GND_net_1, A_ADDR(13) => b9_v_mzCDYXs(11), 
        A_ADDR(12) => b9_v_mzCDYXs(10), A_ADDR(11) => 
        b9_v_mzCDYXs(9), A_ADDR(10) => b9_v_mzCDYXs(8), A_ADDR(9)
         => b9_v_mzCDYXs(7), A_ADDR(8) => b9_v_mzCDYXs(6), 
        A_ADDR(7) => b9_v_mzCDYXs(5), A_ADDR(6) => 
        b9_v_mzCDYXs(4), A_ADDR(5) => b9_v_mzCDYXs(3), A_ADDR(4)
         => b9_v_mzCDYXs(2), A_ADDR(3) => b9_v_mzCDYXs(1), 
        A_ADDR(2) => b9_v_mzCDYXs(0), A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => GND_net_1, A_WEN(0)
         => GND_net_1, B_CLK => CommsFPGA_CCC_0_GL0, B_DOUT_CLK
         => VCC_net_1, B_ARST_N => VCC_net_1, B_DOUT_EN => 
        VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, 
        B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, 
        B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => GND_net_1, 
        B_DIN(16) => GND_net_1, B_DIN(15) => GND_net_1, B_DIN(14)
         => GND_net_1, B_DIN(13) => GND_net_1, B_DIN(12) => 
        GND_net_1, B_DIN(11) => GND_net_1, B_DIN(10) => GND_net_1, 
        B_DIN(9) => GND_net_1, B_DIN(8) => GND_net_1, B_DIN(7)
         => GND_net_1, B_DIN(6) => GND_net_1, B_DIN(5) => 
        GND_net_1, B_DIN(4) => GND_net_1, B_DIN(3) => 
        b11_OFWNT9L_8tZ(23), B_DIN(2) => b11_OFWNT9L_8tZ(22), 
        B_DIN(1) => b11_OFWNT9L_8tZ(21), B_DIN(0) => 
        b11_OFWNT9L_8tZ(20), B_ADDR(13) => b12_2_St6KCa_jHv(11), 
        B_ADDR(12) => b12_2_St6KCa_jHv(10), B_ADDR(11) => 
        b12_2_St6KCa_jHv(9), B_ADDR(10) => b12_2_St6KCa_jHv(8), 
        B_ADDR(9) => b12_2_St6KCa_jHv(7), B_ADDR(8) => 
        b12_2_St6KCa_jHv(6), B_ADDR(7) => b12_2_St6KCa_jHv(5), 
        B_ADDR(6) => b12_2_St6KCa_jHv(4), B_ADDR(5) => 
        b12_2_St6KCa_jHv(3), B_ADDR(4) => b12_2_St6KCa_jHv(2), 
        B_ADDR(3) => b12_2_St6KCa_jHv(1), B_ADDR(2) => 
        b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, B_ADDR(0)
         => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0) => b4_2o_z, 
        A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, A_WIDTH(2)
         => GND_net_1, A_WIDTH(1) => VCC_net_1, A_WIDTH(0) => 
        GND_net_1, A_WMODE => VCC_net_1, B_EN => VCC_net_1, 
        B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => GND_net_1, 
        B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => GND_net_1, B_WMODE
         => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_29 : RAM1K18
      port map(A_DOUT(17) => nc656, A_DOUT(16) => nc1098, 
        A_DOUT(15) => nc471, A_DOUT(14) => nc870, A_DOUT(13) => 
        nc303, A_DOUT(12) => nc405, A_DOUT(11) => nc516, 
        A_DOUT(10) => nc873, A_DOUT(9) => nc149, A_DOUT(8) => 
        nc603, A_DOUT(7) => nc1057, A_DOUT(6) => nc650, A_DOUT(5)
         => nc89, A_DOUT(4) => nc459, A_DOUT(3) => 
        b7_vFW_PlM(119), A_DOUT(2) => b7_vFW_PlM(118), A_DOUT(1)
         => b7_vFW_PlM(117), A_DOUT(0) => b7_vFW_PlM(116), 
        B_DOUT(17) => nc490, B_DOUT(16) => nc261, B_DOUT(15) => 
        nc165, B_DOUT(14) => nc746, B_DOUT(13) => nc1060, 
        B_DOUT(12) => nc313, B_DOUT(11) => nc415, B_DOUT(10) => 
        nc13, B_DOUT(9) => nc881, B_DOUT(8) => nc92, B_DOUT(7)
         => nc1103, B_DOUT(6) => nc764, B_DOUT(5) => nc613, 
        B_DOUT(4) => nc360, B_DOUT(3) => nc632, B_DOUT(2) => 
        nc1325, B_DOUT(1) => nc1253, B_DOUT(0) => nc804, BUSY => 
        OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(119), B_DIN(2) => 
        b11_OFWNT9L_8tZ(118), B_DIN(1) => b11_OFWNT9L_8tZ(117), 
        B_DIN(0) => b11_OFWNT9L_8tZ(116), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_18 : RAM1K18
      port map(A_DOUT(17) => nc285, A_DOUT(16) => nc1116, 
        A_DOUT(15) => nc1302, A_DOUT(14) => nc1176, A_DOUT(13)
         => nc1003, A_DOUT(12) => nc708, A_DOUT(11) => nc877, 
        A_DOUT(10) => nc1200, A_DOUT(9) => nc1092, A_DOUT(8) => 
        nc814, A_DOUT(7) => nc1257, A_DOUT(6) => nc1094, 
        A_DOUT(5) => nc503, A_DOUT(4) => nc4, A_DOUT(3) => 
        b7_vFW_PlM(75), A_DOUT(2) => b7_vFW_PlM(74), A_DOUT(1)
         => b7_vFW_PlM(73), A_DOUT(0) => b7_vFW_PlM(72), 
        B_DOUT(17) => nc1198, B_DOUT(16) => nc718, B_DOUT(15) => 
        nc851, B_DOUT(14) => nc779, B_DOUT(13) => nc1119, 
        B_DOUT(12) => nc1254, B_DOUT(11) => nc1179, B_DOUT(10)
         => nc520, B_DOUT(9) => nc1182, B_DOUT(8) => nc1201, 
        B_DOUT(7) => nc255, B_DOUT(6) => nc1125, B_DOUT(5) => 
        nc513, B_DOUT(4) => nc634, B_DOUT(3) => nc597, B_DOUT(2)
         => nc282, B_DOUT(1) => nc1085, B_DOUT(0) => nc876, BUSY
         => OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => 
        VCC_net_1, A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, 
        A_BLK(2) => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0)
         => VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N
         => VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        GND_net_1, A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, 
        A_DIN(13) => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11)
         => GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => 
        GND_net_1, A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, 
        A_DIN(6) => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4)
         => GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => 
        GND_net_1, A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, 
        A_ADDR(13) => b9_v_mzCDYXs(11), A_ADDR(12) => 
        b9_v_mzCDYXs(10), A_ADDR(11) => b9_v_mzCDYXs(9), 
        A_ADDR(10) => b9_v_mzCDYXs(8), A_ADDR(9) => 
        b9_v_mzCDYXs(7), A_ADDR(8) => b9_v_mzCDYXs(6), A_ADDR(7)
         => b9_v_mzCDYXs(5), A_ADDR(6) => b9_v_mzCDYXs(4), 
        A_ADDR(5) => b9_v_mzCDYXs(3), A_ADDR(4) => 
        b9_v_mzCDYXs(2), A_ADDR(3) => b9_v_mzCDYXs(1), A_ADDR(2)
         => b9_v_mzCDYXs(0), A_ADDR(1) => GND_net_1, A_ADDR(0)
         => GND_net_1, A_WEN(1) => GND_net_1, A_WEN(0) => 
        GND_net_1, B_CLK => CommsFPGA_CCC_0_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => VCC_net_1, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        GND_net_1, B_DIN(15) => GND_net_1, B_DIN(14) => GND_net_1, 
        B_DIN(13) => GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11)
         => GND_net_1, B_DIN(10) => GND_net_1, B_DIN(9) => 
        GND_net_1, B_DIN(8) => GND_net_1, B_DIN(7) => GND_net_1, 
        B_DIN(6) => GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4)
         => GND_net_1, B_DIN(3) => b11_OFWNT9L_8tZ(75), B_DIN(2)
         => b11_OFWNT9L_8tZ(74), B_DIN(1) => b11_OFWNT9L_8tZ(73), 
        B_DIN(0) => b11_OFWNT9L_8tZ(72), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_26 : RAM1K18
      port map(A_DOUT(17) => nc133, A_DOUT(16) => nc605, 
        A_DOUT(15) => nc1205, A_DOUT(14) => nc944, A_DOUT(13) => 
        nc36, A_DOUT(12) => nc1107, A_DOUT(11) => nc365, 
        A_DOUT(10) => nc268, A_DOUT(9) => nc982, A_DOUT(8) => 
        nc501, A_DOUT(7) => nc1100, A_DOUT(6) => nc879, A_DOUT(5)
         => nc1248, A_DOUT(4) => nc790, A_DOUT(3) => 
        b7_vFW_PlM(107), A_DOUT(2) => b7_vFW_PlM(106), A_DOUT(1)
         => b7_vFW_PlM(105), A_DOUT(0) => b7_vFW_PlM(104), 
        B_DOUT(17) => nc615, B_DOUT(16) => nc367, B_DOUT(15) => 
        nc1212, B_DOUT(14) => nc1272, B_DOUT(13) => nc252, 
        B_DOUT(12) => nc1091, B_DOUT(11) => nc747, B_DOUT(10) => 
        nc1080, B_DOUT(9) => nc882, B_DOUT(8) => nc572, B_DOUT(7)
         => nc511, B_DOUT(6) => nc1335, B_DOUT(5) => nc528, 
        B_DOUT(4) => nc733, B_DOUT(3) => nc438, B_DOUT(2) => 
        nc1313, B_DOUT(1) => nc264, B_DOUT(0) => nc199, BUSY => 
        OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(107), B_DIN(2) => 
        b11_OFWNT9L_8tZ(106), B_DIN(1) => b11_OFWNT9L_8tZ(105), 
        B_DIN(0) => b11_OFWNT9L_8tZ(104), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_39 : RAM1K18
      port map(A_DOUT(17) => nc104, A_DOUT(16) => nc1328, 
        A_DOUT(15) => nc1007, A_DOUT(14) => nc952, A_DOUT(13) => 
        nc796, A_DOUT(12) => nc160, A_DOUT(11) => nc220, 
        A_DOUT(10) => nc403, A_DOUT(9) => nc87, A_DOUT(8) => 
        nc608, A_DOUT(7) => nc470, A_DOUT(6) => nc565, A_DOUT(5)
         => nc114, A_DOUT(4) => nc368, A_DOUT(3) => 
        b7_vFW_PlM(159), A_DOUT(2) => b7_vFW_PlM(158), A_DOUT(1)
         => b7_vFW_PlM(157), A_DOUT(0) => b7_vFW_PlM(156), 
        B_DOUT(17) => nc852, B_DOUT(16) => nc504, B_DOUT(15) => 
        nc1203, B_DOUT(14) => nc206, B_DOUT(13) => nc526, 
        B_DOUT(12) => nc413, B_DOUT(11) => nc1058, B_DOUT(10) => 
        nc618, B_DOUT(9) => nc1246, B_DOUT(8) => nc961, B_DOUT(7)
         => nc1135, B_DOUT(6) => nc985, B_DOUT(5) => nc207, 
        B_DOUT(4) => nc241, B_DOUT(3) => nc145, B_DOUT(2) => 
        nc514, B_DOUT(1) => nc323, B_DOUT(0) => nc425, BUSY => 
        OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(159), B_DIN(2) => 
        b11_OFWNT9L_8tZ(158), B_DIN(1) => b11_OFWNT9L_8tZ(157), 
        B_DIN(0) => b11_OFWNT9L_8tZ(156), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_36 : RAM1K18
      port map(A_DOUT(17) => nc216, A_DOUT(16) => nc46, 
        A_DOUT(15) => nc6, A_DOUT(14) => nc1207, A_DOUT(13) => 
        nc989, A_DOUT(12) => nc606, A_DOUT(11) => nc960, 
        A_DOUT(10) => nc623, A_DOUT(9) => nc744, A_DOUT(8) => 
        nc340, A_DOUT(7) => nc217, A_DOUT(6) => nc181, A_DOUT(5)
         => nc93, A_DOUT(4) => nc187, A_DOUT(3) => 
        b7_vFW_PlM(147), A_DOUT(2) => b7_vFW_PlM(146), A_DOUT(1)
         => b7_vFW_PlM(145), A_DOUT(0) => b7_vFW_PlM(144), 
        B_DOUT(17) => nc1204, B_DOUT(16) => nc1123, B_DOUT(15)
         => nc616, B_DOUT(14) => nc600, B_DOUT(13) => nc409, 
        B_DOUT(12) => nc289, B_DOUT(11) => nc577, B_DOUT(10) => 
        nc467, B_DOUT(9) => nc955, B_DOUT(8) => nc824, B_DOUT(7)
         => nc1269, B_DOUT(6) => nc1322, B_DOUT(5) => nc1023, 
        B_DOUT(4) => nc728, B_DOUT(3) => nc1052, B_DOUT(2) => 
        nc994, B_DOUT(1) => nc610, B_DOUT(0) => nc419, BUSY => 
        OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(147), B_DIN(2) => 
        b11_OFWNT9L_8tZ(146), B_DIN(1) => b11_OFWNT9L_8tZ(145), 
        B_DIN(0) => b11_OFWNT9L_8tZ(144), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_24 : RAM1K18
      port map(A_DOUT(17) => nc1054, A_DOUT(16) => nc959, 
        A_DOUT(15) => nc1220, A_DOUT(14) => nc1158, A_DOUT(13)
         => nc151, A_DOUT(12) => nc523, A_DOUT(11) => nc1, 
        A_DOUT(10) => nc157, A_DOUT(9) => nc362, A_DOUT(8) => 
        nc466, A_DOUT(7) => nc530, A_DOUT(6) => nc1338, A_DOUT(5)
         => nc1144, A_DOUT(4) => nc1099, A_DOUT(3) => 
        b7_vFW_PlM(99), A_DOUT(2) => b7_vFW_PlM(98), A_DOUT(1)
         => b7_vFW_PlM(97), A_DOUT(0) => b7_vFW_PlM(96), 
        B_DOUT(17) => nc770, B_DOUT(16) => nc259, B_DOUT(15) => 
        nc1221, B_DOUT(14) => nc797, B_DOUT(13) => nc801, 
        B_DOUT(12) => nc34, B_DOUT(11) => nc369, B_DOUT(10) => 
        nc345, B_DOUT(9) => nc248, B_DOUT(8) => nc205, B_DOUT(7)
         => nc988, B_DOUT(6) => nc625, B_DOUT(5) => nc179, 
        B_DOUT(4) => nc1225, B_DOUT(3) => nc811, B_DOUT(2) => 
        nc1319, B_DOUT(1) => nc1166, B_DOUT(0) => nc347, BUSY => 
        OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(99), B_DIN(2) => 
        b11_OFWNT9L_8tZ(98), B_DIN(1) => b11_OFWNT9L_8tZ(97), 
        B_DIN(0) => b11_OFWNT9L_8tZ(96), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_2 : RAM1K18
      port map(A_DOUT(17) => nc1141, A_DOUT(16) => nc462, 
        A_DOUT(15) => nc1127, A_DOUT(14) => nc967, A_DOUT(13) => 
        nc776, A_DOUT(12) => nc215, A_DOUT(11) => nc521, 
        A_DOUT(10) => nc1120, A_DOUT(9) => nc1051, A_DOUT(8) => 
        nc781, A_DOUT(7) => nc244, A_DOUT(6) => nc1008, A_DOUT(5)
         => nc538, A_DOUT(4) => nc1133, A_DOUT(3) => 
        b7_vFW_PlM(11), A_DOUT(2) => b7_vFW_PlM(10), A_DOUT(1)
         => b7_vFW_PlM(9), A_DOUT(0) => b7_vFW_PlM(8), B_DOUT(17)
         => nc291, B_DOUT(16) => nc195, B_DOUT(15) => nc1169, 
        B_DOUT(14) => nc958, B_DOUT(13) => nc66, B_DOUT(12) => 
        nc140, B_DOUT(11) => nc687, B_DOUT(10) => nc202, 
        B_DOUT(9) => nc1332, B_DOUT(8) => nc661, B_DOUT(7) => 
        nc545, B_DOUT(6) => nc794, B_DOUT(5) => nc390, B_DOUT(4)
         => nc1289, B_DOUT(3) => nc1033, B_DOUT(2) => nc230, 
        B_DOUT(1) => nc124, B_DOUT(0) => nc1027, BUSY => OPEN, 
        A_CLK => IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(11), B_DIN(2) => 
        b11_OFWNT9L_8tZ(10), B_DIN(1) => b11_OFWNT9L_8tZ(9), 
        B_DIN(0) => b11_OFWNT9L_8tZ(8), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_12 : RAM1K18
      port map(A_DOUT(17) => nc348, A_DOUT(16) => nc162, 
        A_DOUT(15) => nc423, A_DOUT(14) => nc751, A_DOUT(13) => 
        nc1230, A_DOUT(12) => nc628, A_DOUT(11) => nc1046, 
        A_DOUT(10) => nc212, A_DOUT(9) => nc283, A_DOUT(8) => 
        nc941, A_DOUT(7) => nc384, A_DOUT(6) => nc902, A_DOUT(5)
         => nc536, A_DOUT(4) => nc524, A_DOUT(3) => 
        b7_vFW_PlM(51), A_DOUT(2) => b7_vFW_PlM(50), A_DOUT(1)
         => b7_vFW_PlM(49), A_DOUT(0) => b7_vFW_PlM(48), 
        B_DOUT(17) => nc1223, B_DOUT(16) => nc226, B_DOUT(15) => 
        nc44, B_DOUT(14) => nc657, B_DOUT(13) => nc1231, 
        B_DOUT(12) => nc940, B_DOUT(11) => nc333, B_DOUT(10) => 
        nc435, B_DOUT(9) => nc1002, B_DOUT(8) => nc227, B_DOUT(7)
         => nc1262, B_DOUT(6) => nc912, B_DOUT(5) => nc802, 
        B_DOUT(4) => nc1004, B_DOUT(3) => nc974, B_DOUT(2) => 
        nc16, B_DOUT(1) => nc633, B_DOUT(0) => nc1108, BUSY => 
        OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(51), B_DIN(2) => 
        b11_OFWNT9L_8tZ(50), B_DIN(1) => b11_OFWNT9L_8tZ(49), 
        B_DIN(0) => b11_OFWNT9L_8tZ(48), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_SoW_b3_SoW_0_34 : RAM1K18
      port map(A_DOUT(17) => nc662, A_DOUT(16) => nc1227, 
        A_DOUT(15) => nc626, A_DOUT(14) => nc253, A_DOUT(13) => 
        nc354, A_DOUT(12) => nc1235, A_DOUT(11) => nc812, 
        A_DOUT(10) => nc447, A_DOUT(9) => nc1224, A_DOUT(8) => 
        nc1186, A_DOUT(7) => nc1137, A_DOUT(6) => nc834, 
        A_DOUT(5) => nc620, A_DOUT(4) => nc429, A_DOUT(3) => 
        b7_vFW_PlM(139), A_DOUT(2) => b7_vFW_PlM(138), A_DOUT(1)
         => b7_vFW_PlM(137), A_DOUT(0) => b7_vFW_PlM(136), 
        B_DOUT(17) => nc1340, B_DOUT(16) => nc1130, B_DOUT(15)
         => nc777, B_DOUT(14) => nc589, B_DOUT(13) => nc39, 
        B_DOUT(12) => nc738, B_DOUT(11) => nc395, B_DOUT(10) => 
        nc298, B_DOUT(9) => nc1218, B_DOUT(8) => nc1278, 
        B_DOUT(7) => nc342, B_DOUT(6) => nc446, B_DOUT(5) => 
        nc397, B_DOUT(4) => nc533, B_DOUT(3) => nc905, B_DOUT(2)
         => nc9, B_DOUT(1) => nc664, B_DOUT(0) => nc1189, BUSY
         => OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => 
        VCC_net_1, A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, 
        A_BLK(2) => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0)
         => VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N
         => VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        GND_net_1, A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, 
        A_DIN(13) => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11)
         => GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => 
        GND_net_1, A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, 
        A_DIN(6) => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4)
         => GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => 
        GND_net_1, A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, 
        A_ADDR(13) => b9_v_mzCDYXs(11), A_ADDR(12) => 
        b9_v_mzCDYXs(10), A_ADDR(11) => b9_v_mzCDYXs(9), 
        A_ADDR(10) => b9_v_mzCDYXs(8), A_ADDR(9) => 
        b9_v_mzCDYXs(7), A_ADDR(8) => b9_v_mzCDYXs(6), A_ADDR(7)
         => b9_v_mzCDYXs(5), A_ADDR(6) => b9_v_mzCDYXs(4), 
        A_ADDR(5) => b9_v_mzCDYXs(3), A_ADDR(4) => 
        b9_v_mzCDYXs(2), A_ADDR(3) => b9_v_mzCDYXs(1), A_ADDR(2)
         => b9_v_mzCDYXs(0), A_ADDR(1) => GND_net_1, A_ADDR(0)
         => GND_net_1, A_WEN(1) => GND_net_1, A_WEN(0) => 
        GND_net_1, B_CLK => CommsFPGA_CCC_0_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => VCC_net_1, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        GND_net_1, B_DIN(15) => GND_net_1, B_DIN(14) => GND_net_1, 
        B_DIN(13) => GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11)
         => GND_net_1, B_DIN(10) => GND_net_1, B_DIN(9) => 
        GND_net_1, B_DIN(8) => GND_net_1, B_DIN(7) => GND_net_1, 
        B_DIN(6) => GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4)
         => GND_net_1, B_DIN(3) => b11_OFWNT9L_8tZ(139), B_DIN(2)
         => b11_OFWNT9L_8tZ(138), B_DIN(1) => 
        b11_OFWNT9L_8tZ(137), B_DIN(0) => b11_OFWNT9L_8tZ(136), 
        B_ADDR(13) => b12_2_St6KCa_jHv(11), B_ADDR(12) => 
        b12_2_St6KCa_jHv(10), B_ADDR(11) => b12_2_St6KCa_jHv(9), 
        B_ADDR(10) => b12_2_St6KCa_jHv(8), B_ADDR(9) => 
        b12_2_St6KCa_jHv(7), B_ADDR(8) => b12_2_St6KCa_jHv(6), 
        B_ADDR(7) => b12_2_St6KCa_jHv(5), B_ADDR(6) => 
        b12_2_St6KCa_jHv(4), B_ADDR(5) => b12_2_St6KCa_jHv(3), 
        B_ADDR(4) => b12_2_St6KCa_jHv(2), B_ADDR(3) => 
        b12_2_St6KCa_jHv(1), B_ADDR(2) => b12_2_St6KCa_jHv(0), 
        B_ADDR(1) => GND_net_1, B_ADDR(0) => GND_net_1, B_WEN(1)
         => GND_net_1, B_WEN(0) => b4_2o_z, A_EN => VCC_net_1, 
        A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => GND_net_1, 
        A_WIDTH(1) => VCC_net_1, A_WIDTH(0) => GND_net_1, A_WMODE
         => VCC_net_1, B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, 
        B_WIDTH(2) => GND_net_1, B_WIDTH(1) => VCC_net_1, 
        B_WIDTH(0) => GND_net_1, B_WMODE => VCC_net_1, SII_LOCK
         => GND_net_1);
    
    b3_SoW_b3_SoW_0_21 : RAM1K18
      port map(A_DOUT(17) => nc1059, A_DOUT(16) => nc909, 
        A_DOUT(15) => nc1037, A_DOUT(14) => nc1001, A_DOUT(13)
         => nc349, A_DOUT(12) => nc294, A_DOUT(11) => nc915, 
        A_DOUT(10) => nc559, A_DOUT(9) => nc163, A_DOUT(8) => 
        nc101, A_DOUT(7) => nc107, A_DOUT(6) => nc821, A_DOUT(5)
         => nc919, A_DOUT(4) => nc186, A_DOUT(3) => 
        b7_vFW_PlM(87), A_DOUT(2) => b7_vFW_PlM(86), A_DOUT(1)
         => b7_vFW_PlM(85), A_DOUT(0) => b7_vFW_PlM(84), 
        B_DOUT(17) => nc190, B_DOUT(16) => nc28, B_DOUT(15) => 
        nc888, B_DOUT(14) => nc271, B_DOUT(13) => nc442, 
        B_DOUT(12) => nc1233, B_DOUT(11) => nc983, B_DOUT(10) => 
        nc175, B_DOUT(9) => nc209, B_DOUT(8) => nc947, B_DOUT(7)
         => nc635, B_DOUT(6) => nc595, B_DOUT(5) => nc225, 
        B_DOUT(4) => nc111, B_DOUT(3) => nc117, B_DOUT(2) => 
        nc398, B_DOUT(1) => nc774, B_DOUT(0) => nc370, BUSY => 
        OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(87), B_DIN(2) => 
        b11_OFWNT9L_8tZ(86), B_DIN(1) => b11_OFWNT9L_8tZ(85), 
        B_DIN(0) => b11_OFWNT9L_8tZ(84), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_3 : RAM1K18
      port map(A_DOUT(17) => nc1216, A_DOUT(16) => nc531, 
        A_DOUT(15) => nc1276, A_DOUT(14) => nc1282, A_DOUT(13)
         => nc991, A_DOUT(12) => nc219, A_DOUT(11) => nc1237, 
        A_DOUT(10) => nc763, A_DOUT(9) => nc468, A_DOUT(8) => 
        nc49, A_DOUT(7) => nc64, A_DOUT(6) => nc782, A_DOUT(5)
         => nc156, A_DOUT(4) => nc1192, A_DOUT(3) => 
        b7_vFW_PlM(15), A_DOUT(2) => b7_vFW_PlM(14), A_DOUT(1)
         => b7_vFW_PlM(13), A_DOUT(0) => b7_vFW_PlM(12), 
        B_DOUT(17) => nc641, B_DOUT(16) => nc25, B_DOUT(15) => 
        nc990, B_DOUT(14) => nc858, B_DOUT(13) => nc1234, 
        B_DOUT(12) => nc1028, B_DOUT(11) => nc953, B_DOUT(10) => 
        nc142, B_DOUT(9) => nc78, B_DOUT(8) => nc58, B_DOUT(7)
         => nc222, B_DOUT(6) => nc134, B_DOUT(5) => nc1095, 
        B_DOUT(4) => nc433, B_DOUT(3) => nc908, B_DOUT(2) => 
        nc638, B_DOUT(1) => nc497, B_DOUT(0) => nc752, BUSY => 
        OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(15), B_DIN(2) => 
        b11_OFWNT9L_8tZ(14), B_DIN(1) => b11_OFWNT9L_8tZ(13), 
        B_DIN(0) => b11_OFWNT9L_8tZ(12), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_13 : RAM1K18
      port map(A_DOUT(17) => nc534, A_DOUT(16) => nc236, 
        A_DOUT(15) => nc922, A_DOUT(14) => nc1304, A_DOUT(13) => 
        nc918, A_DOUT(12) => nc14, A_DOUT(11) => nc701, 
        A_DOUT(10) => nc37, A_DOUT(9) => nc237, A_DOUT(8) => 
        nc642, A_DOUT(7) => nc1114, A_DOUT(6) => nc885, A_DOUT(5)
         => nc375, A_DOUT(4) => nc75, A_DOUT(3) => b7_vFW_PlM(55), 
        A_DOUT(2) => b7_vFW_PlM(54), A_DOUT(1) => b7_vFW_PlM(53), 
        A_DOUT(0) => b7_vFW_PlM(52), B_DOUT(17) => nc278, 
        B_DOUT(16) => nc392, B_DOUT(15) => nc496, B_DOUT(14) => 
        nc1090, B_DOUT(13) => nc55, B_DOUT(12) => nc1174, 
        B_DOUT(11) => nc96, B_DOUT(10) => nc785, B_DOUT(9) => 
        nc1022, B_DOUT(8) => nc822, B_DOUT(7) => nc1024, 
        B_DOUT(6) => nc636, B_DOUT(5) => nc711, B_DOUT(4) => 
        nc377, B_DOUT(3) => nc1128, B_DOUT(2) => nc188, B_DOUT(1)
         => nc607, B_DOUT(0) => nc1009, BUSY => OPEN, A_CLK => 
        IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, A_ARST_N => 
        VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2) => VCC_net_1, 
        A_BLK(1) => VCC_net_1, A_BLK(0) => VCC_net_1, 
        A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => VCC_net_1, 
        A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, A_DIN(15)
         => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13) => 
        GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => GND_net_1, 
        A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, A_DIN(8)
         => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6) => 
        GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => GND_net_1, 
        A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, A_DIN(1)
         => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13) => 
        b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(55), B_DIN(2) => 
        b11_OFWNT9L_8tZ(54), B_DIN(1) => b11_OFWNT9L_8tZ(53), 
        B_DIN(0) => b11_OFWNT9L_8tZ(52), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_31 : RAM1K18
      port map(A_DOUT(17) => nc386, A_DOUT(16) => nc1317, 
        A_DOUT(15) => nc399, A_DOUT(14) => nc630, A_DOUT(13) => 
        nc439, A_DOUT(12) => nc274, A_DOUT(11) => nc617, 
        A_DOUT(10) => nc203, A_DOUT(9) => nc1111, A_DOUT(8) => 
        nc304, A_DOUT(7) => nc855, A_DOUT(6) => nc1171, A_DOUT(5)
         => nc689, A_DOUT(4) => nc492, A_DOUT(3) => 
        b7_vFW_PlM(127), A_DOUT(2) => b7_vFW_PlM(126), A_DOUT(1)
         => b7_vFW_PlM(125), A_DOUT(0) => b7_vFW_PlM(124), 
        B_DOUT(17) => nc755, B_DOUT(16) => nc997, B_DOUT(15) => 
        nc644, B_DOUT(14) => nc1145, B_DOUT(13) => nc170, 
        B_DOUT(12) => nc560, B_DOUT(11) => nc1038, B_DOUT(10) => 
        nc158, B_DOUT(9) => nc213, B_DOUT(8) => nc575, B_DOUT(7)
         => nc314, B_DOUT(6) => nc925, B_DOUT(5) => nc356, 
        B_DOUT(4) => nc378, B_DOUT(3) => nc143, B_DOUT(2) => 
        nc971, B_DOUT(1) => nc986, B_DOUT(0) => nc929, BUSY => 
        OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(127), B_DIN(2) => 
        b11_OFWNT9L_8tZ(126), B_DIN(1) => b11_OFWNT9L_8tZ(125), 
        B_DIN(0) => b11_OFWNT9L_8tZ(124), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_8 : RAM1K18
      port map(A_DOUT(17) => nc69, A_DOUT(16) => nc1021, 
        A_DOUT(15) => nc691, A_DOUT(14) => nc659, A_DOUT(13) => 
        nc831, A_DOUT(12) => nc121, A_DOUT(11) => nc47, 
        A_DOUT(10) => nc127, A_DOUT(9) => nc970, A_DOUT(8) => 
        nc381, A_DOUT(7) => nc235, A_DOUT(6) => nc1016, A_DOUT(5)
         => nc192, A_DOUT(4) => nc509, A_DOUT(3) => 
        b7_vFW_PlM(35), A_DOUT(2) => b7_vFW_PlM(34), A_DOUT(1)
         => b7_vFW_PlM(33), A_DOUT(0) => b7_vFW_PlM(32), 
        B_DOUT(17) => nc1076, B_DOUT(16) => nc229, B_DOUT(15) => 
        nc743, B_DOUT(14) => nc448, B_DOUT(13) => nc484, 
        B_DOUT(12) => nc1306, B_DOUT(11) => nc1032, B_DOUT(10)
         => nc1034, B_DOUT(9) => nc956, B_DOUT(8) => nc1268, 
        B_DOUT(7) => nc519, B_DOUT(6) => nc568, B_DOUT(5) => 
        nc477, B_DOUT(4) => nc1138, B_DOUT(3) => nc1152, 
        B_DOUT(2) => nc19, B_DOUT(1) => nc351, B_DOUT(0) => nc260, 
        BUSY => OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => 
        VCC_net_1, A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, 
        A_BLK(2) => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0)
         => VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N
         => VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        GND_net_1, A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, 
        A_DIN(13) => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11)
         => GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => 
        GND_net_1, A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, 
        A_DIN(6) => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4)
         => GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => 
        GND_net_1, A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, 
        A_ADDR(13) => b9_v_mzCDYXs(11), A_ADDR(12) => 
        b9_v_mzCDYXs(10), A_ADDR(11) => b9_v_mzCDYXs(9), 
        A_ADDR(10) => b9_v_mzCDYXs(8), A_ADDR(9) => 
        b9_v_mzCDYXs(7), A_ADDR(8) => b9_v_mzCDYXs(6), A_ADDR(7)
         => b9_v_mzCDYXs(5), A_ADDR(6) => b9_v_mzCDYXs(4), 
        A_ADDR(5) => b9_v_mzCDYXs(3), A_ADDR(4) => 
        b9_v_mzCDYXs(2), A_ADDR(3) => b9_v_mzCDYXs(1), A_ADDR(2)
         => b9_v_mzCDYXs(0), A_ADDR(1) => GND_net_1, A_ADDR(0)
         => GND_net_1, A_WEN(1) => GND_net_1, A_WEN(0) => 
        GND_net_1, B_CLK => CommsFPGA_CCC_0_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => VCC_net_1, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        GND_net_1, B_DIN(15) => GND_net_1, B_DIN(14) => GND_net_1, 
        B_DIN(13) => GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11)
         => GND_net_1, B_DIN(10) => GND_net_1, B_DIN(9) => 
        GND_net_1, B_DIN(8) => GND_net_1, B_DIN(7) => GND_net_1, 
        B_DIN(6) => GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4)
         => GND_net_1, B_DIN(3) => b11_OFWNT9L_8tZ(35), B_DIN(2)
         => b11_OFWNT9L_8tZ(34), B_DIN(1) => b11_OFWNT9L_8tZ(33), 
        B_DIN(0) => b11_OFWNT9L_8tZ(32), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_0 : RAM1K18
      port map(A_DOUT(17) => nc692, A_DOUT(16) => nc232, 
        A_DOUT(15) => nc372, A_DOUT(14) => nc476, A_DOUT(13) => 
        nc1055, A_DOUT(12) => nc106, A_DOUT(11) => nc454, 
        A_DOUT(10) => nc20, A_DOUT(9) => nc808, A_DOUT(8) => 
        nc566, A_DOUT(7) => nc1310, A_DOUT(6) => nc903, A_DOUT(5)
         => nc481, A_DOUT(4) => nc880, A_DOUT(3) => b7_vFW_PlM(3), 
        A_DOUT(2) => b7_vFW_PlM(2), A_DOUT(1) => b7_vFW_PlM(1), 
        A_DOUT(0) => b7_vFW_PlM(0), B_DOUT(17) => nc928, 
        B_DOUT(16) => nc883, B_DOUT(15) => nc116, B_DOUT(14) => 
        nc363, B_DOUT(13) => nc465, B_DOUT(12) => nc932, 
        B_DOUT(11) => nc379, B_DOUT(10) => nc21, B_DOUT(9) => 
        nc818, B_DOUT(8) => nc913, B_DOUT(7) => nc94, B_DOUT(6)
         => nc663, B_DOUT(5) => nc1266, B_DOUT(4) => nc1324, 
        B_DOUT(3) => nc1050, B_DOUT(2) => nc694, B_DOUT(1) => 
        nc1031, B_DOUT(0) => nc721, BUSY => OPEN, A_CLK => 
        IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, A_ARST_N => 
        VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2) => VCC_net_1, 
        A_BLK(1) => VCC_net_1, A_BLK(0) => VCC_net_1, 
        A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => VCC_net_1, 
        A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, A_DIN(15)
         => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13) => 
        GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => GND_net_1, 
        A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, A_DIN(8)
         => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6) => 
        GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => GND_net_1, 
        A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, A_DIN(1)
         => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13) => 
        b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(3), B_DIN(2) => 
        b11_OFWNT9L_8tZ(2), B_DIN(1) => b11_OFWNT9L_8tZ(1), 
        B_DIN(0) => b11_OFWNT9L_8tZ(0), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_7 : RAM1K18
      port map(A_DOUT(17) => nc1143, A_DOUT(16) => nc702, 
        A_DOUT(15) => nc472, A_DOUT(14) => nc832, A_DOUT(13) => 
        nc977, A_DOUT(12) => nc451, A_DOUT(11) => nc850, 
        A_DOUT(10) => nc1342, A_DOUT(9) => nc193, A_DOUT(8) => 
        nc1043, A_DOUT(7) => nc864, A_DOUT(6) => nc853, A_DOUT(5)
         => nc887, A_DOUT(4) => nc627, A_DOUT(3) => 
        b7_vFW_PlM(31), A_DOUT(2) => b7_vFW_PlM(30), A_DOUT(1)
         => b7_vFW_PlM(29), A_DOUT(0) => b7_vFW_PlM(28), 
        B_DOUT(17) => nc70, B_DOUT(16) => nc712, B_DOUT(15) => 
        nc50, B_DOUT(14) => nc1299, B_DOUT(13) => nc1029, 
        B_DOUT(12) => nc768, B_DOUT(11) => nc1240, B_DOUT(10) => 
        nc1301, B_DOUT(9) => nc67, B_DOUT(8) => nc540, B_DOUT(7)
         => nc789, B_DOUT(6) => nc563, B_DOUT(5) => nc71, 
        B_DOUT(4) => nc1288, B_DOUT(3) => nc671, B_DOUT(2) => 
        nc223, B_DOUT(1) => nc51, B_DOUT(0) => nc324, BUSY => 
        OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(31), B_DIN(2) => 
        b11_OFWNT9L_8tZ(30), B_DIN(1) => b11_OFWNT9L_8tZ(29), 
        B_DIN(0) => b11_OFWNT9L_8tZ(28), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_17 : RAM1K18
      port map(A_DOUT(17) => nc1241, A_DOUT(16) => nc172, 
        A_DOUT(15) => nc935, A_DOUT(14) => nc793, A_DOUT(13) => 
        nc498, A_DOUT(12) => nc857, A_DOUT(11) => nc805, 
        A_DOUT(10) => nc705, A_DOUT(9) => nc886, A_DOUT(8) => 
        nc1164, A_DOUT(7) => nc939, A_DOUT(6) => nc1245, 
        A_DOUT(5) => nc108, A_DOUT(4) => nc1102, A_DOUT(3) => 
        b7_vFW_PlM(71), A_DOUT(2) => b7_vFW_PlM(70), A_DOUT(1)
         => b7_vFW_PlM(69), A_DOUT(0) => b7_vFW_PlM(68), 
        B_DOUT(17) => nc815, B_DOUT(16) => nc759, B_DOUT(15) => 
        nc665, B_DOUT(14) => nc131, B_DOUT(13) => nc1147, 
        B_DOUT(12) => nc306, B_DOUT(11) => nc137, B_DOUT(10) => 
        nc715, B_DOUT(9) => nc889, B_DOUT(8) => nc17, B_DOUT(7)
         => nc1196, B_DOUT(6) => nc1140, B_DOUT(5) => nc672, 
        B_DOUT(4) => nc118, B_DOUT(3) => nc561, B_DOUT(2) => 
        nc239, B_DOUT(1) => nc1334, B_DOUT(0) => nc1005, BUSY => 
        OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(71), B_DIN(2) => 
        b11_OFWNT9L_8tZ(70), B_DIN(1) => b11_OFWNT9L_8tZ(69), 
        B_DIN(0) => b11_OFWNT9L_8tZ(68), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_28 : RAM1K18
      port map(A_DOUT(17) => nc529, A_DOUT(16) => nc609, 
        A_DOUT(15) => nc582, A_DOUT(14) => nc548, A_DOUT(13) => 
        nc316, A_DOUT(12) => nc1286, A_DOUT(11) => nc856, 
        A_DOUT(10) => nc1161, A_DOUT(9) => nc1326, A_DOUT(8) => 
        nc240, A_DOUT(7) => nc1315, A_DOUT(6) => nc1199, 
        A_DOUT(5) => nc619, A_DOUT(4) => nc859, A_DOUT(3) => 
        b7_vFW_PlM(115), A_DOUT(2) => b7_vFW_PlM(114), A_DOUT(1)
         => b7_vFW_PlM(113), A_DOUT(0) => b7_vFW_PlM(112), 
        B_DOUT(17) => nc99, B_DOUT(16) => nc1047, B_DOUT(15) => 
        nc88, B_DOUT(14) => nc480, B_DOUT(13) => nc1039, 
        B_DOUT(12) => nc164, B_DOUT(11) => nc906, B_DOUT(10) => 
        nc1000, B_DOUT(9) => nc463, B_DOUT(8) => nc546, B_DOUT(7)
         => nc674, B_DOUT(6) => nc668, B_DOUT(5) => nc552, 
        B_DOUT(4) => nc1243, B_DOUT(3) => nc301, B_DOUT(2) => 
        nc916, B_DOUT(1) => nc564, B_DOUT(0) => nc126, BUSY => 
        OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(115), B_DIN(2) => 
        b11_OFWNT9L_8tZ(114), B_DIN(1) => b11_OFWNT9L_8tZ(113), 
        B_DIN(0) => b11_OFWNT9L_8tZ(112), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_40 : RAM1K18
      port map(A_DOUT(17) => nc266, A_DOUT(16) => nc343, 
        A_DOUT(15) => nc445, A_DOUT(14) => nc22, A_DOUT(13) => 
        nc938, A_DOUT(12) => nc828, A_DOUT(11) => nc923, 
        A_DOUT(10) => nc173, A_DOUT(9) => nc643, A_DOUT(8) => 
        nc1066, A_DOUT(7) => nc1115, A_DOUT(6) => nc267, 
        A_DOUT(5) => nc85, A_DOUT(4) => nc1175, A_DOUT(3) => 
        b7_vFW_PlM(163), A_DOUT(2) => b7_vFW_PlM(162), A_DOUT(1)
         => b7_vFW_PlM(161), A_DOUT(0) => b7_vFW_PlM(160), 
        B_DOUT(17) => nc404, B_DOUT(16) => nc450, B_DOUT(15) => 
        nc311, B_DOUT(14) => nc1292, B_DOUT(13) => nc1247, 
        B_DOUT(12) => nc590, B_DOUT(11) => nc731, B_DOUT(10) => 
        nc666, B_DOUT(9) => nc1184, B_DOUT(8) => nc1244, 
        B_DOUT(7) => nc844, B_DOUT(6) => nc414, B_DOUT(5) => 
        nc722, B_DOUT(4) => nc587, B_DOUT(3) => nc748, B_DOUT(2)
         => nc660, B_DOUT(1) => nc469, B_DOUT(0) => nc773, BUSY
         => OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => 
        VCC_net_1, A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, 
        A_BLK(2) => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0)
         => VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N
         => VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        GND_net_1, A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, 
        A_DIN(13) => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11)
         => GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => 
        GND_net_1, A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, 
        A_DIN(6) => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4)
         => GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => 
        GND_net_1, A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, 
        A_ADDR(13) => b9_v_mzCDYXs(11), A_ADDR(12) => 
        b9_v_mzCDYXs(10), A_ADDR(11) => b9_v_mzCDYXs(9), 
        A_ADDR(10) => b9_v_mzCDYXs(8), A_ADDR(9) => 
        b9_v_mzCDYXs(7), A_ADDR(8) => b9_v_mzCDYXs(6), A_ADDR(7)
         => b9_v_mzCDYXs(5), A_ADDR(6) => b9_v_mzCDYXs(4), 
        A_ADDR(5) => b9_v_mzCDYXs(3), A_ADDR(4) => 
        b9_v_mzCDYXs(2), A_ADDR(3) => b9_v_mzCDYXs(1), A_ADDR(2)
         => b9_v_mzCDYXs(0), A_ADDR(1) => GND_net_1, A_ADDR(0)
         => GND_net_1, A_WEN(1) => GND_net_1, A_WEN(0) => 
        GND_net_1, B_CLK => CommsFPGA_CCC_0_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => VCC_net_1, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        GND_net_1, B_DIN(15) => GND_net_1, B_DIN(14) => GND_net_1, 
        B_DIN(13) => GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11)
         => GND_net_1, B_DIN(10) => GND_net_1, B_DIN(9) => 
        GND_net_1, B_DIN(8) => GND_net_1, B_DIN(7) => GND_net_1, 
        B_DIN(6) => GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4)
         => GND_net_1, B_DIN(3) => b11_OFWNT9L_8tZ(163), B_DIN(2)
         => b11_OFWNT9L_8tZ(162), B_DIN(1) => 
        b11_OFWNT9L_8tZ(161), B_DIN(0) => b11_OFWNT9L_8tZ(160), 
        B_ADDR(13) => b12_2_St6KCa_jHv(11), B_ADDR(12) => 
        b12_2_St6KCa_jHv(10), B_ADDR(11) => b12_2_St6KCa_jHv(9), 
        B_ADDR(10) => b12_2_St6KCa_jHv(8), B_ADDR(9) => 
        b12_2_St6KCa_jHv(7), B_ADDR(8) => b12_2_St6KCa_jHv(6), 
        B_ADDR(7) => b12_2_St6KCa_jHv(5), B_ADDR(6) => 
        b12_2_St6KCa_jHv(4), B_ADDR(5) => b12_2_St6KCa_jHv(3), 
        B_ADDR(4) => b12_2_St6KCa_jHv(2), B_ADDR(3) => 
        b12_2_St6KCa_jHv(1), B_ADDR(2) => b12_2_St6KCa_jHv(0), 
        B_ADDR(1) => GND_net_1, B_ADDR(0) => GND_net_1, B_WEN(1)
         => GND_net_1, B_WEN(0) => b4_2o_z, A_EN => VCC_net_1, 
        A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => GND_net_1, 
        A_WIDTH(1) => VCC_net_1, A_WIDTH(0) => GND_net_1, A_WMODE
         => VCC_net_1, B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, 
        B_WIDTH(2) => GND_net_1, B_WIDTH(1) => VCC_net_1, 
        B_WIDTH(0) => GND_net_1, B_WMODE => VCC_net_1, SII_LOCK
         => GND_net_1);
    
    b3_SoW_b3_SoW_0_38 : RAM1K18
      port map(A_DOUT(17) => nc637, A_DOUT(16) => nc478, 
        A_DOUT(15) => nc1259, A_DOUT(14) => nc72, A_DOUT(13) => 
        nc52, A_DOUT(12) => nc543, A_DOUT(11) => nc401, 
        A_DOUT(10) => nc800, A_DOUT(9) => nc1181, A_DOUT(8) => 
        nc1336, A_DOUT(7) => nc233, A_DOUT(6) => nc803, A_DOUT(5)
         => nc1321, A_DOUT(4) => nc334, A_DOUT(3) => 
        b7_vFW_PlM(155), A_DOUT(2) => b7_vFW_PlM(154), A_DOUT(1)
         => b7_vFW_PlM(153), A_DOUT(0) => b7_vFW_PlM(152), 
        B_DOUT(17) => nc780, B_DOUT(16) => nc557, B_DOUT(15) => 
        nc411, B_DOUT(14) => nc810, B_DOUT(13) => nc598, 
        B_DOUT(12) => nc1318, B_DOUT(11) => nc813, B_DOUT(10) => 
        nc825, B_DOUT(9) => nc645, B_DOUT(8) => nc861, B_DOUT(7)
         => nc725, B_DOUT(6) => nc290, B_DOUT(5) => nc189, 
        B_DOUT(4) => nc265, B_DOUT(3) => nc128, B_DOUT(2) => 
        nc807, B_DOUT(1) => nc541, B_DOUT(0) => nc1156, BUSY => 
        OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(155), B_DIN(2) => 
        b11_OFWNT9L_8tZ(154), B_DIN(1) => b11_OFWNT9L_8tZ(153), 
        B_DIN(0) => b11_OFWNT9L_8tZ(152), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_15 : RAM1K18
      port map(A_DOUT(17) => nc1122, A_DOUT(16) => nc786, 
        A_DOUT(15) => nc97, A_DOUT(14) => nc750, A_DOUT(13) => 
        nc326, A_DOUT(12) => nc1086, A_DOUT(11) => nc596, 
        A_DOUT(10) => nc539, A_DOUT(9) => nc817, A_DOUT(8) => 
        nc709, A_DOUT(7) => nc1025, A_DOUT(6) => nc393, A_DOUT(5)
         => nc495, A_DOUT(4) => nc629, A_DOUT(3) => 
        b7_vFW_PlM(63), A_DOUT(2) => b7_vFW_PlM(62), A_DOUT(1)
         => b7_vFW_PlM(61), A_DOUT(0) => b7_vFW_PlM(60), 
        B_DOUT(17) => nc1048, B_DOUT(16) => nc693, B_DOUT(15) => 
        nc159, B_DOUT(14) => nc1159, B_DOUT(13) => nc144, 
        B_DOUT(12) => nc719, B_DOUT(11) => nc1113, B_DOUT(10) => 
        nc1173, B_DOUT(9) => nc756, B_DOUT(8) => nc443, B_DOUT(7)
         => nc806, B_DOUT(6) => nc648, B_DOUT(5) => nc262, 
        B_DOUT(4) => nc1312, B_DOUT(3) => nc570, B_DOUT(2) => 
        nc1013, B_DOUT(1) => nc1073, B_DOUT(0) => nc926, BUSY => 
        OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(63), B_DIN(2) => 
        b11_OFWNT9L_8tZ(62), B_DIN(1) => b11_OFWNT9L_8tZ(61), 
        B_DIN(0) => b11_OFWNT9L_8tZ(60), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_10 : RAM1K18
      port map(A_DOUT(17) => nc894, A_DOUT(16) => nc544, 
        A_DOUT(15) => nc1020, A_DOUT(14) => nc246, A_DOUT(13) => 
        nc1331, A_DOUT(12) => nc816, A_DOUT(11) => nc809, 
        A_DOUT(10) => nc1210, A_DOUT(9) => nc798, A_DOUT(8) => 
        nc1270, A_DOUT(7) => nc136, A_DOUT(6) => nc23, A_DOUT(5)
         => nc962, A_DOUT(4) => nc838, A_DOUT(3) => 
        b7_vFW_PlM(43), A_DOUT(2) => b7_vFW_PlM(42), A_DOUT(1)
         => b7_vFW_PlM(41), A_DOUT(0) => b7_vFW_PlM(40), 
        B_DOUT(17) => nc247, B_DOUT(16) => nc933, B_DOUT(15) => 
        nc321, B_DOUT(14) => nc1209, B_DOUT(13) => nc593, 
        B_DOUT(12) => nc502, B_DOUT(11) => nc1042, B_DOUT(10) => 
        nc984, B_DOUT(9) => nc819, B_DOUT(8) => nc646, B_DOUT(7)
         => nc1252, B_DOUT(6) => nc1044, B_DOUT(5) => nc1211, 
        B_DOUT(4) => nc1271, B_DOUT(3) => nc1148, B_DOUT(2) => 
        nc862, B_DOUT(1) => nc424, B_DOUT(0) => nc512, BUSY => 
        OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(43), B_DIN(2) => 
        b11_OFWNT9L_8tZ(42), B_DIN(1) => b11_OFWNT9L_8tZ(41), 
        B_DIN(0) => b11_OFWNT9L_8tZ(40), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_6 : RAM1K18
      port map(A_DOUT(17) => nc640, A_DOUT(16) => nc449, 
        A_DOUT(15) => nc80, A_DOUT(14) => nc732, A_DOUT(13) => 
        nc1132, A_DOUT(12) => nc400, A_DOUT(11) => nc1215, 
        A_DOUT(10) => nc1275, A_DOUT(9) => nc787, A_DOUT(8) => 
        nc578, A_DOUT(7) => nc1117, A_DOUT(6) => nc695, A_DOUT(5)
         => nc1177, A_DOUT(4) => nc954, A_DOUT(3) => 
        b7_vFW_PlM(27), A_DOUT(2) => b7_vFW_PlM(26), A_DOUT(1)
         => b7_vFW_PlM(25), A_DOUT(0) => b7_vFW_PlM(24), 
        B_DOUT(17) => nc73, B_DOUT(16) => nc81, B_DOUT(15) => 
        nc1110, B_DOUT(14) => nc53, B_DOUT(13) => nc410, 
        B_DOUT(12) => nc1170, B_DOUT(11) => nc1035, B_DOUT(10)
         => nc270, B_DOUT(9) => nc591, B_DOUT(8) => nc421, 
        B_DOUT(7) => nc820, B_DOUT(6) => nc1106, B_DOUT(5) => 
        nc965, B_DOUT(4) => nc823, B_DOUT(3) => nc576, B_DOUT(2)
         => nc1165, B_DOUT(1) => nc757, B_DOUT(0) => nc1041, BUSY
         => OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => 
        VCC_net_1, A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, 
        A_BLK(2) => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0)
         => VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N
         => VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        GND_net_1, A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, 
        A_DIN(13) => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11)
         => GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => 
        GND_net_1, A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, 
        A_DIN(6) => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4)
         => GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => 
        GND_net_1, A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, 
        A_ADDR(13) => b9_v_mzCDYXs(11), A_ADDR(12) => 
        b9_v_mzCDYXs(10), A_ADDR(11) => b9_v_mzCDYXs(9), 
        A_ADDR(10) => b9_v_mzCDYXs(8), A_ADDR(9) => 
        b9_v_mzCDYXs(7), A_ADDR(8) => b9_v_mzCDYXs(6), A_ADDR(7)
         => b9_v_mzCDYXs(5), A_ADDR(6) => b9_v_mzCDYXs(4), 
        A_ADDR(5) => b9_v_mzCDYXs(3), A_ADDR(4) => 
        b9_v_mzCDYXs(2), A_ADDR(3) => b9_v_mzCDYXs(1), A_ADDR(2)
         => b9_v_mzCDYXs(0), A_ADDR(1) => GND_net_1, A_ADDR(0)
         => GND_net_1, A_WEN(1) => GND_net_1, A_WEN(0) => 
        GND_net_1, B_CLK => CommsFPGA_CCC_0_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => VCC_net_1, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        GND_net_1, B_DIN(15) => GND_net_1, B_DIN(14) => GND_net_1, 
        B_DIN(13) => GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11)
         => GND_net_1, B_DIN(10) => GND_net_1, B_DIN(9) => 
        GND_net_1, B_DIN(8) => GND_net_1, B_DIN(7) => GND_net_1, 
        B_DIN(6) => GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4)
         => GND_net_1, B_DIN(3) => b11_OFWNT9L_8tZ(27), B_DIN(2)
         => b11_OFWNT9L_8tZ(26), B_DIN(1) => b11_OFWNT9L_8tZ(25), 
        B_DIN(0) => b11_OFWNT9L_8tZ(24), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_22 : RAM1K18
      port map(A_DOUT(17) => nc969, A_DOUT(16) => nc841, 
        A_DOUT(15) => nc1017, A_DOUT(14) => nc1030, A_DOUT(13)
         => nc835, A_DOUT(12) => nc1077, A_DOUT(11) => nc245, 
        A_DOUT(10) => nc161, A_DOUT(9) => nc373, A_DOUT(8) => 
        nc475, A_DOUT(7) => nc735, A_DOUT(6) => nc167, A_DOUT(5)
         => nc281, A_DOUT(4) => nc194, A_DOUT(3) => 
        b7_vFW_PlM(91), A_DOUT(2) => b7_vFW_PlM(90), A_DOUT(1)
         => b7_vFW_PlM(89), A_DOUT(0) => b7_vFW_PlM(88), 
        B_DOUT(17) => nc507, B_DOUT(16) => nc185, B_DOUT(15) => 
        nc1109, B_DOUT(14) => nc673, B_DOUT(13) => nc493, 
        B_DOUT(12) => nc138, B_DOUT(11) => nc698, B_DOUT(10) => 
        nc269, B_DOUT(9) => nc1213, B_DOUT(8) => nc784, B_DOUT(7)
         => nc380, B_DOUT(6) => nc1273, B_DOUT(5) => nc336, 
        B_DOUT(4) => nc827, B_DOUT(3) => nc517, B_DOUT(2) => 
        nc594, B_DOUT(1) => nc296, B_DOUT(0) => nc874, BUSY => 
        OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(91), B_DIN(2) => 
        b11_OFWNT9L_8tZ(90), B_DIN(1) => b11_OFWNT9L_8tZ(89), 
        B_DIN(0) => b11_OFWNT9L_8tZ(88), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_19 : RAM1K18
      port map(A_DOUT(17) => nc1298, A_DOUT(16) => nc639, 
        A_DOUT(15) => nc729, A_DOUT(14) => nc297, A_DOUT(13) => 
        nc1217, A_DOUT(12) => nc778, A_DOUT(11) => nc700, 
        A_DOUT(10) => nc251, A_DOUT(9) => nc1277, A_DOUT(8) => 
        nc155, A_DOUT(7) => nc242, A_DOUT(6) => nc696, A_DOUT(5)
         => nc1214, A_DOUT(4) => nc754, A_DOUT(3) => 
        b7_vFW_PlM(79), A_DOUT(2) => b7_vFW_PlM(78), A_DOUT(1)
         => b7_vFW_PlM(77), A_DOUT(0) => b7_vFW_PlM(76), 
        B_DOUT(17) => nc573, B_DOUT(16) => nc350, B_DOUT(15) => 
        nc1202, B_DOUT(14) => nc1274, B_DOUT(13) => nc710, 
        B_DOUT(12) => nc826, B_DOUT(11) => nc109, B_DOUT(10) => 
        nc936, B_DOUT(9) => nc690, B_DOUT(8) => nc499, B_DOUT(7)
         => nc942, B_DOUT(6) => nc1303, B_DOUT(5) => nc968, 
        B_DOUT(4) => nc706, B_DOUT(3) => nc829, B_DOUT(2) => 
        nc119, B_DOUT(1) => nc331, B_DOUT(0) => nc1344, BUSY => 
        OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(79), B_DIN(2) => 
        b11_OFWNT9L_8tZ(78), B_DIN(1) => b11_OFWNT9L_8tZ(77), 
        B_DIN(0) => b11_OFWNT9L_8tZ(76), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_9 : RAM1K18
      port map(A_DOUT(17) => nc38, A_DOUT(16) => nc842, 
        A_DOUT(15) => nc385, A_DOUT(14) => nc288, A_DOUT(13) => 
        nc1185, A_DOUT(12) => nc675, A_DOUT(11) => nc1229, 
        A_DOUT(10) => nc1296, A_DOUT(9) => nc761, A_DOUT(8) => 
        nc716, A_DOUT(7) => nc522, A_DOUT(6) => nc434, A_DOUT(5)
         => nc387, A_DOUT(4) => nc571, A_DOUT(3) => 
        b7_vFW_PlM(39), A_DOUT(2) => b7_vFW_PlM(38), A_DOUT(1)
         => b7_vFW_PlM(37), A_DOUT(0) => b7_vFW_PlM(36), 
        B_DOUT(17) => nc1049, B_DOUT(16) => nc667, B_DOUT(15) => 
        nc1163, B_DOUT(14) => nc891, B_DOUT(13) => nc2, 
        B_DOUT(12) => nc82, B_DOUT(11) => nc284, B_DOUT(10) => 
        nc420, B_DOUT(9) => nc35, B_DOUT(8) => nc295, B_DOUT(7)
         => nc355, B_DOUT(6) => nc258, B_DOUT(5) => nc1063, 
        B_DOUT(4) => nc263, B_DOUT(3) => nc180, B_DOUT(2) => 
        nc364, B_DOUT(1) => nc357, B_DOUT(0) => nc174, BUSY => 
        OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(39), B_DIN(2) => 
        b11_OFWNT9L_8tZ(38), B_DIN(1) => b11_OFWNT9L_8tZ(37), 
        B_DIN(0) => b11_OFWNT9L_8tZ(36), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_23 : RAM1K18
      port map(A_DOUT(17) => nc945, A_DOUT(16) => nc585, 
        A_DOUT(15) => nc1260, A_DOUT(14) => nc431, A_DOUT(13) => 
        nc830, A_DOUT(12) => nc473, A_DOUT(11) => nc678, 
        A_DOUT(10) => nc388, A_DOUT(9) => nc904, A_DOUT(8) => 
        nc833, A_DOUT(7) => nc1018, A_DOUT(6) => nc949, A_DOUT(5)
         => nc1126, A_DOUT(4) => nc1078, A_DOUT(3) => 
        b7_vFW_PlM(95), A_DOUT(2) => b7_vFW_PlM(94), A_DOUT(1)
         => b7_vFW_PlM(93), A_DOUT(0) => b7_vFW_PlM(92), 
        B_DOUT(17) => nc981, B_DOUT(16) => nc254, B_DOUT(15) => 
        nc574, B_DOUT(14) => nc141, B_DOUT(13) => nc276, 
        B_DOUT(12) => nc1261, B_DOUT(11) => nc147, B_DOUT(10) => 
        nc1194, B_DOUT(9) => nc914, B_DOUT(8) => nc48, B_DOUT(7)
         => nc7, B_DOUT(6) => nc5, B_DOUT(5) => nc150, B_DOUT(4)
         => nc277, B_DOUT(3) => nc292, B_DOUT(2) => nc980, 
        B_DOUT(1) => nc249, B_DOUT(0) => nc707, BUSY => OPEN, 
        A_CLK => IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(95), B_DIN(2) => 
        b11_OFWNT9L_8tZ(94), B_DIN(1) => b11_OFWNT9L_8tZ(93), 
        B_DIN(0) => b11_OFWNT9L_8tZ(92), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_32 : RAM1K18
      port map(A_DOUT(17) => nc555, A_DOUT(16) => nc527, 
        A_DOUT(15) => nc1129, A_DOUT(14) => nc676, A_DOUT(13) => 
        nc1265, A_DOUT(12) => nc358, A_DOUT(11) => nc837, 
        A_DOUT(10) => nc569, A_DOUT(9) => nc1239, A_DOUT(8) => 
        nc1167, A_DOUT(7) => nc951, A_DOUT(6) => nc717, A_DOUT(5)
         => nc992, A_DOUT(4) => nc487, A_DOUT(3) => 
        b7_vFW_PlM(131), A_DOUT(2) => b7_vFW_PlM(130), A_DOUT(1)
         => b7_vFW_PlM(129), A_DOUT(0) => b7_vFW_PlM(128), 
        B_DOUT(17) => nc1160, B_DOUT(16) => nc1191, B_DOUT(15)
         => nc1258, B_DOUT(14) => nc670, B_DOUT(13) => nc479, 
        B_DOUT(12) => nc1012, B_DOUT(11) => nc45, B_DOUT(10) => 
        nc1072, B_DOUT(9) => nc1014, B_DOUT(8) => nc739, 
        B_DOUT(7) => nc1074, B_DOUT(6) => nc1118, B_DOUT(5) => 
        nc950, B_DOUT(4) => nc1309, B_DOUT(3) => nc1178, 
        B_DOUT(2) => nc892, B_DOUT(1) => nc720, B_DOUT(0) => 
        nc1183, BUSY => OPEN, A_CLK => IICE_comm2iice_0, 
        A_DOUT_CLK => VCC_net_1, A_ARST_N => VCC_net_1, A_DOUT_EN
         => VCC_net_1, A_BLK(2) => VCC_net_1, A_BLK(1) => 
        VCC_net_1, A_BLK(0) => VCC_net_1, A_DOUT_ARST_N => 
        VCC_net_1, A_DOUT_SRST_N => VCC_net_1, A_DIN(17) => 
        GND_net_1, A_DIN(16) => GND_net_1, A_DIN(15) => GND_net_1, 
        A_DIN(14) => GND_net_1, A_DIN(13) => GND_net_1, A_DIN(12)
         => GND_net_1, A_DIN(11) => GND_net_1, A_DIN(10) => 
        GND_net_1, A_DIN(9) => GND_net_1, A_DIN(8) => GND_net_1, 
        A_DIN(7) => GND_net_1, A_DIN(6) => GND_net_1, A_DIN(5)
         => GND_net_1, A_DIN(4) => GND_net_1, A_DIN(3) => 
        GND_net_1, A_DIN(2) => GND_net_1, A_DIN(1) => GND_net_1, 
        A_DIN(0) => GND_net_1, A_ADDR(13) => b9_v_mzCDYXs(11), 
        A_ADDR(12) => b9_v_mzCDYXs(10), A_ADDR(11) => 
        b9_v_mzCDYXs(9), A_ADDR(10) => b9_v_mzCDYXs(8), A_ADDR(9)
         => b9_v_mzCDYXs(7), A_ADDR(8) => b9_v_mzCDYXs(6), 
        A_ADDR(7) => b9_v_mzCDYXs(5), A_ADDR(6) => 
        b9_v_mzCDYXs(4), A_ADDR(5) => b9_v_mzCDYXs(3), A_ADDR(4)
         => b9_v_mzCDYXs(2), A_ADDR(3) => b9_v_mzCDYXs(1), 
        A_ADDR(2) => b9_v_mzCDYXs(0), A_ADDR(1) => GND_net_1, 
        A_ADDR(0) => GND_net_1, A_WEN(1) => GND_net_1, A_WEN(0)
         => GND_net_1, B_CLK => CommsFPGA_CCC_0_GL0, B_DOUT_CLK
         => VCC_net_1, B_ARST_N => VCC_net_1, B_DOUT_EN => 
        VCC_net_1, B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, 
        B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, 
        B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => GND_net_1, 
        B_DIN(16) => GND_net_1, B_DIN(15) => GND_net_1, B_DIN(14)
         => GND_net_1, B_DIN(13) => GND_net_1, B_DIN(12) => 
        GND_net_1, B_DIN(11) => GND_net_1, B_DIN(10) => GND_net_1, 
        B_DIN(9) => GND_net_1, B_DIN(8) => GND_net_1, B_DIN(7)
         => GND_net_1, B_DIN(6) => GND_net_1, B_DIN(5) => 
        GND_net_1, B_DIN(4) => GND_net_1, B_DIN(3) => 
        b11_OFWNT9L_8tZ(131), B_DIN(2) => b11_OFWNT9L_8tZ(130), 
        B_DIN(1) => b11_OFWNT9L_8tZ(129), B_DIN(0) => 
        b11_OFWNT9L_8tZ(128), B_ADDR(13) => b12_2_St6KCa_jHv(11), 
        B_ADDR(12) => b12_2_St6KCa_jHv(10), B_ADDR(11) => 
        b12_2_St6KCa_jHv(9), B_ADDR(10) => b12_2_St6KCa_jHv(8), 
        B_ADDR(9) => b12_2_St6KCa_jHv(7), B_ADDR(8) => 
        b12_2_St6KCa_jHv(6), B_ADDR(7) => b12_2_St6KCa_jHv(5), 
        B_ADDR(6) => b12_2_St6KCa_jHv(4), B_ADDR(5) => 
        b12_2_St6KCa_jHv(3), B_ADDR(4) => b12_2_St6KCa_jHv(2), 
        B_ADDR(3) => b12_2_St6KCa_jHv(1), B_ADDR(2) => 
        b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, B_ADDR(0)
         => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0) => b4_2o_z, 
        A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, A_WIDTH(2)
         => GND_net_1, A_WIDTH(1) => VCC_net_1, A_WIDTH(0) => 
        GND_net_1, A_WMODE => VCC_net_1, B_EN => VCC_net_1, 
        B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => GND_net_1, 
        B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => GND_net_1, B_WMODE
         => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_16 : RAM1K18
      port map(A_DOUT(17) => nc382, A_DOUT(16) => nc486, 
        A_DOUT(15) => nc1222, A_DOUT(14) => nc836, A_DOUT(13) => 
        nc201, A_DOUT(12) => nc948, A_DOUT(11) => nc105, 
        A_DOUT(10) => nc1067, A_DOUT(9) => nc1083, A_DOUT(8) => 
        nc457, A_DOUT(7) => nc166, A_DOUT(6) => nc26, A_DOUT(5)
         => nc868, A_DOUT(4) => nc129, A_DOUT(3) => 
        b7_vFW_PlM(67), A_DOUT(2) => b7_vFW_PlM(66), A_DOUT(1)
         => b7_vFW_PlM(65), A_DOUT(0) => b7_vFW_PlM(64), 
        B_DOUT(17) => nc963, B_DOUT(16) => nc704, B_DOUT(15) => 
        nc300, B_DOUT(14) => nc1280, B_DOUT(13) => nc389, 
        B_DOUT(12) => nc1323, B_DOUT(11) => nc839, B_DOUT(10) => 
        nc211, B_DOUT(9) => nc1136, B_DOUT(8) => nc115, B_DOUT(7)
         => nc1096, B_DOUT(6) => nc871, B_DOUT(5) => nc726, 
        B_DOUT(4) => nc1263, B_DOUT(3) => nc741, B_DOUT(2) => 
        nc1256, B_DOUT(1) => nc275, B_DOUT(0) => nc352, BUSY => 
        OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(67), B_DIN(2) => 
        b11_OFWNT9L_8tZ(66), B_DIN(1) => b11_OFWNT9L_8tZ(65), 
        B_DIN(0) => b11_OFWNT9L_8tZ(64), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_4 : RAM1K18
      port map(A_DOUT(17) => nc456, A_DOUT(16) => nc714, 
        A_DOUT(15) => nc310, A_DOUT(14) => nc482, A_DOUT(13) => 
        nc532, A_DOUT(12) => nc1281, A_DOUT(11) => nc995, 
        A_DOUT(10) => nc987, A_DOUT(9) => nc1011, A_DOUT(8) => 
        nc1071, A_DOUT(7) => nc762, A_DOUT(6) => nc647, A_DOUT(5)
         => nc1267, A_DOUT(4) => nc999, A_DOUT(3) => 
        b7_vFW_PlM(19), A_DOUT(2) => b7_vFW_PlM(18), A_DOUT(1)
         => b7_vFW_PlM(17), A_DOUT(0) => b7_vFW_PlM(16), 
        B_DOUT(17) => nc1139, B_DOUT(16) => nc359, B_DOUT(15) => 
        nc191, B_DOUT(14) => nc1285, B_DOUT(13) => nc83, 
        B_DOUT(12) => nc197, B_DOUT(11) => nc1264, B_DOUT(10) => 
        nc430, B_DOUT(9) => nc76, B_DOUT(8) => nc56, B_DOUT(7)
         => nc243, B_DOUT(6) => nc68, B_DOUT(5) => nc1187, 
        B_DOUT(4) => nc344, B_DOUT(3) => nc1341, B_DOUT(2) => 
        nc681, B_DOUT(1) => nc452, B_DOUT(0) => nc299, BUSY => 
        OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(19), B_DIN(2) => 
        b11_OFWNT9L_8tZ(18), B_DIN(1) => b11_OFWNT9L_8tZ(17), 
        B_DIN(0) => b11_OFWNT9L_8tZ(16), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_33 : RAM1K18
      port map(A_DOUT(17) => nc1180, A_DOUT(16) => nc957, 
        A_DOUT(15) => nc272, A_DOUT(14) => nc182, A_DOUT(13) => 
        nc30, A_DOUT(12) => nc305, A_DOUT(11) => nc208, 
        A_DOUT(10) => nc924, A_DOUT(9) => nc865, A_DOUT(8) => 
        nc1232, A_DOUT(7) => nc307, A_DOUT(6) => nc31, A_DOUT(5)
         => nc1208, A_DOUT(4) => nc1154, A_DOUT(3) => 
        b7_vFW_PlM(135), A_DOUT(2) => b7_vFW_PlM(134), A_DOUT(1)
         => b7_vFW_PlM(133), A_DOUT(0) => b7_vFW_PlM(132), 
        B_DOUT(17) => nc972, B_DOUT(16) => nc765, B_DOUT(15) => 
        nc65, B_DOUT(14) => nc315, B_DOUT(13) => nc218, 
        B_DOUT(12) => nc1087, B_DOUT(11) => nc651, B_DOUT(10) => 
        nc1142, B_DOUT(9) => nc168, B_DOUT(8) => nc18, B_DOUT(7)
         => nc1333, B_DOUT(6) => nc317, B_DOUT(5) => nc682, 
        B_DOUT(4) => nc549, B_DOUT(3) => nc366, B_DOUT(2) => 
        nc152, B_DOUT(1) => nc204, B_DOUT(0) => nc872, BUSY => 
        OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(135), B_DIN(2) => 
        b11_OFWNT9L_8tZ(134), B_DIN(1) => b11_OFWNT9L_8tZ(133), 
        B_DIN(0) => b11_OFWNT9L_8tZ(132), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    
    b3_SoW_b3_SoW_0_41 : RAM1K18
      port map(A_DOUT(17) => nc537, A_DOUT(16) => nc727, 
        A_DOUT(15) => nc1283, A_DOUT(14) => nc1045, A_DOUT(13)
         => nc998, A_DOUT(12) => nc100, A_DOUT(11) => nc1314, 
        A_DOUT(10) => nc669, A_DOUT(9) => nc214, A_DOUT(8) => 
        nc1151, A_DOUT(7) => nc505, A_DOUT(6) => nc308, A_DOUT(5)
         => nc1287, A_DOUT(4) => nc791, A_DOUT(3) => 
        b7_vFW_PlM(167), A_DOUT(2) => b7_vFW_PlM(166), A_DOUT(1)
         => b7_vFW_PlM(165), A_DOUT(0) => b7_vFW_PlM(164), 
        B_DOUT(17) => nc15, B_DOUT(16) => nc110, B_DOUT(15) => 
        nc901, B_DOUT(14) => nc730, B_DOUT(13) => nc652, 
        B_DOUT(12) => nc515, B_DOUT(11) => nc1068, B_DOUT(10) => 
        nc1329, B_DOUT(9) => nc1206, B_DOUT(8) => nc1040, 
        B_DOUT(7) => nc684, B_DOUT(6) => nc1284, B_DOUT(5) => 
        nc318, B_DOUT(4) => nc1019, B_DOUT(3) => nc966, B_DOUT(2)
         => nc40, B_DOUT(1) => nc1079, B_DOUT(0) => nc146, BUSY
         => OPEN, A_CLK => IICE_comm2iice_0, A_DOUT_CLK => 
        VCC_net_1, A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, 
        A_BLK(2) => VCC_net_1, A_BLK(1) => VCC_net_1, A_BLK(0)
         => VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N
         => VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => 
        GND_net_1, A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, 
        A_DIN(13) => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11)
         => GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => 
        GND_net_1, A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, 
        A_DIN(6) => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4)
         => GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => 
        GND_net_1, A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, 
        A_ADDR(13) => b9_v_mzCDYXs(11), A_ADDR(12) => 
        b9_v_mzCDYXs(10), A_ADDR(11) => b9_v_mzCDYXs(9), 
        A_ADDR(10) => b9_v_mzCDYXs(8), A_ADDR(9) => 
        b9_v_mzCDYXs(7), A_ADDR(8) => b9_v_mzCDYXs(6), A_ADDR(7)
         => b9_v_mzCDYXs(5), A_ADDR(6) => b9_v_mzCDYXs(4), 
        A_ADDR(5) => b9_v_mzCDYXs(3), A_ADDR(4) => 
        b9_v_mzCDYXs(2), A_ADDR(3) => b9_v_mzCDYXs(1), A_ADDR(2)
         => b9_v_mzCDYXs(0), A_ADDR(1) => GND_net_1, A_ADDR(0)
         => GND_net_1, A_WEN(1) => GND_net_1, A_WEN(0) => 
        GND_net_1, B_CLK => CommsFPGA_CCC_0_GL0, B_DOUT_CLK => 
        VCC_net_1, B_ARST_N => VCC_net_1, B_DOUT_EN => VCC_net_1, 
        B_BLK(2) => VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0)
         => VCC_net_1, B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N
         => VCC_net_1, B_DIN(17) => GND_net_1, B_DIN(16) => 
        GND_net_1, B_DIN(15) => GND_net_1, B_DIN(14) => GND_net_1, 
        B_DIN(13) => GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11)
         => GND_net_1, B_DIN(10) => GND_net_1, B_DIN(9) => 
        GND_net_1, B_DIN(8) => GND_net_1, B_DIN(7) => GND_net_1, 
        B_DIN(6) => GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4)
         => GND_net_1, B_DIN(3) => b11_OFWNT9L_8tZ(167), B_DIN(2)
         => b11_OFWNT9L_8tZ(166), B_DIN(1) => 
        b11_OFWNT9L_8tZ(165), B_DIN(0) => b11_OFWNT9L_8tZ(164), 
        B_ADDR(13) => b12_2_St6KCa_jHv(11), B_ADDR(12) => 
        b12_2_St6KCa_jHv(10), B_ADDR(11) => b12_2_St6KCa_jHv(9), 
        B_ADDR(10) => b12_2_St6KCa_jHv(8), B_ADDR(9) => 
        b12_2_St6KCa_jHv(7), B_ADDR(8) => b12_2_St6KCa_jHv(6), 
        B_ADDR(7) => b12_2_St6KCa_jHv(5), B_ADDR(6) => 
        b12_2_St6KCa_jHv(4), B_ADDR(5) => b12_2_St6KCa_jHv(3), 
        B_ADDR(4) => b12_2_St6KCa_jHv(2), B_ADDR(3) => 
        b12_2_St6KCa_jHv(1), B_ADDR(2) => b12_2_St6KCa_jHv(0), 
        B_ADDR(1) => GND_net_1, B_ADDR(0) => GND_net_1, B_WEN(1)
         => GND_net_1, B_WEN(0) => b4_2o_z, A_EN => VCC_net_1, 
        A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => GND_net_1, 
        A_WIDTH(1) => VCC_net_1, A_WIDTH(0) => GND_net_1, A_WMODE
         => VCC_net_1, B_EN => VCC_net_1, B_DOUT_LAT => VCC_net_1, 
        B_WIDTH(2) => GND_net_1, B_WIDTH(1) => VCC_net_1, 
        B_WIDTH(0) => GND_net_1, B_WMODE => VCC_net_1, SII_LOCK
         => GND_net_1);
    
    b3_SoW_b3_SoW_0_14 : RAM1K18
      port map(A_DOUT(17) => nc975, A_DOUT(16) => nc697, 
        A_DOUT(15) => nc24, A_DOUT(14) => nc848, A_DOUT(13) => 
        nc943, A_DOUT(12) => nc911, A_DOUT(11) => nc900, 
        A_DOUT(10) => nc221, A_DOUT(9) => nc125, A_DOUT(8) => 
        nc183, A_DOUT(7) => nc139, A_DOUT(6) => nc979, A_DOUT(5)
         => nc361, A_DOUT(4) => nc41, A_DOUT(3) => b7_vFW_PlM(59), 
        A_DOUT(2) => b7_vFW_PlM(58), A_DOUT(1) => b7_vFW_PlM(57), 
        A_DOUT(0) => b7_vFW_PlM(56), B_DOUT(17) => nc1056, 
        B_DOUT(16) => nc293, B_DOUT(15) => nc910, B_DOUT(14) => 
        nc736, B_DOUT(13) => nc724, B_DOUT(12) => nc171, 
        B_DOUT(11) => nc320, B_DOUT(10) => nc394, B_DOUT(9) => 
        nc177, B_DOUT(8) => nc407, B_DOUT(7) => nc654, B_DOUT(6)
         => nc464, B_DOUT(5) => nc742, B_DOUT(4) => nc279, 
        B_DOUT(3) => nc1062, B_DOUT(2) => nc1064, B_DOUT(1) => 
        nc417, B_DOUT(0) => nc153, BUSY => OPEN, A_CLK => 
        IICE_comm2iice_0, A_DOUT_CLK => VCC_net_1, A_ARST_N => 
        VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2) => VCC_net_1, 
        A_BLK(1) => VCC_net_1, A_BLK(0) => VCC_net_1, 
        A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => VCC_net_1, 
        A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, A_DIN(15)
         => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13) => 
        GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => GND_net_1, 
        A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, A_DIN(8)
         => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6) => 
        GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => GND_net_1, 
        A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, A_DIN(1)
         => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13) => 
        b9_v_mzCDYXs(11), A_ADDR(12) => b9_v_mzCDYXs(10), 
        A_ADDR(11) => b9_v_mzCDYXs(9), A_ADDR(10) => 
        b9_v_mzCDYXs(8), A_ADDR(9) => b9_v_mzCDYXs(7), A_ADDR(8)
         => b9_v_mzCDYXs(6), A_ADDR(7) => b9_v_mzCDYXs(5), 
        A_ADDR(6) => b9_v_mzCDYXs(4), A_ADDR(5) => 
        b9_v_mzCDYXs(3), A_ADDR(4) => b9_v_mzCDYXs(2), A_ADDR(3)
         => b9_v_mzCDYXs(1), A_ADDR(2) => b9_v_mzCDYXs(0), 
        A_ADDR(1) => GND_net_1, A_ADDR(0) => GND_net_1, A_WEN(1)
         => GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        VCC_net_1, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => VCC_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => b11_OFWNT9L_8tZ(59), B_DIN(2) => 
        b11_OFWNT9L_8tZ(58), B_DIN(1) => b11_OFWNT9L_8tZ(57), 
        B_DIN(0) => b11_OFWNT9L_8tZ(56), B_ADDR(13) => 
        b12_2_St6KCa_jHv(11), B_ADDR(12) => b12_2_St6KCa_jHv(10), 
        B_ADDR(11) => b12_2_St6KCa_jHv(9), B_ADDR(10) => 
        b12_2_St6KCa_jHv(8), B_ADDR(9) => b12_2_St6KCa_jHv(7), 
        B_ADDR(8) => b12_2_St6KCa_jHv(6), B_ADDR(7) => 
        b12_2_St6KCa_jHv(5), B_ADDR(6) => b12_2_St6KCa_jHv(4), 
        B_ADDR(5) => b12_2_St6KCa_jHv(3), B_ADDR(4) => 
        b12_2_St6KCa_jHv(2), B_ADDR(3) => b12_2_St6KCa_jHv(1), 
        B_ADDR(2) => b12_2_St6KCa_jHv(0), B_ADDR(1) => GND_net_1, 
        B_ADDR(0) => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0)
         => b4_2o_z, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => GND_net_1, A_WMODE => VCC_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        GND_net_1, B_WMODE => VCC_net_1, SII_LOCK => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b19_nczQ_DYg_YFaRM_oUoP_32s_1s_x_0 is

    port( IICE_comm2iice_5 : in    std_logic;
          IICE_comm2iice_3 : in    std_logic;
          IICE_comm2iice_0 : in    std_logic;
          IICE_comm2iice_4 : in    std_logic;
          N_1261_i         : out   std_logic;
          ttdo             : in    std_logic;
          b7_yYh03wy5      : in    std_logic;
          b7_yYh03wy4      : in    std_logic
        );

end b19_nczQ_DYg_YFaRM_oUoP_32s_1s_x_0;

architecture DEF_ARCH of b19_nczQ_DYg_YFaRM_oUoP_32s_1s_x_0 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \b13_PLF_2grFt_FH9[24]\, VCC_net_1, 
        \b13_PLF_2grFt_FH9_5[24]\, N_26, GND_net_1, 
        \b13_PLF_2grFt_FH9[25]\, \b13_PLF_2grFt_FH9_5[25]\, 
        \b13_PLF_2grFt_FH9[26]\, \b13_PLF_2grFt_FH9_5[26]\, 
        \b13_PLF_2grFt_FH9[27]\, \b13_PLF_2grFt_FH9_5[27]\, 
        \b13_PLF_2grFt_FH9[28]\, \b13_PLF_2grFt_FH9_5[28]\, 
        \b13_PLF_2grFt_FH9[29]\, \b13_PLF_2grFt_FH9_5[29]\, 
        \b13_PLF_2grFt_FH9[30]\, \b13_PLF_2grFt_FH9_5[30]\, 
        \b13_PLF_2grFt_FH9[31]\, \b13_PLF_2grFt_FH9[9]\, 
        \b13_PLF_2grFt_FH9_5[9]\, \b13_PLF_2grFt_FH9[10]\, 
        \b13_PLF_2grFt_FH9_5[10]\, \b13_PLF_2grFt_FH9[11]\, 
        \b13_PLF_2grFt_FH9_5[11]\, \b13_PLF_2grFt_FH9[12]\, 
        \b13_PLF_2grFt_FH9_5[12]\, \b13_PLF_2grFt_FH9[13]\, 
        \b13_PLF_2grFt_FH9_5[13]\, \b13_PLF_2grFt_FH9[14]\, 
        \b13_PLF_2grFt_FH9_5[14]\, \b13_PLF_2grFt_FH9[15]\, 
        \b13_PLF_2grFt_FH9_5[15]\, \b13_PLF_2grFt_FH9[16]\, 
        \b13_PLF_2grFt_FH9_5[16]\, \b13_PLF_2grFt_FH9[17]\, 
        \b13_PLF_2grFt_FH9_5[17]\, \b13_PLF_2grFt_FH9[18]\, 
        \b13_PLF_2grFt_FH9_5[18]\, \b13_PLF_2grFt_FH9[19]\, 
        \b13_PLF_2grFt_FH9_5[19]\, \b13_PLF_2grFt_FH9[20]\, 
        \b13_PLF_2grFt_FH9_5[20]\, \b13_PLF_2grFt_FH9[21]\, 
        \b13_PLF_2grFt_FH9_5[21]\, \b13_PLF_2grFt_FH9[22]\, 
        \b13_PLF_2grFt_FH9_5[22]\, \b13_PLF_2grFt_FH9[23]\, 
        \b13_PLF_2grFt_FH9_5[23]\, b4_ycsM, 
        \b13_PLF_2grFt_FH9_5[0]\, \b13_PLF_2grFt_FH9[1]\, 
        \b13_PLF_2grFt_FH9_5[1]\, \b13_PLF_2grFt_FH9[2]\, 
        \b13_PLF_2grFt_FH9_5[2]\, \b13_PLF_2grFt_FH9[3]\, 
        \b13_PLF_2grFt_FH9_5[3]\, \b13_PLF_2grFt_FH9[4]\, 
        \b13_PLF_2grFt_FH9_5[4]\, \b13_PLF_2grFt_FH9[5]\, 
        \b13_PLF_2grFt_FH9_5[5]\, \b13_PLF_2grFt_FH9[6]\, 
        \b13_PLF_2grFt_FH9_5[6]\, \b13_PLF_2grFt_FH9[7]\, 
        \b13_PLF_2grFt_FH9_5[7]\, \b13_PLF_2grFt_FH9[8]\, 
        \b13_PLF_2grFt_FH9_5[8]\ : std_logic;

begin 


    \genblk1.b13_PLF_2grFt_FH9[2]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[2]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[2]\);
    
    \genblk1.b13_PLF_2grFt_FH9_5[22]\ : CFG2
      generic map(INIT => x"E")

      port map(A => IICE_comm2iice_3, B => 
        \b13_PLF_2grFt_FH9[23]\, Y => \b13_PLF_2grFt_FH9_5[22]\);
    
    \genblk1.b13_PLF_2grFt_FH9_5[26]\ : CFG2
      generic map(INIT => x"4")

      port map(A => IICE_comm2iice_3, B => 
        \b13_PLF_2grFt_FH9[27]\, Y => \b13_PLF_2grFt_FH9_5[26]\);
    
    \genblk1.b13_PLF_2grFt_FH9_5[5]\ : CFG2
      generic map(INIT => x"E")

      port map(A => IICE_comm2iice_3, B => \b13_PLF_2grFt_FH9[6]\, 
        Y => \b13_PLF_2grFt_FH9_5[5]\);
    
    \genblk1.b13_PLF_2grFt_FH9[5]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[5]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[5]\);
    
    \genblk1.b13_PLF_2grFt_FH9[16]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[16]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[16]\);
    
    \genblk1.b13_PLF_2grFt_FH9_5[3]\ : CFG2
      generic map(INIT => x"E")

      port map(A => IICE_comm2iice_3, B => \b13_PLF_2grFt_FH9[4]\, 
        Y => \b13_PLF_2grFt_FH9_5[3]\);
    
    \genblk1.b13_PLF_2grFt_FH9[10]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[10]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[10]\);
    
    \genblk1.b13_PLF_2grFt_FH9_RNI8O1S[0]\ : CFG4
      generic map(INIT => x"E2C0")

      port map(A => b7_yYh03wy4, B => b7_yYh03wy5, C => ttdo, D
         => b4_ycsM, Y => N_1261_i);
    
    \genblk1.b13_PLF_2grFt_FH9_5[25]\ : CFG2
      generic map(INIT => x"E")

      port map(A => IICE_comm2iice_3, B => 
        \b13_PLF_2grFt_FH9[26]\, Y => \b13_PLF_2grFt_FH9_5[25]\);
    
    \genblk1.b13_PLF_2grFt_FH9[23]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[23]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[23]\);
    
    \genblk1.b13_PLF_2grFt_FH9[0]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[0]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => b4_ycsM);
    
    \genblk1.b13_PLF_2grFt_FH9_5[30]\ : CFG2
      generic map(INIT => x"E")

      port map(A => IICE_comm2iice_3, B => 
        \b13_PLF_2grFt_FH9[31]\, Y => \b13_PLF_2grFt_FH9_5[30]\);
    
    \genblk1.b13_PLF_2grFt_FH9_5[20]\ : CFG2
      generic map(INIT => x"E")

      port map(A => IICE_comm2iice_3, B => 
        \b13_PLF_2grFt_FH9[21]\, Y => \b13_PLF_2grFt_FH9_5[20]\);
    
    \genblk1.b13_PLF_2grFt_FH9[11]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[11]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[11]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \genblk1.b13_PLF_2grFt_FH9_5[21]\ : CFG2
      generic map(INIT => x"E")

      port map(A => IICE_comm2iice_3, B => 
        \b13_PLF_2grFt_FH9[22]\, Y => \b13_PLF_2grFt_FH9_5[21]\);
    
    \genblk1.b13_PLF_2grFt_FH9_5[18]\ : CFG2
      generic map(INIT => x"E")

      port map(A => IICE_comm2iice_3, B => 
        \b13_PLF_2grFt_FH9[19]\, Y => \b13_PLF_2grFt_FH9_5[18]\);
    
    \genblk1.b13_PLF_2grFt_FH9_5[1]\ : CFG2
      generic map(INIT => x"E")

      port map(A => IICE_comm2iice_3, B => \b13_PLF_2grFt_FH9[2]\, 
        Y => \b13_PLF_2grFt_FH9_5[1]\);
    
    \genblk1.b13_PLF_2grFt_FH9[12]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[12]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[12]\);
    
    \genblk1.b13_PLF_2grFt_FH9_5[17]\ : CFG2
      generic map(INIT => x"E")

      port map(A => IICE_comm2iice_3, B => 
        \b13_PLF_2grFt_FH9[18]\, Y => \b13_PLF_2grFt_FH9_5[17]\);
    
    \genblk1.b13_PLF_2grFt_FH9_5[4]\ : CFG2
      generic map(INIT => x"E")

      port map(A => IICE_comm2iice_3, B => \b13_PLF_2grFt_FH9[5]\, 
        Y => \b13_PLF_2grFt_FH9_5[4]\);
    
    \genblk1.b13_PLF_2grFt_FH9[17]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[17]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[17]\);
    
    \genblk1.b13_PLF_2grFt_FH9[26]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[26]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[26]\);
    
    \genblk1.b13_PLF_2grFt_FH9[20]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[20]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[20]\);
    
    \genblk1.b13_PLF_2grFt_FH9_5[24]\ : CFG2
      generic map(INIT => x"4")

      port map(A => IICE_comm2iice_3, B => 
        \b13_PLF_2grFt_FH9[25]\, Y => \b13_PLF_2grFt_FH9_5[24]\);
    
    \genblk1.b13_PLF_2grFt_FH9_5[13]\ : CFG2
      generic map(INIT => x"4")

      port map(A => IICE_comm2iice_3, B => 
        \b13_PLF_2grFt_FH9[14]\, Y => \b13_PLF_2grFt_FH9_5[13]\);
    
    \genblk1.b13_PLF_2grFt_FH9[14]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[14]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[14]\);
    
    \genblk1.b13_PLF_2grFt_FH9_5[29]\ : CFG2
      generic map(INIT => x"4")

      port map(A => IICE_comm2iice_3, B => 
        \b13_PLF_2grFt_FH9[30]\, Y => \b13_PLF_2grFt_FH9_5[29]\);
    
    \genblk1.b13_PLF_2grFt_FH9[6]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[6]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[6]\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \genblk1.b13_PLF_2grFt_FH9[21]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[21]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[21]\);
    
    \genblk1.b13_PLF_2grFt_FH9_5[0]\ : CFG2
      generic map(INIT => x"4")

      port map(A => IICE_comm2iice_3, B => \b13_PLF_2grFt_FH9[1]\, 
        Y => \b13_PLF_2grFt_FH9_5[0]\);
    
    \genblk1.b13_PLF_2grFt_FH9[22]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[22]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[22]\);
    
    \genblk1.b13_PLF_2grFt_FH9[18]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[18]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[18]\);
    
    \genblk1.b13_PLF_2grFt_FH9_5[12]\ : CFG2
      generic map(INIT => x"4")

      port map(A => IICE_comm2iice_3, B => 
        \b13_PLF_2grFt_FH9[13]\, Y => \b13_PLF_2grFt_FH9_5[12]\);
    
    \genblk1.b13_PLF_2grFt_FH9_5[16]\ : CFG2
      generic map(INIT => x"4")

      port map(A => IICE_comm2iice_3, B => 
        \b13_PLF_2grFt_FH9[17]\, Y => \b13_PLF_2grFt_FH9_5[16]\);
    
    \genblk1.b13_PLF_2grFt_FH9[9]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[9]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[9]\);
    
    \genblk1.b13_PLF_2grFt_FH9[4]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[4]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[4]\);
    
    \genblk1.b13_PLF_2grFt_FH9[27]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[27]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[27]\);
    
    \genblk1.b13_PLF_2grFt_FH9[30]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[30]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[30]\);
    
    \genblk1.b13_PLF_2grFt_FH9_5[8]\ : CFG2
      generic map(INIT => x"4")

      port map(A => IICE_comm2iice_3, B => \b13_PLF_2grFt_FH9[9]\, 
        Y => \b13_PLF_2grFt_FH9_5[8]\);
    
    \genblk1.b13_PLF_2grFt_FH9[24]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[24]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[24]\);
    
    \genblk1.b13_PLF_2grFt_FH9_5[15]\ : CFG2
      generic map(INIT => x"E")

      port map(A => IICE_comm2iice_3, B => 
        \b13_PLF_2grFt_FH9[16]\, Y => \b13_PLF_2grFt_FH9_5[15]\);
    
    \genblk1.b13_PLF_2grFt_FH9[15]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[15]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[15]\);
    
    \genblk1.b13_PLF_2grFt_FH9_5[10]\ : CFG2
      generic map(INIT => x"4")

      port map(A => IICE_comm2iice_3, B => 
        \b13_PLF_2grFt_FH9[11]\, Y => \b13_PLF_2grFt_FH9_5[10]\);
    
    \genblk1.b13_PLF_2grFt_FH9[3]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[3]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[3]\);
    
    \genblk1.b13_PLF_2grFt_FH9[31]\ : SLE
      port map(D => IICE_comm2iice_3, CLK => IICE_comm2iice_5, EN
         => N_26, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b13_PLF_2grFt_FH9[31]\);
    
    \genblk1.b13_PLF_2grFt_FH9_5[9]\ : CFG2
      generic map(INIT => x"E")

      port map(A => IICE_comm2iice_3, B => 
        \b13_PLF_2grFt_FH9[10]\, Y => \b13_PLF_2grFt_FH9_5[9]\);
    
    \genblk1.b13_PLF_2grFt_FH9[1]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[1]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[1]\);
    
    \genblk1.b13_PLF_2grFt_FH9_5[11]\ : CFG2
      generic map(INIT => x"E")

      port map(A => IICE_comm2iice_3, B => 
        \b13_PLF_2grFt_FH9[12]\, Y => \b13_PLF_2grFt_FH9_5[11]\);
    
    \genblk1.b13_PLF_2grFt_FH9[7]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[7]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[7]\);
    
    \genblk1.b13_PLF_2grFt_FH9[19]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[19]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[19]\);
    
    \genblk1.b13_PLF_2grFt_FH9_5[6]\ : CFG2
      generic map(INIT => x"E")

      port map(A => IICE_comm2iice_3, B => \b13_PLF_2grFt_FH9[7]\, 
        Y => \b13_PLF_2grFt_FH9_5[6]\);
    
    \genblk1.b13_PLF_2grFt_FH9_5[7]\ : CFG2
      generic map(INIT => x"E")

      port map(A => IICE_comm2iice_3, B => \b13_PLF_2grFt_FH9[8]\, 
        Y => \b13_PLF_2grFt_FH9_5[7]\);
    
    \genblk1.b13_PLF_2grFt_FH9[28]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[28]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[28]\);
    
    \genblk1.b13_PLF_2grFt_FH9_5[28]\ : CFG2
      generic map(INIT => x"4")

      port map(A => IICE_comm2iice_3, B => 
        \b13_PLF_2grFt_FH9[29]\, Y => \b13_PLF_2grFt_FH9_5[28]\);
    
    \genblk1.b13_PLF_2grFt_FH9[8]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[8]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[8]\);
    
    \genblk1.b13_PLF_2grFt_FH9_5[27]\ : CFG2
      generic map(INIT => x"E")

      port map(A => IICE_comm2iice_3, B => 
        \b13_PLF_2grFt_FH9[28]\, Y => \b13_PLF_2grFt_FH9_5[27]\);
    
    un1_b13_PLF_2grFt_FH911_i_a2 : CFG4
      generic map(INIT => x"A080")

      port map(A => IICE_comm2iice_0, B => IICE_comm2iice_3, C
         => b7_yYh03wy4, D => IICE_comm2iice_4, Y => N_26);
    
    \genblk1.b13_PLF_2grFt_FH9_5[14]\ : CFG2
      generic map(INIT => x"E")

      port map(A => IICE_comm2iice_3, B => 
        \b13_PLF_2grFt_FH9[15]\, Y => \b13_PLF_2grFt_FH9_5[14]\);
    
    \genblk1.b13_PLF_2grFt_FH9_5[2]\ : CFG2
      generic map(INIT => x"E")

      port map(A => IICE_comm2iice_3, B => \b13_PLF_2grFt_FH9[3]\, 
        Y => \b13_PLF_2grFt_FH9_5[2]\);
    
    \genblk1.b13_PLF_2grFt_FH9[25]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[25]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[25]\);
    
    \genblk1.b13_PLF_2grFt_FH9_5[19]\ : CFG2
      generic map(INIT => x"E")

      port map(A => IICE_comm2iice_3, B => 
        \b13_PLF_2grFt_FH9[20]\, Y => \b13_PLF_2grFt_FH9_5[19]\);
    
    \genblk1.b13_PLF_2grFt_FH9_5[23]\ : CFG2
      generic map(INIT => x"E")

      port map(A => IICE_comm2iice_3, B => 
        \b13_PLF_2grFt_FH9[24]\, Y => \b13_PLF_2grFt_FH9_5[23]\);
    
    \genblk1.b13_PLF_2grFt_FH9[29]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[29]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[29]\);
    
    \genblk1.b13_PLF_2grFt_FH9[13]\ : SLE
      port map(D => \b13_PLF_2grFt_FH9_5[13]\, CLK => 
        IICE_comm2iice_5, EN => N_26, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b13_PLF_2grFt_FH9[13]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b11_SoWyP0zEFKY_Z2_x_0 is

    port( mdiclink_reg        : in    std_logic_vector(167 downto 0);
          b11_OFWNT9L_8tZ     : out   std_logic_vector(167 downto 0);
          N_145_i             : in    std_logic;
          b4_2o_z             : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic
        );

end b11_SoWyP0zEFKY_Z2_x_0;

architecture DEF_ARCH of b11_SoWyP0zEFKY_Z2_x_0 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;

begin 


    \genblk2.b5_oRB_C[72]\ : SLE
      port map(D => mdiclink_reg(95), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(72));
    
    \genblk2.b5_oRB_C[164]\ : SLE
      port map(D => mdiclink_reg(3), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(164));
    
    \genblk2.b5_oRB_C[61]\ : SLE
      port map(D => mdiclink_reg(106), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(61));
    
    \genblk2.b5_oRB_C[131]\ : SLE
      port map(D => mdiclink_reg(36), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(131));
    
    \genblk2.b5_oRB_C[82]\ : SLE
      port map(D => mdiclink_reg(85), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(82));
    
    \genblk2.b5_oRB_C[122]\ : SLE
      port map(D => mdiclink_reg(45), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(122));
    
    \genblk2.b5_oRB_C[17]\ : SLE
      port map(D => mdiclink_reg(150), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(17));
    
    \genblk2.b5_oRB_C[18]\ : SLE
      port map(D => mdiclink_reg(149), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(18));
    
    \genblk2.b5_oRB_C[66]\ : SLE
      port map(D => mdiclink_reg(101), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(66));
    
    \genblk2.b5_oRB_C[137]\ : SLE
      port map(D => mdiclink_reg(30), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(137));
    
    \genblk2.b5_oRB_C[105]\ : SLE
      port map(D => mdiclink_reg(62), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(105));
    
    \genblk2.b5_oRB_C[121]\ : SLE
      port map(D => mdiclink_reg(46), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(121));
    
    \genblk2.b5_oRB_C[166]\ : SLE
      port map(D => mdiclink_reg(1), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(166));
    
    \genblk2.b5_oRB_C[20]\ : SLE
      port map(D => mdiclink_reg(147), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(20));
    
    \genblk2.b5_oRB_C[43]\ : SLE
      port map(D => mdiclink_reg(124), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(43));
    
    \genblk2.b5_oRB_C[93]\ : SLE
      port map(D => mdiclink_reg(74), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(93));
    
    \genblk2.b5_oRB_C[11]\ : SLE
      port map(D => mdiclink_reg(156), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(11));
    
    \genblk2.b5_oRB_C[127]\ : SLE
      port map(D => mdiclink_reg(40), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(127));
    
    \genblk2.b5_oRB_C[30]\ : SLE
      port map(D => mdiclink_reg(137), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(30));
    
    \genblk2.b5_oRB_C[16]\ : SLE
      port map(D => mdiclink_reg(151), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(16));
    
    \genblk2.b5_oRB_C[45]\ : SLE
      port map(D => mdiclink_reg(122), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(45));
    
    \genblk2.b5_oRB_C[95]\ : SLE
      port map(D => mdiclink_reg(72), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(95));
    
    \genblk2.b5_oRB_C[70]\ : SLE
      port map(D => mdiclink_reg(97), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(70));
    
    \genblk2.b5_oRB_C[5]\ : SLE
      port map(D => mdiclink_reg(162), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(5));
    
    \genblk2.b5_oRB_C[80]\ : SLE
      port map(D => mdiclink_reg(87), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(80));
    
    \genblk2.b5_oRB_C[0]\ : SLE
      port map(D => mdiclink_reg(167), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(0));
    
    \genblk2.b5_oRB_C[104]\ : SLE
      port map(D => mdiclink_reg(63), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(104));
    
    \genblk2.b5_oRB_C[57]\ : SLE
      port map(D => mdiclink_reg(110), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(57));
    
    \genblk2.b5_oRB_C[58]\ : SLE
      port map(D => mdiclink_reg(109), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(58));
    
    \genblk2.b5_oRB_C[63]\ : SLE
      port map(D => mdiclink_reg(104), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(63));
    
    \genblk2.b5_oRB_C[106]\ : SLE
      port map(D => mdiclink_reg(61), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(106));
    
    \genblk2.b5_oRB_C[65]\ : SLE
      port map(D => mdiclink_reg(102), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(65));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \genblk2.b5_oRB_C[51]\ : SLE
      port map(D => mdiclink_reg(116), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(51));
    
    \genblk2.b5_oRB_C[115]\ : SLE
      port map(D => mdiclink_reg(52), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(115));
    
    \genblk2.b5_oRB_C[13]\ : SLE
      port map(D => mdiclink_reg(154), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(13));
    
    \genblk2.b5_oRB_C[56]\ : SLE
      port map(D => mdiclink_reg(111), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(56));
    
    \genblk2.b5_oRB_C[160]\ : SLE
      port map(D => mdiclink_reg(7), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(160));
    
    \genblk2.b5_oRB_C[155]\ : SLE
      port map(D => mdiclink_reg(12), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(155));
    
    \genblk2.b5_oRB_C[163]\ : SLE
      port map(D => mdiclink_reg(4), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(163));
    
    \genblk2.b5_oRB_C[44]\ : SLE
      port map(D => mdiclink_reg(123), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(44));
    
    \genblk2.b5_oRB_C[94]\ : SLE
      port map(D => mdiclink_reg(73), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(94));
    
    \genblk2.b5_oRB_C[15]\ : SLE
      port map(D => mdiclink_reg(152), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(15));
    
    \genblk2.b5_oRB_C[3]\ : SLE
      port map(D => mdiclink_reg(164), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(3));
    
    \genblk2.b5_oRB_C[114]\ : SLE
      port map(D => mdiclink_reg(53), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(114));
    
    \genblk2.b5_oRB_C[108]\ : SLE
      port map(D => mdiclink_reg(59), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(108));
    
    \genblk2.b5_oRB_C[154]\ : SLE
      port map(D => mdiclink_reg(13), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(154));
    
    \genblk2.b5_oRB_C[53]\ : SLE
      port map(D => mdiclink_reg(114), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(53));
    
    \genblk2.b5_oRB_C[64]\ : SLE
      port map(D => mdiclink_reg(103), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(64));
    
    \genblk2.b5_oRB_C[116]\ : SLE
      port map(D => mdiclink_reg(51), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(116));
    
    \genblk2.b5_oRB_C[49]\ : SLE
      port map(D => mdiclink_reg(118), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(49));
    
    \genblk2.b5_oRB_C[99]\ : SLE
      port map(D => mdiclink_reg(68), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(99));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \genblk2.b5_oRB_C[100]\ : SLE
      port map(D => mdiclink_reg(67), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(100));
    
    \genblk2.b5_oRB_C[103]\ : SLE
      port map(D => mdiclink_reg(64), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(103));
    
    \genblk2.b5_oRB_C[156]\ : SLE
      port map(D => mdiclink_reg(11), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(156));
    
    \genblk2.b5_oRB_C[145]\ : SLE
      port map(D => mdiclink_reg(22), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(145));
    
    \genblk2.b5_oRB_C[55]\ : SLE
      port map(D => mdiclink_reg(112), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(55));
    
    \genblk2.b5_oRB_C[162]\ : SLE
      port map(D => mdiclink_reg(5), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(162));
    
    \genblk2.b5_oRB_C[27]\ : SLE
      port map(D => mdiclink_reg(140), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(27));
    
    \genblk2.b5_oRB_C[28]\ : SLE
      port map(D => mdiclink_reg(139), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(28));
    
    \genblk2.b5_oRB_C[14]\ : SLE
      port map(D => mdiclink_reg(153), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(14));
    
    \genblk2.b5_oRB_C[37]\ : SLE
      port map(D => mdiclink_reg(130), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(37));
    
    \genblk2.b5_oRB_C[161]\ : SLE
      port map(D => mdiclink_reg(6), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(161));
    
    \genblk2.b5_oRB_C[38]\ : SLE
      port map(D => mdiclink_reg(129), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(38));
    
    \genblk2.b5_oRB_C[69]\ : SLE
      port map(D => mdiclink_reg(98), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(69));
    
    \genblk2.b5_oRB_C[109]\ : SLE
      port map(D => mdiclink_reg(58), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(109));
    
    \genblk2.b5_oRB_C[1]\ : SLE
      port map(D => mdiclink_reg(166), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(1));
    
    \genblk2.b5_oRB_C[21]\ : SLE
      port map(D => mdiclink_reg(146), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(21));
    
    \genblk2.b5_oRB_C[167]\ : SLE
      port map(D => mdiclink_reg(0), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(167));
    
    \genblk2.b5_oRB_C[77]\ : SLE
      port map(D => mdiclink_reg(90), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(77));
    
    \genblk2.b5_oRB_C[144]\ : SLE
      port map(D => mdiclink_reg(23), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(144));
    
    \genblk2.b5_oRB_C[78]\ : SLE
      port map(D => mdiclink_reg(89), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(78));
    
    \genblk2.b5_oRB_C[87]\ : SLE
      port map(D => mdiclink_reg(80), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(87));
    
    \genblk2.b5_oRB_C[88]\ : SLE
      port map(D => mdiclink_reg(79), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(88));
    
    \genblk2.b5_oRB_C[42]\ : SLE
      port map(D => mdiclink_reg(125), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(42));
    
    \genblk2.b5_oRB_C[92]\ : SLE
      port map(D => mdiclink_reg(75), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(92));
    
    \genblk2.b5_oRB_C[118]\ : SLE
      port map(D => mdiclink_reg(49), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(118));
    
    \genblk2.b5_oRB_C[26]\ : SLE
      port map(D => mdiclink_reg(141), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(26));
    
    \genblk2.b5_oRB_C[31]\ : SLE
      port map(D => mdiclink_reg(136), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(31));
    
    \genblk2.b5_oRB_C[158]\ : SLE
      port map(D => mdiclink_reg(9), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(158));
    
    \genblk2.b5_oRB_C[36]\ : SLE
      port map(D => mdiclink_reg(131), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(36));
    
    \genblk2.b5_oRB_C[146]\ : SLE
      port map(D => mdiclink_reg(21), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(146));
    
    \genblk2.b5_oRB_C[19]\ : SLE
      port map(D => mdiclink_reg(148), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(19));
    
    \genblk2.b5_oRB_C[9]\ : SLE
      port map(D => mdiclink_reg(158), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(9));
    
    \genblk2.b5_oRB_C[71]\ : SLE
      port map(D => mdiclink_reg(96), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(71));
    
    \genblk2.b5_oRB_C[102]\ : SLE
      port map(D => mdiclink_reg(65), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(102));
    
    \genblk2.b5_oRB_C[54]\ : SLE
      port map(D => mdiclink_reg(113), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(54));
    
    \genblk2.b5_oRB_C[81]\ : SLE
      port map(D => mdiclink_reg(86), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(81));
    
    \genblk2.b5_oRB_C[110]\ : SLE
      port map(D => mdiclink_reg(57), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(110));
    
    \genblk2.b5_oRB_C[113]\ : SLE
      port map(D => mdiclink_reg(54), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(113));
    
    \genblk2.b5_oRB_C[76]\ : SLE
      port map(D => mdiclink_reg(91), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(76));
    
    \genblk2.b5_oRB_C[86]\ : SLE
      port map(D => mdiclink_reg(81), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(86));
    
    \genblk2.b5_oRB_C[150]\ : SLE
      port map(D => mdiclink_reg(17), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(150));
    
    \genblk2.b5_oRB_C[153]\ : SLE
      port map(D => mdiclink_reg(14), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(153));
    
    \genblk2.b5_oRB_C[101]\ : SLE
      port map(D => mdiclink_reg(66), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(101));
    
    \genblk2.b5_oRB_C[62]\ : SLE
      port map(D => mdiclink_reg(105), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(62));
    
    \genblk2.b5_oRB_C[135]\ : SLE
      port map(D => mdiclink_reg(32), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(135));
    
    \genblk2.b5_oRB_C[40]\ : SLE
      port map(D => mdiclink_reg(127), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(40));
    
    \genblk2.b5_oRB_C[107]\ : SLE
      port map(D => mdiclink_reg(60), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(107));
    
    \genblk2.b5_oRB_C[90]\ : SLE
      port map(D => mdiclink_reg(77), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(90));
    
    \genblk2.b5_oRB_C[23]\ : SLE
      port map(D => mdiclink_reg(144), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(23));
    
    \genblk2.b5_oRB_C[125]\ : SLE
      port map(D => mdiclink_reg(42), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(125));
    
    \genblk2.b5_oRB_C[119]\ : SLE
      port map(D => mdiclink_reg(48), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(119));
    
    \genblk2.b5_oRB_C[33]\ : SLE
      port map(D => mdiclink_reg(134), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(33));
    
    \genblk2.b5_oRB_C[59]\ : SLE
      port map(D => mdiclink_reg(108), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(59));
    
    \genblk2.b5_oRB_C[12]\ : SLE
      port map(D => mdiclink_reg(155), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(12));
    
    \genblk2.b5_oRB_C[159]\ : SLE
      port map(D => mdiclink_reg(8), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(159));
    
    \genblk2.b5_oRB_C[7]\ : SLE
      port map(D => mdiclink_reg(160), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(7));
    
    \genblk2.b5_oRB_C[25]\ : SLE
      port map(D => mdiclink_reg(142), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(25));
    
    \genblk2.b5_oRB_C[148]\ : SLE
      port map(D => mdiclink_reg(19), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(148));
    
    \genblk2.b5_oRB_C[134]\ : SLE
      port map(D => mdiclink_reg(33), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(134));
    
    \genblk2.b5_oRB_C[73]\ : SLE
      port map(D => mdiclink_reg(94), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(73));
    
    \genblk2.b5_oRB_C[83]\ : SLE
      port map(D => mdiclink_reg(84), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(83));
    
    \genblk2.b5_oRB_C[35]\ : SLE
      port map(D => mdiclink_reg(132), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(35));
    
    \genblk2.b5_oRB_C[60]\ : SLE
      port map(D => mdiclink_reg(107), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(60));
    
    \genblk2.b5_oRB_C[112]\ : SLE
      port map(D => mdiclink_reg(55), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(112));
    
    \genblk2.b5_oRB_C[140]\ : SLE
      port map(D => mdiclink_reg(27), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(140));
    
    \genblk2.b13_oRB_MqCD2_EdR_0_\ : SLE
      port map(D => N_145_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b4_2o_z);
    
    \genblk2.b5_oRB_C[143]\ : SLE
      port map(D => mdiclink_reg(24), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(143));
    
    \genblk2.b5_oRB_C[124]\ : SLE
      port map(D => mdiclink_reg(43), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(124));
    
    \genblk2.b5_oRB_C[75]\ : SLE
      port map(D => mdiclink_reg(92), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(75));
    
    \genblk2.b5_oRB_C[136]\ : SLE
      port map(D => mdiclink_reg(31), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(136));
    
    \genblk2.b5_oRB_C[85]\ : SLE
      port map(D => mdiclink_reg(82), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(85));
    
    \genblk2.b5_oRB_C[152]\ : SLE
      port map(D => mdiclink_reg(15), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(152));
    
    \genblk2.b5_oRB_C[111]\ : SLE
      port map(D => mdiclink_reg(56), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(111));
    
    \genblk2.b5_oRB_C[8]\ : SLE
      port map(D => mdiclink_reg(159), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(8));
    
    \genblk2.b5_oRB_C[2]\ : SLE
      port map(D => mdiclink_reg(165), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(2));
    
    \genblk2.b5_oRB_C[126]\ : SLE
      port map(D => mdiclink_reg(41), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(126));
    
    \genblk2.b5_oRB_C[10]\ : SLE
      port map(D => mdiclink_reg(157), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(10));
    
    \genblk2.b5_oRB_C[52]\ : SLE
      port map(D => mdiclink_reg(115), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(52));
    
    \genblk2.b5_oRB_C[151]\ : SLE
      port map(D => mdiclink_reg(16), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(151));
    
    \genblk2.b5_oRB_C[117]\ : SLE
      port map(D => mdiclink_reg(50), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(117));
    
    \genblk2.b5_oRB_C[149]\ : SLE
      port map(D => mdiclink_reg(18), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(149));
    
    \genblk2.b5_oRB_C[157]\ : SLE
      port map(D => mdiclink_reg(10), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(157));
    
    \genblk2.b5_oRB_C[24]\ : SLE
      port map(D => mdiclink_reg(143), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(24));
    
    \genblk2.b5_oRB_C[34]\ : SLE
      port map(D => mdiclink_reg(133), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(34));
    
    \genblk2.b5_oRB_C[4]\ : SLE
      port map(D => mdiclink_reg(163), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(4));
    
    \genblk2.b5_oRB_C[138]\ : SLE
      port map(D => mdiclink_reg(29), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(138));
    
    \genblk2.b5_oRB_C[142]\ : SLE
      port map(D => mdiclink_reg(25), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(142));
    
    \genblk2.b5_oRB_C[74]\ : SLE
      port map(D => mdiclink_reg(93), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(74));
    
    \genblk2.b5_oRB_C[84]\ : SLE
      port map(D => mdiclink_reg(83), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(84));
    
    \genblk2.b5_oRB_C[50]\ : SLE
      port map(D => mdiclink_reg(117), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(50));
    
    \genblk2.b5_oRB_C[128]\ : SLE
      port map(D => mdiclink_reg(39), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(128));
    
    \genblk2.b5_oRB_C[130]\ : SLE
      port map(D => mdiclink_reg(37), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(130));
    
    \genblk2.b5_oRB_C[141]\ : SLE
      port map(D => mdiclink_reg(26), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(141));
    
    \genblk2.b5_oRB_C[133]\ : SLE
      port map(D => mdiclink_reg(34), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(133));
    
    \genblk2.b5_oRB_C[29]\ : SLE
      port map(D => mdiclink_reg(138), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(29));
    
    \genblk2.b5_oRB_C[147]\ : SLE
      port map(D => mdiclink_reg(20), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(147));
    
    \genblk2.b5_oRB_C[39]\ : SLE
      port map(D => mdiclink_reg(128), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(39));
    
    \genblk2.b5_oRB_C[120]\ : SLE
      port map(D => mdiclink_reg(47), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(120));
    
    \genblk2.b5_oRB_C[123]\ : SLE
      port map(D => mdiclink_reg(44), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(123));
    
    \genblk2.b5_oRB_C[47]\ : SLE
      port map(D => mdiclink_reg(120), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(47));
    
    \genblk2.b5_oRB_C[97]\ : SLE
      port map(D => mdiclink_reg(70), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(97));
    
    \genblk2.b5_oRB_C[48]\ : SLE
      port map(D => mdiclink_reg(119), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(48));
    
    \genblk2.b5_oRB_C[98]\ : SLE
      port map(D => mdiclink_reg(69), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(98));
    
    \genblk2.b5_oRB_C[79]\ : SLE
      port map(D => mdiclink_reg(88), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(79));
    
    \genblk2.b5_oRB_C[89]\ : SLE
      port map(D => mdiclink_reg(78), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(89));
    
    \genblk2.b5_oRB_C[139]\ : SLE
      port map(D => mdiclink_reg(28), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(139));
    
    \genblk2.b5_oRB_C[165]\ : SLE
      port map(D => mdiclink_reg(2), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(165));
    
    \genblk2.b5_oRB_C[6]\ : SLE
      port map(D => mdiclink_reg(161), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(6));
    
    \genblk2.b5_oRB_C[41]\ : SLE
      port map(D => mdiclink_reg(126), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(41));
    
    \genblk2.b5_oRB_C[91]\ : SLE
      port map(D => mdiclink_reg(76), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(91));
    
    \genblk2.b5_oRB_C[129]\ : SLE
      port map(D => mdiclink_reg(38), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(129));
    
    \genblk2.b5_oRB_C[22]\ : SLE
      port map(D => mdiclink_reg(145), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(22));
    
    \genblk2.b5_oRB_C[46]\ : SLE
      port map(D => mdiclink_reg(121), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(46));
    
    \genblk2.b5_oRB_C[96]\ : SLE
      port map(D => mdiclink_reg(71), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(96));
    
    \genblk2.b5_oRB_C[67]\ : SLE
      port map(D => mdiclink_reg(100), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(67));
    
    \genblk2.b5_oRB_C[68]\ : SLE
      port map(D => mdiclink_reg(99), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(68));
    
    \genblk2.b5_oRB_C[32]\ : SLE
      port map(D => mdiclink_reg(135), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(32));
    
    \genblk2.b5_oRB_C[132]\ : SLE
      port map(D => mdiclink_reg(35), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_OFWNT9L_8tZ(132));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b11_OFWNT9s_8tZ_Z3_x is

    port( mdiclink_reg        : in    std_logic_vector(167 downto 0);
          b11_OFWNT9L_8tZ     : out   std_logic_vector(167 downto 0);
          IICE_comm2iice      : in    std_logic_vector(11 downto 0);
          N_145_i             : in    std_logic;
          N_1261_i            : out   std_logic;
          b5_voSc3            : in    std_logic;
          b9_OFWNT9_ab        : in    std_logic;
          b13_wRBtT_ME83hHx   : in    std_logic;
          b5_voSc3_i          : in    std_logic;
          b10_OFWNT9_Y2x      : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic
        );

end b11_OFWNT9s_8tZ_Z3_x;

architecture DEF_ARCH of b11_OFWNT9s_8tZ_Z3_x is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component b19_nczQ_DYg_YFaRM_oUoP_28s_1s_x_0
    port( b8_FZFFLXYE      : in    std_logic_vector(11 downto 0) := (others => 'U');
          b12_PSyi_KyDbLbb : in    std_logic_vector(11 downto 0) := (others => 'U');
          IICE_comm2iice_5 : in    std_logic := 'U';
          IICE_comm2iice_3 : in    std_logic := 'U';
          IICE_comm2iice_0 : in    std_logic := 'U';
          IICE_comm2iice_4 : in    std_logic := 'U';
          b7_yYh03wy5      : in    std_logic := 'U';
          b8_jAA_KlCO      : in    std_logic := 'U';
          ttdo             : out   std_logic
        );
  end component;

  component b13_vFW_xNywD_EdR_174s_12s_4096s_0s_x_0
    port( b11_OFWNT9L_8tZ     : in    std_logic_vector(167 downto 0) := (others => 'U');
          b7_vFW_PlM          : out   std_logic_vector(167 downto 0);
          b12_2_St6KCa_jHv    : in    std_logic_vector(11 downto 0) := (others => 'U');
          b9_v_mzCDYXs        : in    std_logic_vector(11 downto 0) := (others => 'U');
          IICE_comm2iice_0    : in    std_logic := 'U';
          b4_2o_z             : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U'
        );
  end component;

  component b19_nczQ_DYg_YFaRM_oUoP_32s_1s_x_0
    port( IICE_comm2iice_5 : in    std_logic := 'U';
          IICE_comm2iice_3 : in    std_logic := 'U';
          IICE_comm2iice_0 : in    std_logic := 'U';
          IICE_comm2iice_4 : in    std_logic := 'U';
          N_1261_i         : out   std_logic;
          ttdo             : in    std_logic := 'U';
          b7_yYh03wy5      : in    std_logic := 'U';
          b7_yYh03wy4      : in    std_logic := 'U'
        );
  end component;

  component b11_SoWyP0zEFKY_Z2_x_0
    port( mdiclink_reg        : in    std_logic_vector(167 downto 0) := (others => 'U');
          b11_OFWNT9L_8tZ     : out   std_logic_vector(167 downto 0);
          N_145_i             : in    std_logic := 'U';
          b4_2o_z             : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \b12_2_St6KCa_jHv[0]_net_1\, \b12_2_St6KCa_jHv_s[0]\, 
        \b9_v_mzCDYXs[0]\, \b9_v_mzCDYXs_s[0]\, \b3_PfG[156]\, 
        VCC_net_1, \b3_PfG_6[156]\, un1_b7_nYJ_BFM8, GND_net_1, 
        \b3_PfG[157]\, \b3_PfG_6[157]\, \b3_PfG[158]\, 
        \b3_PfG_6[158]\, \b3_PfG[159]\, \b3_PfG_6[159]\, 
        \b3_PfG[160]\, \b3_PfG_6[160]\, \b3_PfG[161]\, 
        \b3_PfG_6[161]\, \b3_PfG[162]\, \b3_PfG_6[162]\, 
        \b3_PfG[163]\, \b3_PfG_6[163]\, \b3_PfG[164]\, 
        \b3_PfG_6[164]\, \b3_PfG[165]\, \b3_PfG_6[165]\, 
        \b3_PfG[166]\, \b3_PfG_6[166]\, \b3_PfG[167]\, 
        \b3_PfG_6[167]\, \b3_PfG[168]\, \b3_PfG_6[168]\, 
        \b3_PfG[141]\, \b3_PfG_6[141]\, \b3_PfG[142]\, 
        \b3_PfG_6[142]\, \b3_PfG[143]\, \b3_PfG_6[143]\, 
        \b3_PfG[144]\, \b3_PfG_6[144]\, \b3_PfG[145]\, 
        \b3_PfG_6[145]\, \b3_PfG[146]\, \b3_PfG_6[146]\, 
        \b3_PfG[147]\, \b3_PfG_6[147]\, \b3_PfG[148]\, 
        \b3_PfG_6[148]\, \b3_PfG[149]\, \b3_PfG_6[149]\, 
        \b3_PfG[150]\, \b3_PfG_6[150]\, \b3_PfG[151]\, 
        \b3_PfG_6[151]\, \b3_PfG[152]\, \b3_PfG_6[152]\, 
        \b3_PfG[153]\, \b3_PfG_6[153]\, \b3_PfG[154]\, 
        \b3_PfG_6[154]\, \b3_PfG[155]\, \b3_PfG_6[155]\, 
        \b3_PfG[126]\, \b3_PfG_6[126]\, \b3_PfG[127]\, 
        \b3_PfG_6[127]\, \b3_PfG[128]\, \b3_PfG_6[128]\, 
        \b3_PfG[129]\, \b3_PfG_6[129]\, \b3_PfG[130]\, 
        \b3_PfG_6[130]\, \b3_PfG[131]\, \b3_PfG_6[131]\, 
        \b3_PfG[132]\, \b3_PfG_6[132]\, \b3_PfG[133]\, 
        \b3_PfG_6[133]\, \b3_PfG[134]\, \b3_PfG_6[134]\, 
        \b3_PfG[135]\, \b3_PfG_6[135]\, \b3_PfG[136]\, 
        \b3_PfG_6[136]\, \b3_PfG[137]\, \b3_PfG_6[137]\, 
        \b3_PfG[138]\, \b3_PfG_6[138]\, \b3_PfG[139]\, 
        \b3_PfG_6[139]\, \b3_PfG[140]\, \b3_PfG_6[140]\, 
        \b3_PfG[111]\, \b3_PfG_6[111]\, \b3_PfG[112]\, 
        \b3_PfG_6[112]\, \b3_PfG[113]\, \b3_PfG_6[113]\, 
        \b3_PfG[114]\, \b3_PfG_6[114]\, \b3_PfG[115]\, 
        \b3_PfG_6[115]\, \b3_PfG[116]\, \b3_PfG_6[116]\, 
        \b3_PfG[117]\, \b3_PfG_6[117]\, \b3_PfG[118]\, 
        \b3_PfG_6[118]\, \b3_PfG[119]\, \b3_PfG_6[119]\, 
        \b3_PfG[120]\, \b3_PfG_6[120]\, \b3_PfG[121]\, 
        \b3_PfG_6[121]\, \b3_PfG[122]\, \b3_PfG_6[122]\, 
        \b3_PfG[123]\, \b3_PfG_6[123]\, \b3_PfG[124]\, 
        \b3_PfG_6[124]\, \b3_PfG[125]\, \b3_PfG_6[125]\, 
        \b3_PfG[96]\, \b3_PfG_6[96]\, \b3_PfG[97]\, 
        \b3_PfG_6[97]\, \b3_PfG[98]\, \b3_PfG_6[98]\, 
        \b3_PfG[99]\, \b3_PfG_6[99]\, \b3_PfG[100]\, 
        \b3_PfG_6[100]\, \b3_PfG[101]\, \b3_PfG_6[101]\, 
        \b3_PfG[102]\, \b3_PfG_6[102]\, \b3_PfG[103]\, 
        \b3_PfG_6[103]\, \b3_PfG[104]\, \b3_PfG_6[104]\, 
        \b3_PfG[105]\, \b3_PfG_6[105]\, \b3_PfG[106]\, 
        \b3_PfG_6[106]\, \b3_PfG[107]\, \b3_PfG_6[107]\, 
        \b3_PfG[108]\, \b3_PfG_6[108]\, \b3_PfG[109]\, 
        \b3_PfG_6[109]\, \b3_PfG[110]\, \b3_PfG_6[110]\, 
        \b3_PfG[81]\, \b3_PfG_6[81]\, \b3_PfG[82]\, 
        \b3_PfG_6[82]\, \b3_PfG[83]\, \b3_PfG_6[83]\, 
        \b3_PfG[84]\, \b3_PfG_6[84]\, \b3_PfG[85]\, 
        \b3_PfG_6[85]\, \b3_PfG[86]\, \b3_PfG_6[86]\, 
        \b3_PfG[87]\, \b3_PfG_6[87]\, \b3_PfG[88]\, 
        \b3_PfG_6[88]\, \b3_PfG[89]\, \b3_PfG_6[89]\, 
        \b3_PfG[90]\, \b3_PfG_6[90]\, \b3_PfG[91]\, 
        \b3_PfG_6[91]\, \b3_PfG[92]\, \b3_PfG_6[92]\, 
        \b3_PfG[93]\, \b3_PfG_6[93]\, \b3_PfG[94]\, 
        \b3_PfG_6[94]\, \b3_PfG[95]\, \b3_PfG_6[95]\, 
        \b3_PfG[66]\, \b3_PfG_6[66]\, \b3_PfG[67]\, 
        \b3_PfG_6[67]\, \b3_PfG[68]\, \b3_PfG_6[68]\, 
        \b3_PfG[69]\, \b3_PfG_6[69]\, \b3_PfG[70]\, 
        \b3_PfG_6[70]\, \b3_PfG[71]\, \b3_PfG_6[71]\, 
        \b3_PfG[72]\, \b3_PfG_6[72]\, \b3_PfG[73]\, 
        \b3_PfG_6[73]\, \b3_PfG[74]\, \b3_PfG_6[74]\, 
        \b3_PfG[75]\, \b3_PfG_6[75]\, \b3_PfG[76]\, 
        \b3_PfG_6[76]\, \b3_PfG[77]\, \b3_PfG_6[77]\, 
        \b3_PfG[78]\, \b3_PfG_6[78]\, \b3_PfG[79]\, 
        \b3_PfG_6[79]\, \b3_PfG[80]\, \b3_PfG_6[80]\, 
        \b3_PfG[51]\, \b3_PfG_6[51]\, \b3_PfG[52]\, 
        \b3_PfG_6[52]\, \b3_PfG[53]\, \b3_PfG_6[53]\, 
        \b3_PfG[54]\, \b3_PfG_6[54]\, \b3_PfG[55]\, 
        \b3_PfG_6[55]\, \b3_PfG[56]\, \b3_PfG_6[56]\, 
        \b3_PfG[57]\, \b3_PfG_6[57]\, \b3_PfG[58]\, 
        \b3_PfG_6[58]\, \b3_PfG[59]\, \b3_PfG_6[59]\, 
        \b3_PfG[60]\, \b3_PfG_6[60]\, \b3_PfG[61]\, 
        \b3_PfG_6[61]\, \b3_PfG[62]\, \b3_PfG_6[62]\, 
        \b3_PfG[63]\, \b3_PfG_6[63]\, \b3_PfG[64]\, 
        \b3_PfG_6[64]\, \b3_PfG[65]\, \b3_PfG_6[65]\, 
        \b3_PfG[36]\, \b3_PfG_6[36]\, \b3_PfG[37]\, 
        \b3_PfG_6[37]\, \b3_PfG[38]\, \b3_PfG_6[38]\, 
        \b3_PfG[39]\, \b3_PfG_6[39]\, \b3_PfG[40]\, 
        \b3_PfG_6[40]\, \b3_PfG[41]\, \b3_PfG_6[41]\, 
        \b3_PfG[42]\, \b3_PfG_6[42]\, \b3_PfG[43]\, 
        \b3_PfG_6[43]\, \b3_PfG[44]\, \b3_PfG_6[44]\, 
        \b3_PfG[45]\, \b3_PfG_6[45]\, \b3_PfG[46]\, 
        \b3_PfG_6[46]\, \b3_PfG[47]\, \b3_PfG_6[47]\, 
        \b3_PfG[48]\, \b3_PfG_6[48]\, \b3_PfG[49]\, 
        \b3_PfG_6[49]\, \b3_PfG[50]\, \b3_PfG_6[50]\, 
        \b3_PfG[21]\, \b3_PfG_6[21]\, \b3_PfG[22]\, 
        \b3_PfG_6[22]\, \b3_PfG[23]\, \b3_PfG_6[23]\, 
        \b3_PfG[24]\, \b3_PfG_6[24]\, \b3_PfG[25]\, 
        \b3_PfG_6[25]\, \b3_PfG[26]\, \b3_PfG_6[26]\, 
        \b3_PfG[27]\, \b3_PfG_6[27]\, \b3_PfG[28]\, 
        \b3_PfG_6[28]\, \b3_PfG[29]\, \b3_PfG_6[29]\, 
        \b3_PfG[30]\, \b3_PfG_6[30]\, \b3_PfG[31]\, 
        \b3_PfG_6[31]\, \b3_PfG[32]\, \b3_PfG_6[32]\, 
        \b3_PfG[33]\, \b3_PfG_6[33]\, \b3_PfG[34]\, 
        \b3_PfG_6[34]\, \b3_PfG[35]\, \b3_PfG_6[35]\, \b3_PfG[6]\, 
        \b3_PfG_6[6]\, \b3_PfG[7]\, \b3_PfG_6[7]\, \b3_PfG[8]\, 
        \b3_PfG_6[8]\, \b3_PfG[9]\, \b3_PfG_6[9]\, \b3_PfG[10]\, 
        \b3_PfG_6[10]\, \b3_PfG[11]\, \b3_PfG_6[11]\, 
        \b3_PfG[12]\, \b3_PfG_6[12]\, \b3_PfG[13]\, 
        \b3_PfG_6[13]\, \b3_PfG[14]\, \b3_PfG_6[14]\, 
        \b3_PfG[15]\, \b3_PfG_6[15]\, \b3_PfG[16]\, 
        \b3_PfG_6[16]\, \b3_PfG[17]\, \b3_PfG_6[17]\, 
        \b3_PfG[18]\, \b3_PfG_6[18]\, \b3_PfG[19]\, 
        \b3_PfG_6[19]\, \b3_PfG[20]\, \b3_PfG_6[20]\, 
        \b12_PSyi_KyDbLbb[3]_net_1\, \b12_2_St6KCa_jHv[3]_net_1\, 
        \b12_PSyi_KyDbLbb_0_sqmuxa\, \b12_PSyi_KyDbLbb[4]_net_1\, 
        \b12_2_St6KCa_jHv[4]_net_1\, \b12_PSyi_KyDbLbb[5]_net_1\, 
        \b12_2_St6KCa_jHv[5]_net_1\, \b12_PSyi_KyDbLbb[6]_net_1\, 
        \b12_2_St6KCa_jHv[6]_net_1\, \b12_PSyi_KyDbLbb[7]_net_1\, 
        \b12_2_St6KCa_jHv[7]_net_1\, \b12_PSyi_KyDbLbb[8]_net_1\, 
        \b12_2_St6KCa_jHv[8]_net_1\, \b12_PSyi_KyDbLbb[9]_net_1\, 
        \b12_2_St6KCa_jHv[9]_net_1\, \b12_PSyi_KyDbLbb[10]_net_1\, 
        \b12_2_St6KCa_jHv[10]_net_1\, 
        \b12_PSyi_KyDbLbb[11]_net_1\, 
        \b12_2_St6KCa_jHv[11]_net_1\, \b3_PfG_6[0]\, \b3_PfG[1]\, 
        \b3_PfG_6[1]\, \b3_PfG[2]\, \b3_PfG_6[2]\, \b3_PfG[3]\, 
        \b3_PfG_6[3]\, \b3_PfG[4]\, \b3_PfG_6[4]\, \b3_PfG[5]\, 
        \b3_PfG_6[5]\, \b8_FZFFLXYE[0]_net_1\, b4_2o_z, 
        \b8_FZFFLXYE[1]_net_1\, \b12_2_St6KCa_jHv[1]_net_1\, 
        \b8_FZFFLXYE[2]_net_1\, \b12_2_St6KCa_jHv[2]_net_1\, 
        \b8_FZFFLXYE[3]_net_1\, \b8_FZFFLXYE[4]_net_1\, 
        \b8_FZFFLXYE[5]_net_1\, \b8_FZFFLXYE[6]_net_1\, 
        \b8_FZFFLXYE[7]_net_1\, \b8_FZFFLXYE[8]_net_1\, 
        \b8_FZFFLXYE[9]_net_1\, \b8_FZFFLXYE[10]_net_1\, 
        \b8_FZFFLXYE[11]_net_1\, \b12_PSyi_KyDbLbb[0]_net_1\, 
        \b12_PSyi_KyDbLbb[1]_net_1\, \b12_PSyi_KyDbLbb[2]_net_1\, 
        \b7_nYJ_BFM[171]\, \b7_nYJ_BFM[170]\, \N_15_i\, 
        \b7_nYJ_BFM[172]\, \b7_nYJ_BFM[173]\, \b7_nYJ_BFM[174]\, 
        \b7_nYJ_BFM[156]\, \b7_nYJ_BFM[155]\, \b7_nYJ_BFM[157]\, 
        \b7_nYJ_BFM[158]\, \b7_nYJ_BFM[159]\, \b7_nYJ_BFM[160]\, 
        \b7_nYJ_BFM[161]\, \b7_nYJ_BFM[162]\, \b7_nYJ_BFM[163]\, 
        \b7_nYJ_BFM[164]\, \b7_nYJ_BFM[165]\, \b7_nYJ_BFM[166]\, 
        \b7_nYJ_BFM[167]\, \b7_nYJ_BFM[168]\, \b7_nYJ_BFM[169]\, 
        \b7_nYJ_BFM[141]\, \b7_nYJ_BFM[140]\, \b7_nYJ_BFM[142]\, 
        \b7_nYJ_BFM[143]\, \b7_nYJ_BFM[144]\, \b7_nYJ_BFM[145]\, 
        \b7_nYJ_BFM[146]\, \b7_nYJ_BFM[147]\, \b7_nYJ_BFM[148]\, 
        \b7_nYJ_BFM[149]\, \b7_nYJ_BFM[150]\, \b7_nYJ_BFM[151]\, 
        \b7_nYJ_BFM[152]\, \b7_nYJ_BFM[153]\, \b7_nYJ_BFM[154]\, 
        \b7_nYJ_BFM[126]\, \b7_nYJ_BFM[125]\, \b7_nYJ_BFM[127]\, 
        \b7_nYJ_BFM[128]\, \b7_nYJ_BFM[129]\, \b7_nYJ_BFM[130]\, 
        \b7_nYJ_BFM[131]\, \b7_nYJ_BFM[132]\, \b7_nYJ_BFM[133]\, 
        \b7_nYJ_BFM[134]\, \b7_nYJ_BFM[135]\, \b7_nYJ_BFM[136]\, 
        \b7_nYJ_BFM[137]\, \b7_nYJ_BFM[138]\, \b7_nYJ_BFM[139]\, 
        \b7_nYJ_BFM[111]\, \b7_nYJ_BFM[110]\, \b7_nYJ_BFM[112]\, 
        \b7_nYJ_BFM[113]\, \b7_nYJ_BFM[114]\, \b7_nYJ_BFM[115]\, 
        \b7_nYJ_BFM[116]\, \b7_nYJ_BFM[117]\, \b7_nYJ_BFM[118]\, 
        \b7_nYJ_BFM[119]\, \b7_nYJ_BFM[120]\, \b7_nYJ_BFM[121]\, 
        \b7_nYJ_BFM[122]\, \b7_nYJ_BFM[123]\, \b7_nYJ_BFM[124]\, 
        \b7_nYJ_BFM[96]\, \b7_nYJ_BFM[95]\, \b7_nYJ_BFM[97]\, 
        \b7_nYJ_BFM[98]\, \b7_nYJ_BFM[99]\, \b7_nYJ_BFM[100]\, 
        \b7_nYJ_BFM[101]\, \b7_nYJ_BFM[102]\, \b7_nYJ_BFM[103]\, 
        \b7_nYJ_BFM[104]\, \b7_nYJ_BFM[105]\, \b7_nYJ_BFM[106]\, 
        \b7_nYJ_BFM[107]\, \b7_nYJ_BFM[108]\, \b7_nYJ_BFM[109]\, 
        \b7_nYJ_BFM[81]\, \b7_nYJ_BFM[80]\, \b7_nYJ_BFM[82]\, 
        \b7_nYJ_BFM[83]\, \b7_nYJ_BFM[84]\, \b7_nYJ_BFM[85]\, 
        \b7_nYJ_BFM[86]\, \b7_nYJ_BFM[87]\, \b7_nYJ_BFM[88]\, 
        \b7_nYJ_BFM[89]\, \b7_nYJ_BFM[90]\, \b7_nYJ_BFM[91]\, 
        \b7_nYJ_BFM[92]\, \b7_nYJ_BFM[93]\, \b7_nYJ_BFM[94]\, 
        \b7_nYJ_BFM[66]\, \b7_nYJ_BFM[65]\, \b7_nYJ_BFM[67]\, 
        \b7_nYJ_BFM[68]\, \b7_nYJ_BFM[69]\, \b7_nYJ_BFM[70]\, 
        \b7_nYJ_BFM[71]\, \b7_nYJ_BFM[72]\, \b7_nYJ_BFM[73]\, 
        \b7_nYJ_BFM[74]\, \b7_nYJ_BFM[75]\, \b7_nYJ_BFM[76]\, 
        \b7_nYJ_BFM[77]\, \b7_nYJ_BFM[78]\, \b7_nYJ_BFM[79]\, 
        \b7_nYJ_BFM[51]\, \b7_nYJ_BFM[50]\, \b7_nYJ_BFM[52]\, 
        \b7_nYJ_BFM[53]\, \b7_nYJ_BFM[54]\, \b7_nYJ_BFM[55]\, 
        \b7_nYJ_BFM[56]\, \b7_nYJ_BFM[57]\, \b7_nYJ_BFM[58]\, 
        \b7_nYJ_BFM[59]\, \b7_nYJ_BFM[60]\, \b7_nYJ_BFM[61]\, 
        \b7_nYJ_BFM[62]\, \b7_nYJ_BFM[63]\, \b7_nYJ_BFM[64]\, 
        \b7_nYJ_BFM[36]\, \b7_nYJ_BFM[35]\, \b7_nYJ_BFM[37]\, 
        \b7_nYJ_BFM[38]\, \b7_nYJ_BFM[39]\, \b7_nYJ_BFM[40]\, 
        \b7_nYJ_BFM[41]\, \b7_nYJ_BFM[42]\, \b7_nYJ_BFM[43]\, 
        \b7_nYJ_BFM[44]\, \b7_nYJ_BFM[45]\, \b7_nYJ_BFM[46]\, 
        \b7_nYJ_BFM[47]\, \b7_nYJ_BFM[48]\, \b7_nYJ_BFM[49]\, 
        \b7_nYJ_BFM[21]\, \b7_nYJ_BFM[20]\, \b7_nYJ_BFM[22]\, 
        \b7_nYJ_BFM[23]\, \b7_nYJ_BFM[24]\, \b7_nYJ_BFM[25]\, 
        \b7_nYJ_BFM[26]\, \b7_nYJ_BFM[27]\, \b7_nYJ_BFM[28]\, 
        \b7_nYJ_BFM[29]\, \b7_nYJ_BFM[30]\, \b7_nYJ_BFM[31]\, 
        \b7_nYJ_BFM[32]\, \b7_nYJ_BFM[33]\, \b7_nYJ_BFM[34]\, 
        \b7_nYJ_BFM[6]\, \b7_nYJ_BFM[5]\, \b7_nYJ_BFM[7]\, 
        \b7_nYJ_BFM[8]\, \b7_nYJ_BFM[9]\, \b7_nYJ_BFM[10]\, 
        \b7_nYJ_BFM[11]\, \b7_nYJ_BFM[12]\, \b7_nYJ_BFM[13]\, 
        \b7_nYJ_BFM[14]\, \b7_nYJ_BFM[15]\, \b7_nYJ_BFM[16]\, 
        \b7_nYJ_BFM[17]\, \b7_nYJ_BFM[18]\, \b7_nYJ_BFM[19]\, 
        \b8_jAA_KlCO\, \b8_jAA_KlCO_0_sqmuxa\, \b7_nYJ_BFM[0]\, 
        \b7_nYJ_BFM[1]\, \b7_nYJ_BFM[2]\, \b7_nYJ_BFM[3]\, 
        \b7_nYJ_BFM[4]\, \b9_PSyil9s_2\, b11_nFG0rDY_9e2, 
        b11_nFG0rDY_9e2_2, b9_v_mzCDYXs13, \b9_v_mzCDYXs[1]\, 
        \b9_v_mzCDYXs_s[1]\, \b9_v_mzCDYXs[2]\, 
        \b9_v_mzCDYXs_s[2]\, \b9_v_mzCDYXs[3]\, 
        \b9_v_mzCDYXs_s[3]\, \b9_v_mzCDYXs[4]\, 
        \b9_v_mzCDYXs_s[4]\, \b9_v_mzCDYXs[5]\, 
        \b9_v_mzCDYXs_s[5]\, \b9_v_mzCDYXs[6]\, 
        \b9_v_mzCDYXs_s[6]\, \b9_v_mzCDYXs[7]\, 
        \b9_v_mzCDYXs_s[7]\, \b9_v_mzCDYXs[8]\, 
        \b9_v_mzCDYXs_s[8]\, \b9_v_mzCDYXs[9]\, 
        \b9_v_mzCDYXs_s[9]\, \b9_v_mzCDYXs[10]\, 
        \b9_v_mzCDYXs_s[10]\, \b9_v_mzCDYXs[11]\, 
        \b9_v_mzCDYXs_s[11]\, \b12_2_St6KCa_jHv_s[1]\, 
        \b12_2_St6KCa_jHv_s[2]\, \b12_2_St6KCa_jHv_s[3]\, 
        \b12_2_St6KCa_jHv_s[4]\, \b12_2_St6KCa_jHv_s[5]\, 
        \b12_2_St6KCa_jHv_s[6]\, \b12_2_St6KCa_jHv_s[7]\, 
        \b12_2_St6KCa_jHv_s[8]\, \b12_2_St6KCa_jHv_s[9]\, 
        \b12_2_St6KCa_jHv_s[10]\, \b12_2_St6KCa_jHv_s[11]_net_1\, 
        b12_2_St6KCa_jHv_s_900_FCO, 
        \b12_2_St6KCa_jHv_cry[1]_net_1\, 
        \b12_2_St6KCa_jHv_cry[2]_net_1\, 
        \b12_2_St6KCa_jHv_cry[3]_net_1\, 
        \b12_2_St6KCa_jHv_cry[4]_net_1\, 
        \b12_2_St6KCa_jHv_cry[5]_net_1\, 
        \b12_2_St6KCa_jHv_cry[6]_net_1\, 
        \b12_2_St6KCa_jHv_cry[7]_net_1\, 
        \b12_2_St6KCa_jHv_cry[8]_net_1\, 
        \b12_2_St6KCa_jHv_cry[9]_net_1\, 
        \b12_2_St6KCa_jHv_cry[10]_net_1\, b9_v_mzCDYXs_s_901_FCO, 
        \b9_v_mzCDYXs_cry[1]\, \b9_v_mzCDYXs_cry[2]\, 
        \b9_v_mzCDYXs_cry[3]\, \b9_v_mzCDYXs_cry[4]\, 
        \b9_v_mzCDYXs_cry[5]\, \b9_v_mzCDYXs_cry[6]\, 
        \b9_v_mzCDYXs_cry[7]\, \b9_v_mzCDYXs_cry[8]\, 
        \b9_v_mzCDYXs_cry[9]\, \b9_v_mzCDYXs_cry[10]\, 
        \b7_vFW_PlM[167]\, \b7_vFW_PlM[166]\, \b7_vFW_PlM[165]\, 
        \b7_vFW_PlM[164]\, \b7_vFW_PlM[163]\, \b7_vFW_PlM[162]\, 
        \b7_vFW_PlM[161]\, \b7_vFW_PlM[160]\, \b7_vFW_PlM[159]\, 
        \b7_vFW_PlM[158]\, \b7_vFW_PlM[157]\, \b7_vFW_PlM[156]\, 
        \b7_vFW_PlM[155]\, \b7_vFW_PlM[154]\, \b7_vFW_PlM[153]\, 
        \b7_vFW_PlM[152]\, \b7_vFW_PlM[151]\, \b7_vFW_PlM[150]\, 
        \b7_vFW_PlM[149]\, \b7_vFW_PlM[148]\, \b7_vFW_PlM[147]\, 
        \b7_vFW_PlM[146]\, \b7_vFW_PlM[145]\, \b7_vFW_PlM[144]\, 
        \b7_vFW_PlM[143]\, \b7_vFW_PlM[142]\, \b7_vFW_PlM[141]\, 
        \b7_vFW_PlM[140]\, \b7_vFW_PlM[139]\, \b7_vFW_PlM[138]\, 
        \b7_vFW_PlM[137]\, \b7_vFW_PlM[136]\, \b7_vFW_PlM[135]\, 
        \b7_vFW_PlM[134]\, \b7_vFW_PlM[133]\, \b7_vFW_PlM[132]\, 
        \b7_vFW_PlM[131]\, \b7_vFW_PlM[130]\, \b7_vFW_PlM[129]\, 
        \b7_vFW_PlM[128]\, \b7_vFW_PlM[127]\, \b7_vFW_PlM[126]\, 
        \b7_vFW_PlM[125]\, \b7_vFW_PlM[124]\, \b7_vFW_PlM[123]\, 
        \b7_vFW_PlM[122]\, \b7_vFW_PlM[121]\, \b7_vFW_PlM[120]\, 
        \b7_vFW_PlM[119]\, \b7_vFW_PlM[118]\, \b7_vFW_PlM[117]\, 
        \b7_vFW_PlM[116]\, \b7_vFW_PlM[115]\, \b7_vFW_PlM[114]\, 
        \b7_vFW_PlM[113]\, \b7_vFW_PlM[112]\, \b7_vFW_PlM[111]\, 
        \b7_vFW_PlM[110]\, \b7_vFW_PlM[109]\, \b7_vFW_PlM[108]\, 
        \b7_vFW_PlM[107]\, \b7_vFW_PlM[106]\, \b7_vFW_PlM[105]\, 
        \b7_vFW_PlM[104]\, \b7_vFW_PlM[103]\, \b7_vFW_PlM[102]\, 
        \b7_vFW_PlM[101]\, \b7_vFW_PlM[100]\, \b7_vFW_PlM[99]\, 
        \b7_vFW_PlM[98]\, \b7_vFW_PlM[97]\, \b7_vFW_PlM[96]\, 
        \b7_vFW_PlM[95]\, \b7_vFW_PlM[94]\, \b7_vFW_PlM[93]\, 
        \b7_vFW_PlM[92]\, \b7_vFW_PlM[91]\, \b7_vFW_PlM[90]\, 
        \b7_vFW_PlM[89]\, \b7_vFW_PlM[88]\, \b7_vFW_PlM[87]\, 
        \b7_vFW_PlM[86]\, \b7_vFW_PlM[85]\, \b7_vFW_PlM[84]\, 
        \b7_vFW_PlM[83]\, \b7_vFW_PlM[82]\, \b7_vFW_PlM[81]\, 
        \b7_vFW_PlM[80]\, \b7_vFW_PlM[79]\, \b7_vFW_PlM[78]\, 
        \b7_vFW_PlM[77]\, \b7_vFW_PlM[76]\, \b7_vFW_PlM[75]\, 
        \b7_vFW_PlM[74]\, \b7_vFW_PlM[73]\, \b7_vFW_PlM[72]\, 
        \b7_vFW_PlM[71]\, \b7_vFW_PlM[70]\, \b7_vFW_PlM[69]\, 
        \b7_vFW_PlM[68]\, \b7_vFW_PlM[67]\, \b7_vFW_PlM[66]\, 
        \b7_vFW_PlM[65]\, \b7_vFW_PlM[64]\, \b7_vFW_PlM[63]\, 
        \b7_vFW_PlM[62]\, \b7_vFW_PlM[61]\, \b7_vFW_PlM[60]\, 
        \b7_vFW_PlM[59]\, \b7_vFW_PlM[58]\, \b7_vFW_PlM[57]\, 
        \b7_vFW_PlM[56]\, \b7_vFW_PlM[55]\, \b7_vFW_PlM[54]\, 
        \b7_vFW_PlM[53]\, \b7_vFW_PlM[52]\, \b7_vFW_PlM[51]\, 
        \b7_vFW_PlM[50]\, \b7_vFW_PlM[49]\, \b7_vFW_PlM[48]\, 
        \b7_vFW_PlM[47]\, \b7_vFW_PlM[46]\, \b7_vFW_PlM[45]\, 
        \b7_vFW_PlM[44]\, \b7_vFW_PlM[43]\, \b7_vFW_PlM[42]\, 
        \b7_vFW_PlM[41]\, \b7_vFW_PlM[40]\, \b7_vFW_PlM[39]\, 
        \b7_vFW_PlM[38]\, \b7_vFW_PlM[37]\, \b7_vFW_PlM[36]\, 
        \b7_vFW_PlM[35]\, \b7_vFW_PlM[34]\, \b7_vFW_PlM[33]\, 
        \b7_vFW_PlM[32]\, \b7_vFW_PlM[31]\, \b7_vFW_PlM[30]\, 
        \b7_vFW_PlM[29]\, \b7_vFW_PlM[28]\, \b7_vFW_PlM[27]\, 
        \b7_vFW_PlM[26]\, \b7_vFW_PlM[25]\, \b7_vFW_PlM[24]\, 
        \b7_vFW_PlM[23]\, \b7_vFW_PlM[22]\, \b7_vFW_PlM[21]\, 
        \b7_vFW_PlM[20]\, \b7_vFW_PlM[19]\, \b7_vFW_PlM[18]\, 
        \b7_vFW_PlM[17]\, \b7_vFW_PlM[16]\, \b7_vFW_PlM[15]\, 
        \b7_vFW_PlM[14]\, \b7_vFW_PlM[13]\, \b7_vFW_PlM[12]\, 
        \b7_vFW_PlM[11]\, \b7_vFW_PlM[10]\, \b7_vFW_PlM[9]\, 
        \b7_vFW_PlM[8]\, \b7_vFW_PlM[7]\, \b7_vFW_PlM[6]\, 
        \b7_vFW_PlM[5]\, \b7_vFW_PlM[4]\, \b7_vFW_PlM[3]\, 
        \b7_vFW_PlM[2]\, \b7_vFW_PlM[1]\, \b7_vFW_PlM[0]\, 
        \b8_jAA_KlCO_0_sqmuxa_8\, \b8_jAA_KlCO_0_sqmuxa_7\, 
        \b8_jAA_KlCO_0_sqmuxa_1\, \b7_yYh03wy4_0_a2_0_2\, 
        b7_yYh03wy5, b7_yYh03wy4, ttdo, \b11_OFWNT9L_8tZ[0]\, 
        \b11_OFWNT9L_8tZ[1]\, \b11_OFWNT9L_8tZ[2]\, 
        \b11_OFWNT9L_8tZ[3]\, \b11_OFWNT9L_8tZ[4]\, 
        \b11_OFWNT9L_8tZ[5]\, \b11_OFWNT9L_8tZ[6]\, 
        \b11_OFWNT9L_8tZ[7]\, \b11_OFWNT9L_8tZ[8]\, 
        \b11_OFWNT9L_8tZ[9]\, \b11_OFWNT9L_8tZ[10]\, 
        \b11_OFWNT9L_8tZ[11]\, \b11_OFWNT9L_8tZ[12]\, 
        \b11_OFWNT9L_8tZ[13]\, \b11_OFWNT9L_8tZ[14]\, 
        \b11_OFWNT9L_8tZ[15]\, \b11_OFWNT9L_8tZ[16]\, 
        \b11_OFWNT9L_8tZ[17]\, \b11_OFWNT9L_8tZ[18]\, 
        \b11_OFWNT9L_8tZ[19]\, \b11_OFWNT9L_8tZ[20]\, 
        \b11_OFWNT9L_8tZ[21]\, \b11_OFWNT9L_8tZ[22]\, 
        \b11_OFWNT9L_8tZ[23]\, \b11_OFWNT9L_8tZ[24]\, 
        \b11_OFWNT9L_8tZ[25]\, \b11_OFWNT9L_8tZ[26]\, 
        \b11_OFWNT9L_8tZ[27]\, \b11_OFWNT9L_8tZ[28]\, 
        \b11_OFWNT9L_8tZ[29]\, \b11_OFWNT9L_8tZ[30]\, 
        \b11_OFWNT9L_8tZ[31]\, \b11_OFWNT9L_8tZ[32]\, 
        \b11_OFWNT9L_8tZ[33]\, \b11_OFWNT9L_8tZ[34]\, 
        \b11_OFWNT9L_8tZ[35]\, \b11_OFWNT9L_8tZ[36]\, 
        \b11_OFWNT9L_8tZ[37]\, \b11_OFWNT9L_8tZ[38]\, 
        \b11_OFWNT9L_8tZ[39]\, \b11_OFWNT9L_8tZ[40]\, 
        \b11_OFWNT9L_8tZ[41]\, \b11_OFWNT9L_8tZ[42]\, 
        \b11_OFWNT9L_8tZ[43]\, \b11_OFWNT9L_8tZ[44]\, 
        \b11_OFWNT9L_8tZ[45]\, \b11_OFWNT9L_8tZ[46]\, 
        \b11_OFWNT9L_8tZ[47]\, \b11_OFWNT9L_8tZ[48]\, 
        \b11_OFWNT9L_8tZ[49]\, \b11_OFWNT9L_8tZ[50]\, 
        \b11_OFWNT9L_8tZ[51]\, \b11_OFWNT9L_8tZ[52]\, 
        \b11_OFWNT9L_8tZ[53]\, \b11_OFWNT9L_8tZ[54]\, 
        \b11_OFWNT9L_8tZ[55]\, \b11_OFWNT9L_8tZ[56]\, 
        \b11_OFWNT9L_8tZ[57]\, \b11_OFWNT9L_8tZ[58]\, 
        \b11_OFWNT9L_8tZ[59]\, \b11_OFWNT9L_8tZ[60]\, 
        \b11_OFWNT9L_8tZ[61]\, \b11_OFWNT9L_8tZ[62]\, 
        \b11_OFWNT9L_8tZ[63]\, \b11_OFWNT9L_8tZ[64]\, 
        \b11_OFWNT9L_8tZ[65]\, \b11_OFWNT9L_8tZ[66]\, 
        \b11_OFWNT9L_8tZ[67]\, \b11_OFWNT9L_8tZ[68]\, 
        \b11_OFWNT9L_8tZ[69]\, \b11_OFWNT9L_8tZ[70]\, 
        \b11_OFWNT9L_8tZ[71]\, \b11_OFWNT9L_8tZ[72]\, 
        \b11_OFWNT9L_8tZ[73]\, \b11_OFWNT9L_8tZ[74]\, 
        \b11_OFWNT9L_8tZ[75]\, \b11_OFWNT9L_8tZ[76]\, 
        \b11_OFWNT9L_8tZ[77]\, \b11_OFWNT9L_8tZ[78]\, 
        \b11_OFWNT9L_8tZ[79]\, \b11_OFWNT9L_8tZ[80]\, 
        \b11_OFWNT9L_8tZ[81]\, \b11_OFWNT9L_8tZ[82]\, 
        \b11_OFWNT9L_8tZ[83]\, \b11_OFWNT9L_8tZ[84]\, 
        \b11_OFWNT9L_8tZ[85]\, \b11_OFWNT9L_8tZ[86]\, 
        \b11_OFWNT9L_8tZ[87]\, \b11_OFWNT9L_8tZ[88]\, 
        \b11_OFWNT9L_8tZ[89]\, \b11_OFWNT9L_8tZ[90]\, 
        \b11_OFWNT9L_8tZ[91]\, \b11_OFWNT9L_8tZ[92]\, 
        \b11_OFWNT9L_8tZ[93]\, \b11_OFWNT9L_8tZ[94]\, 
        \b11_OFWNT9L_8tZ[95]\, \b11_OFWNT9L_8tZ[96]\, 
        \b11_OFWNT9L_8tZ[97]\, \b11_OFWNT9L_8tZ[98]\, 
        \b11_OFWNT9L_8tZ[99]\, \b11_OFWNT9L_8tZ[100]\, 
        \b11_OFWNT9L_8tZ[101]\, \b11_OFWNT9L_8tZ[102]\, 
        \b11_OFWNT9L_8tZ[103]\, \b11_OFWNT9L_8tZ[104]\, 
        \b11_OFWNT9L_8tZ[105]\, \b11_OFWNT9L_8tZ[106]\, 
        \b11_OFWNT9L_8tZ[107]\, \b11_OFWNT9L_8tZ[108]\, 
        \b11_OFWNT9L_8tZ[109]\, \b11_OFWNT9L_8tZ[110]\, 
        \b11_OFWNT9L_8tZ[111]\, \b11_OFWNT9L_8tZ[112]\, 
        \b11_OFWNT9L_8tZ[113]\, \b11_OFWNT9L_8tZ[114]\, 
        \b11_OFWNT9L_8tZ[115]\, \b11_OFWNT9L_8tZ[116]\, 
        \b11_OFWNT9L_8tZ[117]\, \b11_OFWNT9L_8tZ[118]\, 
        \b11_OFWNT9L_8tZ[119]\, \b11_OFWNT9L_8tZ[120]\, 
        \b11_OFWNT9L_8tZ[121]\, \b11_OFWNT9L_8tZ[122]\, 
        \b11_OFWNT9L_8tZ[123]\, \b11_OFWNT9L_8tZ[124]\, 
        \b11_OFWNT9L_8tZ[125]\, \b11_OFWNT9L_8tZ[126]\, 
        \b11_OFWNT9L_8tZ[127]\, \b11_OFWNT9L_8tZ[128]\, 
        \b11_OFWNT9L_8tZ[129]\, \b11_OFWNT9L_8tZ[130]\, 
        \b11_OFWNT9L_8tZ[131]\, \b11_OFWNT9L_8tZ[132]\, 
        \b11_OFWNT9L_8tZ[133]\, \b11_OFWNT9L_8tZ[134]\, 
        \b11_OFWNT9L_8tZ[135]\, \b11_OFWNT9L_8tZ[136]\, 
        \b11_OFWNT9L_8tZ[137]\, \b11_OFWNT9L_8tZ[138]\, 
        \b11_OFWNT9L_8tZ[139]\, \b11_OFWNT9L_8tZ[140]\, 
        \b11_OFWNT9L_8tZ[141]\, \b11_OFWNT9L_8tZ[142]\, 
        \b11_OFWNT9L_8tZ[143]\, \b11_OFWNT9L_8tZ[144]\, 
        \b11_OFWNT9L_8tZ[145]\, \b11_OFWNT9L_8tZ[146]\, 
        \b11_OFWNT9L_8tZ[147]\, \b11_OFWNT9L_8tZ[148]\, 
        \b11_OFWNT9L_8tZ[149]\, \b11_OFWNT9L_8tZ[150]\, 
        \b11_OFWNT9L_8tZ[151]\, \b11_OFWNT9L_8tZ[152]\, 
        \b11_OFWNT9L_8tZ[153]\, \b11_OFWNT9L_8tZ[154]\, 
        \b11_OFWNT9L_8tZ[155]\, \b11_OFWNT9L_8tZ[156]\, 
        \b11_OFWNT9L_8tZ[157]\, \b11_OFWNT9L_8tZ[158]\, 
        \b11_OFWNT9L_8tZ[159]\, \b11_OFWNT9L_8tZ[160]\, 
        \b11_OFWNT9L_8tZ[161]\, \b11_OFWNT9L_8tZ[162]\, 
        \b11_OFWNT9L_8tZ[163]\, \b11_OFWNT9L_8tZ[164]\, 
        \b11_OFWNT9L_8tZ[165]\, \b11_OFWNT9L_8tZ[166]\, 
        \b11_OFWNT9L_8tZ[167]\ : std_logic;

    for all : b19_nczQ_DYg_YFaRM_oUoP_28s_1s_x_0
	Use entity work.b19_nczQ_DYg_YFaRM_oUoP_28s_1s_x_0(DEF_ARCH);
    for all : b13_vFW_xNywD_EdR_174s_12s_4096s_0s_x_0
	Use entity work.
        b13_vFW_xNywD_EdR_174s_12s_4096s_0s_x_0(DEF_ARCH);
    for all : b19_nczQ_DYg_YFaRM_oUoP_32s_1s_x_0
	Use entity work.b19_nczQ_DYg_YFaRM_oUoP_32s_1s_x_0(DEF_ARCH);
    for all : b11_SoWyP0zEFKY_Z2_x_0
	Use entity work.b11_SoWyP0zEFKY_Z2_x_0(DEF_ARCH);
begin 

    b11_OFWNT9L_8tZ(167) <= \b11_OFWNT9L_8tZ[167]\;
    b11_OFWNT9L_8tZ(166) <= \b11_OFWNT9L_8tZ[166]\;
    b11_OFWNT9L_8tZ(165) <= \b11_OFWNT9L_8tZ[165]\;
    b11_OFWNT9L_8tZ(164) <= \b11_OFWNT9L_8tZ[164]\;
    b11_OFWNT9L_8tZ(163) <= \b11_OFWNT9L_8tZ[163]\;
    b11_OFWNT9L_8tZ(162) <= \b11_OFWNT9L_8tZ[162]\;
    b11_OFWNT9L_8tZ(161) <= \b11_OFWNT9L_8tZ[161]\;
    b11_OFWNT9L_8tZ(160) <= \b11_OFWNT9L_8tZ[160]\;
    b11_OFWNT9L_8tZ(159) <= \b11_OFWNT9L_8tZ[159]\;
    b11_OFWNT9L_8tZ(158) <= \b11_OFWNT9L_8tZ[158]\;
    b11_OFWNT9L_8tZ(157) <= \b11_OFWNT9L_8tZ[157]\;
    b11_OFWNT9L_8tZ(156) <= \b11_OFWNT9L_8tZ[156]\;
    b11_OFWNT9L_8tZ(155) <= \b11_OFWNT9L_8tZ[155]\;
    b11_OFWNT9L_8tZ(154) <= \b11_OFWNT9L_8tZ[154]\;
    b11_OFWNT9L_8tZ(153) <= \b11_OFWNT9L_8tZ[153]\;
    b11_OFWNT9L_8tZ(152) <= \b11_OFWNT9L_8tZ[152]\;
    b11_OFWNT9L_8tZ(151) <= \b11_OFWNT9L_8tZ[151]\;
    b11_OFWNT9L_8tZ(150) <= \b11_OFWNT9L_8tZ[150]\;
    b11_OFWNT9L_8tZ(149) <= \b11_OFWNT9L_8tZ[149]\;
    b11_OFWNT9L_8tZ(148) <= \b11_OFWNT9L_8tZ[148]\;
    b11_OFWNT9L_8tZ(147) <= \b11_OFWNT9L_8tZ[147]\;
    b11_OFWNT9L_8tZ(146) <= \b11_OFWNT9L_8tZ[146]\;
    b11_OFWNT9L_8tZ(145) <= \b11_OFWNT9L_8tZ[145]\;
    b11_OFWNT9L_8tZ(144) <= \b11_OFWNT9L_8tZ[144]\;
    b11_OFWNT9L_8tZ(143) <= \b11_OFWNT9L_8tZ[143]\;
    b11_OFWNT9L_8tZ(142) <= \b11_OFWNT9L_8tZ[142]\;
    b11_OFWNT9L_8tZ(141) <= \b11_OFWNT9L_8tZ[141]\;
    b11_OFWNT9L_8tZ(140) <= \b11_OFWNT9L_8tZ[140]\;
    b11_OFWNT9L_8tZ(139) <= \b11_OFWNT9L_8tZ[139]\;
    b11_OFWNT9L_8tZ(138) <= \b11_OFWNT9L_8tZ[138]\;
    b11_OFWNT9L_8tZ(137) <= \b11_OFWNT9L_8tZ[137]\;
    b11_OFWNT9L_8tZ(136) <= \b11_OFWNT9L_8tZ[136]\;
    b11_OFWNT9L_8tZ(135) <= \b11_OFWNT9L_8tZ[135]\;
    b11_OFWNT9L_8tZ(134) <= \b11_OFWNT9L_8tZ[134]\;
    b11_OFWNT9L_8tZ(133) <= \b11_OFWNT9L_8tZ[133]\;
    b11_OFWNT9L_8tZ(132) <= \b11_OFWNT9L_8tZ[132]\;
    b11_OFWNT9L_8tZ(131) <= \b11_OFWNT9L_8tZ[131]\;
    b11_OFWNT9L_8tZ(130) <= \b11_OFWNT9L_8tZ[130]\;
    b11_OFWNT9L_8tZ(129) <= \b11_OFWNT9L_8tZ[129]\;
    b11_OFWNT9L_8tZ(128) <= \b11_OFWNT9L_8tZ[128]\;
    b11_OFWNT9L_8tZ(127) <= \b11_OFWNT9L_8tZ[127]\;
    b11_OFWNT9L_8tZ(126) <= \b11_OFWNT9L_8tZ[126]\;
    b11_OFWNT9L_8tZ(125) <= \b11_OFWNT9L_8tZ[125]\;
    b11_OFWNT9L_8tZ(124) <= \b11_OFWNT9L_8tZ[124]\;
    b11_OFWNT9L_8tZ(123) <= \b11_OFWNT9L_8tZ[123]\;
    b11_OFWNT9L_8tZ(122) <= \b11_OFWNT9L_8tZ[122]\;
    b11_OFWNT9L_8tZ(121) <= \b11_OFWNT9L_8tZ[121]\;
    b11_OFWNT9L_8tZ(120) <= \b11_OFWNT9L_8tZ[120]\;
    b11_OFWNT9L_8tZ(119) <= \b11_OFWNT9L_8tZ[119]\;
    b11_OFWNT9L_8tZ(118) <= \b11_OFWNT9L_8tZ[118]\;
    b11_OFWNT9L_8tZ(117) <= \b11_OFWNT9L_8tZ[117]\;
    b11_OFWNT9L_8tZ(116) <= \b11_OFWNT9L_8tZ[116]\;
    b11_OFWNT9L_8tZ(115) <= \b11_OFWNT9L_8tZ[115]\;
    b11_OFWNT9L_8tZ(114) <= \b11_OFWNT9L_8tZ[114]\;
    b11_OFWNT9L_8tZ(113) <= \b11_OFWNT9L_8tZ[113]\;
    b11_OFWNT9L_8tZ(112) <= \b11_OFWNT9L_8tZ[112]\;
    b11_OFWNT9L_8tZ(111) <= \b11_OFWNT9L_8tZ[111]\;
    b11_OFWNT9L_8tZ(110) <= \b11_OFWNT9L_8tZ[110]\;
    b11_OFWNT9L_8tZ(109) <= \b11_OFWNT9L_8tZ[109]\;
    b11_OFWNT9L_8tZ(108) <= \b11_OFWNT9L_8tZ[108]\;
    b11_OFWNT9L_8tZ(107) <= \b11_OFWNT9L_8tZ[107]\;
    b11_OFWNT9L_8tZ(106) <= \b11_OFWNT9L_8tZ[106]\;
    b11_OFWNT9L_8tZ(105) <= \b11_OFWNT9L_8tZ[105]\;
    b11_OFWNT9L_8tZ(104) <= \b11_OFWNT9L_8tZ[104]\;
    b11_OFWNT9L_8tZ(103) <= \b11_OFWNT9L_8tZ[103]\;
    b11_OFWNT9L_8tZ(102) <= \b11_OFWNT9L_8tZ[102]\;
    b11_OFWNT9L_8tZ(101) <= \b11_OFWNT9L_8tZ[101]\;
    b11_OFWNT9L_8tZ(100) <= \b11_OFWNT9L_8tZ[100]\;
    b11_OFWNT9L_8tZ(99) <= \b11_OFWNT9L_8tZ[99]\;
    b11_OFWNT9L_8tZ(98) <= \b11_OFWNT9L_8tZ[98]\;
    b11_OFWNT9L_8tZ(97) <= \b11_OFWNT9L_8tZ[97]\;
    b11_OFWNT9L_8tZ(96) <= \b11_OFWNT9L_8tZ[96]\;
    b11_OFWNT9L_8tZ(95) <= \b11_OFWNT9L_8tZ[95]\;
    b11_OFWNT9L_8tZ(94) <= \b11_OFWNT9L_8tZ[94]\;
    b11_OFWNT9L_8tZ(93) <= \b11_OFWNT9L_8tZ[93]\;
    b11_OFWNT9L_8tZ(92) <= \b11_OFWNT9L_8tZ[92]\;
    b11_OFWNT9L_8tZ(91) <= \b11_OFWNT9L_8tZ[91]\;
    b11_OFWNT9L_8tZ(90) <= \b11_OFWNT9L_8tZ[90]\;
    b11_OFWNT9L_8tZ(89) <= \b11_OFWNT9L_8tZ[89]\;
    b11_OFWNT9L_8tZ(88) <= \b11_OFWNT9L_8tZ[88]\;
    b11_OFWNT9L_8tZ(87) <= \b11_OFWNT9L_8tZ[87]\;
    b11_OFWNT9L_8tZ(86) <= \b11_OFWNT9L_8tZ[86]\;
    b11_OFWNT9L_8tZ(85) <= \b11_OFWNT9L_8tZ[85]\;
    b11_OFWNT9L_8tZ(84) <= \b11_OFWNT9L_8tZ[84]\;
    b11_OFWNT9L_8tZ(83) <= \b11_OFWNT9L_8tZ[83]\;
    b11_OFWNT9L_8tZ(82) <= \b11_OFWNT9L_8tZ[82]\;
    b11_OFWNT9L_8tZ(81) <= \b11_OFWNT9L_8tZ[81]\;
    b11_OFWNT9L_8tZ(80) <= \b11_OFWNT9L_8tZ[80]\;
    b11_OFWNT9L_8tZ(79) <= \b11_OFWNT9L_8tZ[79]\;
    b11_OFWNT9L_8tZ(78) <= \b11_OFWNT9L_8tZ[78]\;
    b11_OFWNT9L_8tZ(77) <= \b11_OFWNT9L_8tZ[77]\;
    b11_OFWNT9L_8tZ(76) <= \b11_OFWNT9L_8tZ[76]\;
    b11_OFWNT9L_8tZ(75) <= \b11_OFWNT9L_8tZ[75]\;
    b11_OFWNT9L_8tZ(74) <= \b11_OFWNT9L_8tZ[74]\;
    b11_OFWNT9L_8tZ(73) <= \b11_OFWNT9L_8tZ[73]\;
    b11_OFWNT9L_8tZ(72) <= \b11_OFWNT9L_8tZ[72]\;
    b11_OFWNT9L_8tZ(71) <= \b11_OFWNT9L_8tZ[71]\;
    b11_OFWNT9L_8tZ(70) <= \b11_OFWNT9L_8tZ[70]\;
    b11_OFWNT9L_8tZ(69) <= \b11_OFWNT9L_8tZ[69]\;
    b11_OFWNT9L_8tZ(68) <= \b11_OFWNT9L_8tZ[68]\;
    b11_OFWNT9L_8tZ(67) <= \b11_OFWNT9L_8tZ[67]\;
    b11_OFWNT9L_8tZ(66) <= \b11_OFWNT9L_8tZ[66]\;
    b11_OFWNT9L_8tZ(65) <= \b11_OFWNT9L_8tZ[65]\;
    b11_OFWNT9L_8tZ(64) <= \b11_OFWNT9L_8tZ[64]\;
    b11_OFWNT9L_8tZ(63) <= \b11_OFWNT9L_8tZ[63]\;
    b11_OFWNT9L_8tZ(62) <= \b11_OFWNT9L_8tZ[62]\;
    b11_OFWNT9L_8tZ(61) <= \b11_OFWNT9L_8tZ[61]\;
    b11_OFWNT9L_8tZ(60) <= \b11_OFWNT9L_8tZ[60]\;
    b11_OFWNT9L_8tZ(59) <= \b11_OFWNT9L_8tZ[59]\;
    b11_OFWNT9L_8tZ(58) <= \b11_OFWNT9L_8tZ[58]\;
    b11_OFWNT9L_8tZ(57) <= \b11_OFWNT9L_8tZ[57]\;
    b11_OFWNT9L_8tZ(56) <= \b11_OFWNT9L_8tZ[56]\;
    b11_OFWNT9L_8tZ(55) <= \b11_OFWNT9L_8tZ[55]\;
    b11_OFWNT9L_8tZ(54) <= \b11_OFWNT9L_8tZ[54]\;
    b11_OFWNT9L_8tZ(53) <= \b11_OFWNT9L_8tZ[53]\;
    b11_OFWNT9L_8tZ(52) <= \b11_OFWNT9L_8tZ[52]\;
    b11_OFWNT9L_8tZ(51) <= \b11_OFWNT9L_8tZ[51]\;
    b11_OFWNT9L_8tZ(50) <= \b11_OFWNT9L_8tZ[50]\;
    b11_OFWNT9L_8tZ(49) <= \b11_OFWNT9L_8tZ[49]\;
    b11_OFWNT9L_8tZ(48) <= \b11_OFWNT9L_8tZ[48]\;
    b11_OFWNT9L_8tZ(47) <= \b11_OFWNT9L_8tZ[47]\;
    b11_OFWNT9L_8tZ(46) <= \b11_OFWNT9L_8tZ[46]\;
    b11_OFWNT9L_8tZ(45) <= \b11_OFWNT9L_8tZ[45]\;
    b11_OFWNT9L_8tZ(44) <= \b11_OFWNT9L_8tZ[44]\;
    b11_OFWNT9L_8tZ(43) <= \b11_OFWNT9L_8tZ[43]\;
    b11_OFWNT9L_8tZ(42) <= \b11_OFWNT9L_8tZ[42]\;
    b11_OFWNT9L_8tZ(41) <= \b11_OFWNT9L_8tZ[41]\;
    b11_OFWNT9L_8tZ(40) <= \b11_OFWNT9L_8tZ[40]\;
    b11_OFWNT9L_8tZ(39) <= \b11_OFWNT9L_8tZ[39]\;
    b11_OFWNT9L_8tZ(38) <= \b11_OFWNT9L_8tZ[38]\;
    b11_OFWNT9L_8tZ(37) <= \b11_OFWNT9L_8tZ[37]\;
    b11_OFWNT9L_8tZ(36) <= \b11_OFWNT9L_8tZ[36]\;
    b11_OFWNT9L_8tZ(35) <= \b11_OFWNT9L_8tZ[35]\;
    b11_OFWNT9L_8tZ(34) <= \b11_OFWNT9L_8tZ[34]\;
    b11_OFWNT9L_8tZ(33) <= \b11_OFWNT9L_8tZ[33]\;
    b11_OFWNT9L_8tZ(32) <= \b11_OFWNT9L_8tZ[32]\;
    b11_OFWNT9L_8tZ(31) <= \b11_OFWNT9L_8tZ[31]\;
    b11_OFWNT9L_8tZ(30) <= \b11_OFWNT9L_8tZ[30]\;
    b11_OFWNT9L_8tZ(29) <= \b11_OFWNT9L_8tZ[29]\;
    b11_OFWNT9L_8tZ(28) <= \b11_OFWNT9L_8tZ[28]\;
    b11_OFWNT9L_8tZ(27) <= \b11_OFWNT9L_8tZ[27]\;
    b11_OFWNT9L_8tZ(26) <= \b11_OFWNT9L_8tZ[26]\;
    b11_OFWNT9L_8tZ(25) <= \b11_OFWNT9L_8tZ[25]\;
    b11_OFWNT9L_8tZ(24) <= \b11_OFWNT9L_8tZ[24]\;
    b11_OFWNT9L_8tZ(23) <= \b11_OFWNT9L_8tZ[23]\;
    b11_OFWNT9L_8tZ(22) <= \b11_OFWNT9L_8tZ[22]\;
    b11_OFWNT9L_8tZ(21) <= \b11_OFWNT9L_8tZ[21]\;
    b11_OFWNT9L_8tZ(20) <= \b11_OFWNT9L_8tZ[20]\;
    b11_OFWNT9L_8tZ(19) <= \b11_OFWNT9L_8tZ[19]\;
    b11_OFWNT9L_8tZ(18) <= \b11_OFWNT9L_8tZ[18]\;
    b11_OFWNT9L_8tZ(17) <= \b11_OFWNT9L_8tZ[17]\;
    b11_OFWNT9L_8tZ(16) <= \b11_OFWNT9L_8tZ[16]\;
    b11_OFWNT9L_8tZ(15) <= \b11_OFWNT9L_8tZ[15]\;
    b11_OFWNT9L_8tZ(14) <= \b11_OFWNT9L_8tZ[14]\;
    b11_OFWNT9L_8tZ(13) <= \b11_OFWNT9L_8tZ[13]\;
    b11_OFWNT9L_8tZ(12) <= \b11_OFWNT9L_8tZ[12]\;
    b11_OFWNT9L_8tZ(11) <= \b11_OFWNT9L_8tZ[11]\;
    b11_OFWNT9L_8tZ(10) <= \b11_OFWNT9L_8tZ[10]\;
    b11_OFWNT9L_8tZ(9) <= \b11_OFWNT9L_8tZ[9]\;
    b11_OFWNT9L_8tZ(8) <= \b11_OFWNT9L_8tZ[8]\;
    b11_OFWNT9L_8tZ(7) <= \b11_OFWNT9L_8tZ[7]\;
    b11_OFWNT9L_8tZ(6) <= \b11_OFWNT9L_8tZ[6]\;
    b11_OFWNT9L_8tZ(5) <= \b11_OFWNT9L_8tZ[5]\;
    b11_OFWNT9L_8tZ(4) <= \b11_OFWNT9L_8tZ[4]\;
    b11_OFWNT9L_8tZ(3) <= \b11_OFWNT9L_8tZ[3]\;
    b11_OFWNT9L_8tZ(2) <= \b11_OFWNT9L_8tZ[2]\;
    b11_OFWNT9L_8tZ(1) <= \b11_OFWNT9L_8tZ[1]\;
    b11_OFWNT9L_8tZ(0) <= \b11_OFWNT9L_8tZ[0]\;

    \genblk9.b3_PfG_RNO[101]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[102]\, C => 
        \b7_vFW_PlM[100]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[101]\);
    
    \genblk9.b7_nYJ_BFM[34]\ : SLE
      port map(D => \b7_nYJ_BFM[33]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[34]\);
    
    \genblk9.b3_PfG_RNO[61]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[62]\, C => 
        \b7_vFW_PlM[60]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[61]\);
    
    \genblk9.b3_PfG[14]\ : SLE
      port map(D => \b3_PfG_6[14]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[14]\);
    
    \genblk9.b3_PfG_RNO[60]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[61]\, C => 
        \b7_vFW_PlM[59]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[60]\);
    
    \genblk9.b3_PfG[2]\ : SLE
      port map(D => \b3_PfG_6[2]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[2]\);
    
    \genblk9.b3_PfG_RNO[104]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[105]\, C => 
        \b7_vFW_PlM[103]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[104]\);
    
    \genblk9.b7_nYJ_BFM[48]\ : SLE
      port map(D => \b7_nYJ_BFM[47]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[48]\);
    
    \genblk9.b3_PfG_RNO[41]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[42]\, C => 
        \b7_vFW_PlM[40]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[41]\);
    
    \genblk9.b3_PfG_RNO[57]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[58]\, C => 
        \b7_vFW_PlM[56]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[57]\);
    
    \genblk9.b3_PfG_RNO[139]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[140]\, C => 
        \b7_vFW_PlM[138]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[139]\);
    
    \genblk9.b3_PfG_RNO[40]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[41]\, C => 
        \b7_vFW_PlM[39]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[40]\);
    
    \genblk9.b3_PfG_RNO[133]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[134]\, C => 
        \b7_vFW_PlM[132]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[133]\);
    
    \genblk9.b3_PfG_RNO[92]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[93]\, C => 
        \b7_vFW_PlM[91]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[92]\);
    
    \genblk9.b3_PfG[6]\ : SLE
      port map(D => \b3_PfG_6[6]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[6]\);
    
    \genblk9.b7_nYJ_BFM[158]\ : SLE
      port map(D => \b7_nYJ_BFM[157]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[158]\);
    
    \genblk9.b7_nYJ_BFM[27]\ : SLE
      port map(D => \b7_nYJ_BFM[26]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[27]\);
    
    \genblk9.b9_v_mzCDYXs[3]\ : SLE
      port map(D => \b9_v_mzCDYXs_s[3]\, CLK => 
        IICE_comm2iice(11), EN => b9_v_mzCDYXs13, ALn => 
        b5_voSc3_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \b9_v_mzCDYXs[3]\);
    
    \genblk9.b3_PfG[116]\ : SLE
      port map(D => \b3_PfG_6[116]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[116]\);
    
    \genblk9.b7_nYJ_BFM[95]\ : SLE
      port map(D => \b7_nYJ_BFM[94]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[95]\);
    
    \genblk9.b7_nYJ_BFM[167]\ : SLE
      port map(D => \b7_nYJ_BFM[166]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[167]\);
    
    \genblk9.b7_nYJ_BFM[147]\ : SLE
      port map(D => \b7_nYJ_BFM[146]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[147]\);
    
    \genblk9.b7_nYJ_BFM[71]\ : SLE
      port map(D => \b7_nYJ_BFM[70]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[71]\);
    
    \genblk9.b3_PfG_RNO[109]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[110]\, C => 
        \b7_vFW_PlM[108]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[109]\);
    
    \genblk9.b3_PfG_RNO[6]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[7]\, C => 
        \b7_vFW_PlM[5]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[6]\);
    
    \genblk9.b3_PfG_RNO[103]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[104]\, C => 
        \b7_vFW_PlM[102]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[103]\);
    
    \genblk9.b3_PfG[131]\ : SLE
      port map(D => \b3_PfG_6[131]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[131]\);
    
    \genblk9.b7_nYJ_BFM[61]\ : SLE
      port map(D => \b7_nYJ_BFM[60]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[61]\);
    
    \genblk9.b3_PfG[90]\ : SLE
      port map(D => \b3_PfG_6[90]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[90]\);
    
    \genblk9.b3_PfG[78]\ : SLE
      port map(D => \b3_PfG_6[78]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[78]\);
    
    \genblk9.b3_PfG[11]\ : SLE
      port map(D => \b3_PfG_6[11]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[11]\);
    
    \genblk9.b3_PfG[127]\ : SLE
      port map(D => \b3_PfG_6[127]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[127]\);
    
    \genblk9.b9_v_mzCDYXs[2]\ : SLE
      port map(D => \b9_v_mzCDYXs_s[2]\, CLK => 
        IICE_comm2iice(11), EN => b9_v_mzCDYXs13, ALn => 
        b5_voSc3_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \b9_v_mzCDYXs[2]\);
    
    \genblk9.b7_nYJ_BFM[80]\ : SLE
      port map(D => \b7_nYJ_BFM[79]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[80]\);
    
    \genblk9.b9_v_mzCDYXs_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \b9_v_mzCDYXs[2]\, C => 
        GND_net_1, D => GND_net_1, FCI => \b9_v_mzCDYXs_cry[1]\, 
        S => \b9_v_mzCDYXs_s[2]\, Y => OPEN, FCO => 
        \b9_v_mzCDYXs_cry[2]\);
    
    \genblk9.b3_PfG_RNO[150]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[151]\, C => 
        \b7_vFW_PlM[149]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[150]\);
    
    \genblk9.b3_PfG[34]\ : SLE
      port map(D => \b3_PfG_6[34]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[34]\);
    
    \genblk9.b3_PfG[107]\ : SLE
      port map(D => \b3_PfG_6[107]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[107]\);
    
    \genblk9.b7_nYJ_BFM[120]\ : SLE
      port map(D => \b7_nYJ_BFM[119]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[120]\);
    
    \genblk9.b3_PfG[68]\ : SLE
      port map(D => \b3_PfG_6[68]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[68]\);
    
    \genblk9.b3_PfG[145]\ : SLE
      port map(D => \b3_PfG_6[145]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[145]\);
    
    \b12_PSyi_KyDbLbb[7]\ : SLE
      port map(D => \b12_2_St6KCa_jHv[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \b12_PSyi_KyDbLbb_0_sqmuxa\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \b12_PSyi_KyDbLbb[7]_net_1\);
    
    \genblk9.b7_nYJ_BFM[91]\ : SLE
      port map(D => \b7_nYJ_BFM[90]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[91]\);
    
    \genblk9.b3_PfG[136]\ : SLE
      port map(D => \b3_PfG_6[136]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[136]\);
    
    \genblk9.b3_PfG_RNO[28]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[29]\, C => 
        \b7_vFW_PlM[27]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[28]\);
    
    \genblk9.b7_nYJ_BFM[170]\ : SLE
      port map(D => \b7_nYJ_BFM[169]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[170]\);
    
    \genblk9.b7_nYJ_BFM[56]\ : SLE
      port map(D => \b7_nYJ_BFM[55]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[56]\);
    
    \genblk9.b7_nYJ_BFM[12]\ : SLE
      port map(D => \b7_nYJ_BFM[11]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[12]\);
    
    \genblk9.b3_PfG_RNO[93]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[94]\, C => 
        \b7_vFW_PlM[92]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[93]\);
    
    \genblk9.b3_PfG[25]\ : SLE
      port map(D => \b3_PfG_6[25]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[25]\);
    
    \genblk9.b3_PfG_RNO[12]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[13]\, C => 
        \b7_vFW_PlM[11]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[12]\);
    
    \genblk9.b3_PfG[151]\ : SLE
      port map(D => \b3_PfG_6[151]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[151]\);
    
    \genblk9.b7_nYJ_BFM[36]\ : SLE
      port map(D => \b7_nYJ_BFM[35]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[36]\);
    
    \b12_2_St6KCa_jHv_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \b12_2_St6KCa_jHv[0]_net_1\, Y => 
        \b12_2_St6KCa_jHv_s[0]\);
    
    \genblk9.b3_PfG[31]\ : SLE
      port map(D => \b3_PfG_6[31]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[31]\);
    
    \genblk9.b3_PfG_RNO[86]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[87]\, C => 
        \b7_vFW_PlM[85]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[86]\);
    
    \genblk9.b7_nYJ_BFM[110]\ : SLE
      port map(D => \b7_nYJ_BFM[109]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[110]\);
    
    \genblk9.b3_PfG_RNO[31]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[32]\, C => 
        \b7_vFW_PlM[30]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[31]\);
    
    \genblk9.b3_PfG_RNO[68]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[69]\, C => 
        \b7_vFW_PlM[67]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[68]\);
    
    \genblk9.b3_PfG_RNO[30]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[31]\, C => 
        \b7_vFW_PlM[29]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[30]\);
    
    \genblk9.b7_nYJ_BFM[161]\ : SLE
      port map(D => \b7_nYJ_BFM[160]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[161]\);
    
    \b12_2_St6KCa_jHv[5]\ : SLE
      port map(D => \b12_2_St6KCa_jHv_s[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b4_2o_z, ALn => b5_voSc3_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b12_2_St6KCa_jHv[5]_net_1\);
    
    \genblk9.b9_v_mzCDYXs[4]\ : SLE
      port map(D => \b9_v_mzCDYXs_s[4]\, CLK => 
        IICE_comm2iice(11), EN => b9_v_mzCDYXs13, ALn => 
        b5_voSc3_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \b9_v_mzCDYXs[4]\);
    
    \genblk9.b7_nYJ_BFM[141]\ : SLE
      port map(D => \b7_nYJ_BFM[140]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[141]\);
    
    \genblk9.b3_PfG[165]\ : SLE
      port map(D => \b3_PfG_6[165]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[165]\);
    
    \genblk9.b3_PfG[40]\ : SLE
      port map(D => \b3_PfG_6[40]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[40]\);
    
    \genblk9.b3_PfG_RNO[48]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[49]\, C => 
        \b7_vFW_PlM[47]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[48]\);
    
    \genblk9.b3_PfG[16]\ : SLE
      port map(D => \b3_PfG_6[16]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[16]\);
    
    \genblk9.b3_PfG[122]\ : SLE
      port map(D => \b3_PfG_6[122]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[122]\);
    
    \genblk9.b3_PfG[77]\ : SLE
      port map(D => \b3_PfG_6[77]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[77]\);
    
    \genblk9.b3_PfG[143]\ : SLE
      port map(D => \b3_PfG_6[143]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[143]\);
    
    \b8_FZFFLXYE[4]\ : SLE
      port map(D => \b12_2_St6KCa_jHv[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b4_2o_z, ALn => b5_voSc3_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b8_FZFFLXYE[4]_net_1\);
    
    \genblk9.b3_PfG[156]\ : SLE
      port map(D => \b3_PfG_6[156]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[156]\);
    
    \b8_FZFFLXYE[0]\ : SLE
      port map(D => \b12_2_St6KCa_jHv[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b4_2o_z, ALn => b5_voSc3_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b8_FZFFLXYE[0]_net_1\);
    
    \genblk9.b9_v_mzCDYXs[7]\ : SLE
      port map(D => \b9_v_mzCDYXs_s[7]\, CLK => 
        IICE_comm2iice(11), EN => b9_v_mzCDYXs13, ALn => 
        b5_voSc3_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \b9_v_mzCDYXs[7]\);
    
    \genblk9.b3_PfG[102]\ : SLE
      port map(D => \b3_PfG_6[102]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[102]\);
    
    \genblk9.b3_PfG[54]\ : SLE
      port map(D => \b3_PfG_6[54]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[54]\);
    
    \genblk9.b3_PfG[140]\ : SLE
      port map(D => \b3_PfG_6[140]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[140]\);
    
    \genblk9.b3_PfG[67]\ : SLE
      port map(D => \b3_PfG_6[67]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[67]\);
    
    \b8_FZFFLXYE[2]\ : SLE
      port map(D => \b12_2_St6KCa_jHv[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b4_2o_z, ALn => b5_voSc3_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b8_FZFFLXYE[2]_net_1\);
    
    \genblk9.b11_nFG0rDY_9e2\ : SLE
      port map(D => b11_nFG0rDY_9e2_2, CLK => IICE_comm2iice(11), 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_nFG0rDY_9e2);
    
    \b8_FZFFLXYE[8]\ : SLE
      port map(D => \b12_2_St6KCa_jHv[8]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b4_2o_z, ALn => b5_voSc3_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b8_FZFFLXYE[8]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \genblk9.b7_nYJ_BFM[25]\ : SLE
      port map(D => \b7_nYJ_BFM[24]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[25]\);
    
    \genblk9.b7_nYJ_BFM[166]\ : SLE
      port map(D => \b7_nYJ_BFM[165]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[166]\);
    
    \genblk9.b3_PfG[85]\ : SLE
      port map(D => \b3_PfG_6[85]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[85]\);
    
    \genblk9.b7_nYJ_BFM[146]\ : SLE
      port map(D => \b7_nYJ_BFM[145]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[146]\);
    
    \genblk9.b7_nYJ_BFM[129]\ : SLE
      port map(D => \b7_nYJ_BFM[128]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[129]\);
    
    \genblk9.b7_nYJ_BFM[72]\ : SLE
      port map(D => \b7_nYJ_BFM[71]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[72]\);
    
    \genblk9.b3_PfG_RNO[97]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[98]\, C => 
        \b7_vFW_PlM[96]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[97]\);
    
    \genblk9.b7_nYJ_BFM[130]\ : SLE
      port map(D => \b7_nYJ_BFM[129]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[130]\);
    
    \genblk9.b3_PfG_RNO[13]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[14]\, C => 
        \b7_vFW_PlM[12]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[13]\);
    
    \genblk9.b3_PfG_RNO[1]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[2]\, C => 
        \b7_vFW_PlM[0]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[1]\);
    
    \genblk9.b7_nYJ_BFM[83]\ : SLE
      port map(D => \b7_nYJ_BFM[82]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[83]\);
    
    \genblk9.b3_PfG[163]\ : SLE
      port map(D => \b3_PfG_6[163]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[163]\);
    
    \genblk9.b3_PfG[36]\ : SLE
      port map(D => \b3_PfG_6[36]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[36]\);
    
    \genblk9.b7_nYJ_BFM[19]\ : SLE
      port map(D => \b7_nYJ_BFM[18]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[19]\);
    
    \genblk9.b3_PfG[72]\ : SLE
      port map(D => \b3_PfG_6[72]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[72]\);
    
    \genblk9.b7_nYJ_BFM[62]\ : SLE
      port map(D => \b7_nYJ_BFM[61]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[62]\);
    
    \b12_2_St6KCa_jHv[0]\ : SLE
      port map(D => \b12_2_St6KCa_jHv_s[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b4_2o_z, ALn => b5_voSc3_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b12_2_St6KCa_jHv[0]_net_1\);
    
    \genblk9.b3_PfG_RNO[76]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[77]\, C => 
        \b7_vFW_PlM[75]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[76]\);
    
    \b12_2_St6KCa_jHv[6]\ : SLE
      port map(D => \b12_2_St6KCa_jHv_s[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b4_2o_z, ALn => b5_voSc3_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b12_2_St6KCa_jHv[6]_net_1\);
    
    \b12_2_St6KCa_jHv_s[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \b12_2_St6KCa_jHv[11]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \b12_2_St6KCa_jHv_cry[10]_net_1\, S => 
        \b12_2_St6KCa_jHv_s[11]_net_1\, Y => OPEN, FCO => OPEN);
    
    \genblk9.b3_PfG_RNO[165]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[166]\, C => 
        \b7_vFW_PlM[164]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[165]\);
    
    \genblk9.b3_PfG[51]\ : SLE
      port map(D => \b3_PfG_6[51]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[51]\);
    
    \genblk9.b3_PfG_RNO[85]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[86]\, C => 
        \b7_vFW_PlM[84]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[85]\);
    
    b9_PSyil9s_2 : SLE
      port map(D => b13_wRBtT_ME83hHx, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b9_PSyil9s_2\);
    
    \genblk9.b3_PfG[79]\ : SLE
      port map(D => \b3_PfG_6[79]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[79]\);
    
    \genblk9.b3_PfG[160]\ : SLE
      port map(D => \b3_PfG_6[160]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[160]\);
    
    \genblk9.b7_nYJ_BFM[40]\ : SLE
      port map(D => \b7_nYJ_BFM[39]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[40]\);
    
    \genblk9.b7_nYJ_BFM[57]\ : SLE
      port map(D => \b7_nYJ_BFM[56]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[57]\);
    
    \genblk9.b7_nYJ_BFM[125]\ : SLE
      port map(D => \b7_nYJ_BFM[124]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[125]\);
    
    \genblk9.b3_PfG[62]\ : SLE
      port map(D => \b3_PfG_6[62]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[62]\);
    
    \genblk9.b7_nYJ_BFM[119]\ : SLE
      port map(D => \b7_nYJ_BFM[118]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[119]\);
    
    \genblk9.b7_nYJ_BFM[123]\ : SLE
      port map(D => \b7_nYJ_BFM[122]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[123]\);
    
    \b12_2_St6KCa_jHv_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \b12_2_St6KCa_jHv[1]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        b12_2_St6KCa_jHv_s_900_FCO, S => \b12_2_St6KCa_jHv_s[1]\, 
        Y => OPEN, FCO => \b12_2_St6KCa_jHv_cry[1]_net_1\);
    
    \genblk9.b7_nYJ_BFM[37]\ : SLE
      port map(D => \b7_nYJ_BFM[36]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[37]\);
    
    \genblk9.b3_PfG_RNO[161]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[162]\, C => 
        \b7_vFW_PlM[160]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[161]\);
    
    \genblk9.b7_nYJ_BFM[21]\ : SLE
      port map(D => \b7_nYJ_BFM[20]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[21]\);
    
    \b8_FZFFLXYE[11]\ : SLE
      port map(D => \b12_2_St6KCa_jHv[11]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b4_2o_z, ALn => b5_voSc3_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b8_FZFFLXYE[11]_net_1\);
    
    \genblk9.b7_nYJ_BFM[84]\ : SLE
      port map(D => \b7_nYJ_BFM[83]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[84]\);
    
    \b12_2_St6KCa_jHv_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \b12_2_St6KCa_jHv[3]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \b12_2_St6KCa_jHv_cry[2]_net_1\, S => 
        \b12_2_St6KCa_jHv_s[3]\, Y => OPEN, FCO => 
        \b12_2_St6KCa_jHv_cry[3]_net_1\);
    
    \genblk9.b7_nYJ_BFM[92]\ : SLE
      port map(D => \b7_nYJ_BFM[91]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[92]\);
    
    \genblk9.b3_PfG[69]\ : SLE
      port map(D => \b3_PfG_6[69]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[69]\);
    
    \genblk9.b7_nYJ_BFM[18]\ : SLE
      port map(D => \b7_nYJ_BFM[17]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[18]\);
    
    \genblk9.b7_nYJ_BFM[173]\ : SLE
      port map(D => \b7_nYJ_BFM[172]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[173]\);
    
    \genblk9.b3_PfG_RNO[38]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[39]\, C => 
        \b7_vFW_PlM[37]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[38]\);
    
    \b12_PSyi_KyDbLbb[11]\ : SLE
      port map(D => \b12_2_St6KCa_jHv[11]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \b12_PSyi_KyDbLbb_0_sqmuxa\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \b12_PSyi_KyDbLbb[11]_net_1\);
    
    \genblk9.b3_PfG_RNO[164]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[165]\, C => 
        \b7_vFW_PlM[163]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[164]\);
    
    \genblk9.b9_v_mzCDYXs[1]\ : SLE
      port map(D => \b9_v_mzCDYXs_s[1]\, CLK => 
        IICE_comm2iice(11), EN => b9_v_mzCDYXs13, ALn => 
        b5_voSc3_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \b9_v_mzCDYXs[1]\);
    
    \genblk9.b7_nYJ_BFM[124]\ : SLE
      port map(D => \b7_nYJ_BFM[123]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[124]\);
    
    \genblk9.b3_PfG_RNO[156]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[157]\, C => 
        \b7_vFW_PlM[155]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[156]\);
    
    \genblk9.b3_PfG[9]\ : SLE
      port map(D => \b3_PfG_6[9]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[9]\);
    
    \genblk9.b3_PfG[94]\ : SLE
      port map(D => \b3_PfG_6[94]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[94]\);
    
    \genblk9.b7_nYJ_BFM[107]\ : SLE
      port map(D => \b7_nYJ_BFM[106]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[107]\);
    
    \genblk9.b9_v_mzCDYXs_s_901\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \b9_v_mzCDYXs[0]\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => b9_v_mzCDYXs_s_901_FCO);
    
    \genblk9.b7_nYJ_BFM[115]\ : SLE
      port map(D => \b7_nYJ_BFM[114]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[115]\);
    
    N_15_i : CFG2
      generic map(INIT => x"8")

      port map(A => b9_OFWNT9_ab, B => IICE_comm2iice(10), Y => 
        \N_15_i\);
    
    \genblk9.b7_nYJ_BFM[174]\ : SLE
      port map(D => \b7_nYJ_BFM[173]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[174]\);
    
    \b12_2_St6KCa_jHv[10]\ : SLE
      port map(D => \b12_2_St6KCa_jHv_s[10]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b4_2o_z, ALn => b5_voSc3_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b12_2_St6KCa_jHv[10]_net_1\);
    
    \genblk9.b7_nYJ_BFM[113]\ : SLE
      port map(D => \b7_nYJ_BFM[112]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[113]\);
    
    \genblk9.b3_PfG_RNO[17]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[18]\, C => 
        \b7_vFW_PlM[16]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[17]\);
    
    \genblk9.b3_PfG[121]\ : SLE
      port map(D => \b3_PfG_6[121]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[121]\);
    
    \genblk9.b3_PfG[18]\ : SLE
      port map(D => \b3_PfG_6[18]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[18]\);
    
    \genblk9.b3_PfG_RNO[145]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[146]\, C => 
        \b7_vFW_PlM[144]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[145]\);
    
    \genblk9.b3_PfG_RNO[163]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[164]\, C => 
        \b7_vFW_PlM[162]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[163]\);
    
    \genblk9.b3_PfG_RNO[4]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[5]\, C => 
        \b7_vFW_PlM[3]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[4]\);
    
    \genblk9.b3_PfG_RNO[56]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[57]\, C => 
        \b7_vFW_PlM[55]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[56]\);
    
    \genblk9.b3_PfG_RNO[22]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[23]\, C => 
        \b7_vFW_PlM[21]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[22]\);
    
    \genblk9.b9_v_mzCDYXs_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \b9_v_mzCDYXs[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => \b9_v_mzCDYXs_cry[3]\, 
        S => \b9_v_mzCDYXs_s[4]\, Y => OPEN, FCO => 
        \b9_v_mzCDYXs_cry[4]\);
    
    \genblk9.b9_v_mzCDYXs[0]\ : SLE
      port map(D => \b9_v_mzCDYXs_s[0]\, CLK => 
        IICE_comm2iice(11), EN => b9_v_mzCDYXs13, ALn => 
        b5_voSc3_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \b9_v_mzCDYXs[0]\);
    
    \genblk9.b7_nYJ_BFM[79]\ : SLE
      port map(D => \b7_nYJ_BFM[78]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[79]\);
    
    \genblk9.b3_PfG_RNO[7]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[8]\, C => 
        \b7_vFW_PlM[6]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[7]\);
    
    \genblk9.b3_PfG_RNO[132]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[133]\, C => 
        \b7_vFW_PlM[131]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[132]\);
    
    \genblk9.b3_PfG[56]\ : SLE
      port map(D => \b3_PfG_6[56]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[56]\);
    
    \genblk9.b3_PfG[101]\ : SLE
      port map(D => \b3_PfG_6[101]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[101]\);
    
    \genblk9.b3_PfG[73]\ : SLE
      port map(D => \b3_PfG_6[73]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[73]\);
    
    \genblk9.b7_nYJ_BFM[139]\ : SLE
      port map(D => \b7_nYJ_BFM[138]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[139]\);
    
    \genblk9.b7_nYJ_BFM[114]\ : SLE
      port map(D => \b7_nYJ_BFM[113]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[114]\);
    
    b7_yYh03wy4_0_a2_0_2 : CFG3
      generic map(INIT => x"20")

      port map(A => IICE_comm2iice(0), B => IICE_comm2iice(3), C
         => IICE_comm2iice(1), Y => \b7_yYh03wy4_0_a2_0_2\);
    
    \genblk9.b7_nYJ_BFM[69]\ : SLE
      port map(D => \b7_nYJ_BFM[68]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[69]\);
    
    \genblk9.b7_nYJ_BFM[122]\ : SLE
      port map(D => \b7_nYJ_BFM[121]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[122]\);
    
    \b12_PSyi_KyDbLbb[9]\ : SLE
      port map(D => \b12_2_St6KCa_jHv[9]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \b12_PSyi_KyDbLbb_0_sqmuxa\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \b12_PSyi_KyDbLbb[9]_net_1\);
    
    \genblk9.b3_PfG_RNO[141]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[142]\, C => 
        \b7_vFW_PlM[140]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[141]\);
    
    \genblk9.b3_PfG_RNO[75]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[76]\, C => 
        \b7_vFW_PlM[74]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[75]\);
    
    \genblk9.b3_PfG[91]\ : SLE
      port map(D => \b3_PfG_6[91]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[91]\);
    
    \genblk9.b3_PfG[144]\ : SLE
      port map(D => \b3_PfG_6[144]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[144]\);
    
    \genblk9.b3_PfG_RNO[125]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[126]\, C => 
        \b7_vFW_PlM[124]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[125]\);
    
    b8_jAA_KlCO_0_sqmuxa_7 : CFG4
      generic map(INIT => x"8000")

      port map(A => \b12_2_St6KCa_jHv[11]_net_1\, B => 
        \b12_2_St6KCa_jHv[10]_net_1\, C => 
        \b12_2_St6KCa_jHv[9]_net_1\, D => 
        \b12_2_St6KCa_jHv[8]_net_1\, Y => 
        \b8_jAA_KlCO_0_sqmuxa_7\);
    
    \b8_FZFFLXYE[3]\ : SLE
      port map(D => \b12_2_St6KCa_jHv[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b4_2o_z, ALn => b5_voSc3_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b8_FZFFLXYE[3]_net_1\);
    
    \b12_2_St6KCa_jHv_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \b12_2_St6KCa_jHv[8]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \b12_2_St6KCa_jHv_cry[7]_net_1\, S => 
        \b12_2_St6KCa_jHv_s[8]\, Y => OPEN, FCO => 
        \b12_2_St6KCa_jHv_cry[8]_net_1\);
    
    \genblk9.b3_PfG_RNO[102]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[103]\, C => 
        \b7_vFW_PlM[101]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[102]\);
    
    \b8_FZFFLXYE[7]\ : SLE
      port map(D => \b12_2_St6KCa_jHv[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b4_2o_z, ALn => b5_voSc3_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b8_FZFFLXYE[7]_net_1\);
    
    \genblk9.b3_PfG[63]\ : SLE
      port map(D => \b3_PfG_6[63]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[63]\);
    
    \genblk9.b3_PfG[126]\ : SLE
      port map(D => \b3_PfG_6[126]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[126]\);
    
    \genblk9.b7_nYJ_BFM[172]\ : SLE
      port map(D => \b7_nYJ_BFM[171]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[172]\);
    
    \genblk9.b3_PfG_RNO[144]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[145]\, C => 
        \b7_vFW_PlM[143]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[144]\);
    
    \genblk9.b3_PfG_RNO[9]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[10]\, C => 
        \b7_vFW_PlM[8]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[9]\);
    
    \genblk9.b3_PfG[20]\ : SLE
      port map(D => \b3_PfG_6[20]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[20]\);
    
    \genblk9.b3_PfG_RNO[62]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[63]\, C => 
        \b7_vFW_PlM[61]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[62]\);
    
    \genblk9.b3_PfG_RNO[89]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[90]\, C => 
        \b7_vFW_PlM[88]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[89]\);
    
    \genblk9.b3_PfG_RNO[138]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[139]\, C => 
        \b7_vFW_PlM[137]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[138]\);
    
    \b12_2_St6KCa_jHv[4]\ : SLE
      port map(D => \b12_2_St6KCa_jHv_s[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b4_2o_z, ALn => b5_voSc3_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b12_2_St6KCa_jHv[4]_net_1\);
    
    \genblk9.b3_PfG_RNO[121]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[122]\, C => 
        \b7_vFW_PlM[120]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[121]\);
    
    \genblk9.b7_nYJ_BFM[78]\ : SLE
      port map(D => \b7_nYJ_BFM[77]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[78]\);
    
    \genblk9.b7_nYJ_BFM[135]\ : SLE
      port map(D => \b7_nYJ_BFM[134]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[135]\);
    
    \genblk9.b3_PfG_RNO[42]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[43]\, C => 
        \b7_vFW_PlM[41]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[42]\);
    
    \genblk9.b3_PfG_RNO[137]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[138]\, C => 
        \b7_vFW_PlM[136]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[137]\);
    
    \genblk9.b3_PfG[106]\ : SLE
      port map(D => \b3_PfG_6[106]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[106]\);
    
    \genblk9.b3_PfG[38]\ : SLE
      port map(D => \b3_PfG_6[38]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[38]\);
    
    \genblk9.b7_nYJ_BFM[99]\ : SLE
      port map(D => \b7_nYJ_BFM[98]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[99]\);
    
    \genblk9.b7_nYJ_BFM[133]\ : SLE
      port map(D => \b7_nYJ_BFM[132]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[133]\);
    
    \genblk9.b3_PfG[44]\ : SLE
      port map(D => \b3_PfG_6[44]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[44]\);
    
    \genblk9.b3_PfG_RNO[149]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[150]\, C => 
        \b7_vFW_PlM[148]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[149]\);
    
    \genblk9.b7_nYJ_BFM[112]\ : SLE
      port map(D => \b7_nYJ_BFM[111]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[112]\);
    
    \genblk9.b7_nYJ_BFM[68]\ : SLE
      port map(D => \b7_nYJ_BFM[67]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[68]\);
    
    \genblk9.b7_nYJ_BFM[43]\ : SLE
      port map(D => \b7_nYJ_BFM[42]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[43]\);
    
    \genblk9.b3_PfG_RNO[124]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[125]\, C => 
        \b7_vFW_PlM[123]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[124]\);
    
    \genblk9.b3_PfG_RNO[143]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[144]\, C => 
        \b7_vFW_PlM[142]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[143]\);
    
    \genblk9.b3_PfG_RNO[108]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[109]\, C => 
        \b7_vFW_PlM[107]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[108]\);
    
    \genblk9.b3_PfG[115]\ : SLE
      port map(D => \b3_PfG_6[115]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[115]\);
    
    \genblk9.b7_nYJ_BFM[86]\ : SLE
      port map(D => \b7_nYJ_BFM[85]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[86]\);
    
    \genblk9.b3_PfG_RNO[84]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[85]\, C => 
        \b7_vFW_PlM[83]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[84]\);
    
    \b12_PSyi_KyDbLbb[6]\ : SLE
      port map(D => \b12_2_St6KCa_jHv[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \b12_PSyi_KyDbLbb_0_sqmuxa\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \b12_PSyi_KyDbLbb[6]_net_1\);
    
    \genblk9.b3_PfG_RNO[107]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[108]\, C => 
        \b7_vFW_PlM[106]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[107]\);
    
    \genblk9.b3_PfG[148]\ : SLE
      port map(D => \b3_PfG_6[148]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[148]\);
    
    \genblk9.b9_v_mzCDYXs_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \b9_v_mzCDYXs[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => \b9_v_mzCDYXs_cry[4]\, 
        S => \b9_v_mzCDYXs_s[5]\, Y => OPEN, FCO => 
        \b9_v_mzCDYXs_cry[5]\);
    
    \genblk9.b3_PfG[164]\ : SLE
      port map(D => \b3_PfG_6[164]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[164]\);
    
    \genblk9.b7_nYJ_BFM[134]\ : SLE
      port map(D => \b7_nYJ_BFM[133]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[134]\);
    
    \genblk9.b7_nYJ_BFM[157]\ : SLE
      port map(D => \b7_nYJ_BFM[156]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[157]\);
    
    \genblk9.b3_PfG_RNO[23]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[24]\, C => 
        \b7_vFW_PlM[22]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[23]\);
    
    \genblk9.b3_PfG[17]\ : SLE
      port map(D => \b3_PfG_6[17]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[17]\);
    
    \genblk9.b7_nYJ_BFM[101]\ : SLE
      port map(D => \b7_nYJ_BFM[100]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[101]\);
    
    \genblk9.b7_nYJ_BFM[1]\ : SLE
      port map(D => \b7_nYJ_BFM[0]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[1]\);
    
    \genblk9.b3_PfG[5]\ : SLE
      port map(D => \b3_PfG_6[5]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[5]\);
    
    \genblk9.b3_PfG_RNO[115]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[116]\, C => 
        \b7_vFW_PlM[114]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[115]\);
    
    \genblk9.b3_PfG_RNO[129]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[130]\, C => 
        \b7_vFW_PlM[128]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[129]\);
    
    \genblk9.b7_nYJ_BFM[128]\ : SLE
      port map(D => \b7_nYJ_BFM[127]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[128]\);
    
    \genblk9.b7_nYJ_BFM[55]\ : SLE
      port map(D => \b7_nYJ_BFM[54]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[55]\);
    
    \genblk9.b3_PfG_RNO[123]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[124]\, C => 
        \b7_vFW_PlM[122]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[123]\);
    
    \genblk9.b3_PfG_RNO[55]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[56]\, C => 
        \b7_vFW_PlM[54]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[55]\);
    
    \genblk9.un1_b7_nYJ_BFM8\ : CFG3
      generic map(INIT => x"EC")

      port map(A => b9_OFWNT9_ab, B => b11_nFG0rDY_9e2, C => 
        IICE_comm2iice(10), Y => un1_b7_nYJ_BFM8);
    
    \genblk9.b7_nYJ_BFM[98]\ : SLE
      port map(D => \b7_nYJ_BFM[97]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[98]\);
    
    \genblk9.b7_nYJ_BFM[35]\ : SLE
      port map(D => \b7_nYJ_BFM[34]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[35]\);
    
    \genblk9.b3_PfG[96]\ : SLE
      port map(D => \b3_PfG_6[96]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[96]\);
    
    \genblk9.b7_nYJ_BFM[44]\ : SLE
      port map(D => \b7_nYJ_BFM[43]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[44]\);
    
    \genblk9.b3_PfG[41]\ : SLE
      port map(D => \b3_PfG_6[41]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[41]\);
    
    \genblk9.b7_nYJ_BFM[22]\ : SLE
      port map(D => \b7_nYJ_BFM[21]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[22]\);
    
    \genblk9.b3_PfG_RNO[111]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[112]\, C => 
        \b7_vFW_PlM[110]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[111]\);
    
    \genblk9.b3_PfG[80]\ : SLE
      port map(D => \b3_PfG_6[80]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[80]\);
    
    \genblk9.b3_PfG_RNO[63]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[64]\, C => 
        \b7_vFW_PlM[62]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[63]\);
    
    \genblk9.b3_PfG[168]\ : SLE
      port map(D => \b3_PfG_6[168]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[168]\);
    
    \genblk9.b3_PfG[135]\ : SLE
      port map(D => \b3_PfG_6[135]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[135]\);
    
    \b8_FZFFLXYE[6]\ : SLE
      port map(D => \b12_2_St6KCa_jHv[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b4_2o_z, ALn => b5_voSc3_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b8_FZFFLXYE[6]_net_1\);
    
    \genblk9.b7_nYJ_BFM[132]\ : SLE
      port map(D => \b7_nYJ_BFM[131]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[132]\);
    
    \genblk9.b3_PfG_RNO[79]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[80]\, C => 
        \b7_vFW_PlM[78]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[79]\);
    
    \genblk9.b3_PfG_RNO[114]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[115]\, C => 
        \b7_vFW_PlM[113]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[114]\);
    
    \b12_PSyi_KyDbLbb[1]\ : SLE
      port map(D => \b12_2_St6KCa_jHv[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \b12_PSyi_KyDbLbb_0_sqmuxa\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \b12_PSyi_KyDbLbb[1]_net_1\);
    
    \genblk9.b3_PfG[113]\ : SLE
      port map(D => \b3_PfG_6[113]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[113]\);
    
    \genblk9.b3_PfG_RNO[43]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[44]\, C => 
        \b7_vFW_PlM[42]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[43]\);
    
    \genblk9.b7_nYJ_BFM[106]\ : SLE
      port map(D => \b7_nYJ_BFM[105]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[106]\);
    
    \genblk9.b7_nYJ_BFM[118]\ : SLE
      port map(D => \b7_nYJ_BFM[117]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[118]\);
    
    \genblk9.b7_nYJ_BFM[4]\ : SLE
      port map(D => \b7_nYJ_BFM[3]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[4]\);
    
    \genblk9.b3_PfG[12]\ : SLE
      port map(D => \b3_PfG_6[12]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[12]\);
    
    \genblk9.b3_PfG[37]\ : SLE
      port map(D => \b3_PfG_6[37]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[37]\);
    
    \genblk9.b3_PfG[58]\ : SLE
      port map(D => \b3_PfG_6[58]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[58]\);
    
    \genblk9.b7_nYJ_BFM[51]\ : SLE
      port map(D => \b7_nYJ_BFM[50]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[51]\);
    
    \genblk9.b3_PfG[110]\ : SLE
      port map(D => \b3_PfG_6[110]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[110]\);
    
    \genblk9.b3_PfG_RNO[119]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[120]\, C => 
        \b7_vFW_PlM[118]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[119]\);
    
    \genblk9.b3_PfG_RNO[74]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[75]\, C => 
        \b7_vFW_PlM[73]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[74]\);
    
    \genblk9.b3_PfG[19]\ : SLE
      port map(D => \b3_PfG_6[19]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[19]\);
    
    \genblk9.b3_PfG_RNO[113]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[114]\, C => 
        \b7_vFW_PlM[112]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[113]\);
    
    \genblk9.b3_PfG_RNO[32]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[33]\, C => 
        \b7_vFW_PlM[31]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[32]\);
    
    \b12_PSyi_KyDbLbb[4]\ : SLE
      port map(D => \b12_2_St6KCa_jHv[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \b12_PSyi_KyDbLbb_0_sqmuxa\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \b12_PSyi_KyDbLbb[4]_net_1\);
    
    \genblk9.b7_nYJ_BFM[31]\ : SLE
      port map(D => \b7_nYJ_BFM[30]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[31]\);
    
    \genblk9.b3_PfG_RNO[27]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[28]\, C => 
        \b7_vFW_PlM[26]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[27]\);
    
    \genblk9.b7_nYJ_BFM[3]\ : SLE
      port map(D => \b7_nYJ_BFM[2]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[3]\);
    
    \genblk9.b7_nYJ_BFM[10]\ : SLE
      port map(D => \b7_nYJ_BFM[9]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[10]\);
    
    \genblk9.b3_PfG_RNO[96]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[97]\, C => 
        \b7_vFW_PlM[95]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[96]\);
    
    \b12_2_St6KCa_jHv[3]\ : SLE
      port map(D => \b12_2_St6KCa_jHv_s[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b4_2o_z, ALn => b5_voSc3_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b12_2_St6KCa_jHv[3]_net_1\);
    
    \b12_PSyi_KyDbLbb[2]\ : SLE
      port map(D => \b12_2_St6KCa_jHv[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \b12_PSyi_KyDbLbb_0_sqmuxa\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \b12_PSyi_KyDbLbb[2]_net_1\);
    
    \genblk9.b7_nYJ_BFM[151]\ : SLE
      port map(D => \b7_nYJ_BFM[150]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[151]\);
    
    \genblk9.b7_nYJ_BFM[87]\ : SLE
      port map(D => \b7_nYJ_BFM[86]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[87]\);
    
    \genblk9.b3_PfG[46]\ : SLE
      port map(D => \b3_PfG_6[46]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[46]\);
    
    \genblk9.b3_PfG[133]\ : SLE
      port map(D => \b3_PfG_6[133]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[133]\);
    
    \genblk9.b3_PfG[155]\ : SLE
      port map(D => \b3_PfG_6[155]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[155]\);
    
    \genblk9.b3_PfG_RNO[130]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[131]\, C => 
        \b7_vFW_PlM[129]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[130]\);
    
    \genblk9.b3_PfG[32]\ : SLE
      port map(D => \b3_PfG_6[32]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[32]\);
    
    \b12_2_St6KCa_jHv[11]\ : SLE
      port map(D => \b12_2_St6KCa_jHv_s[11]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b4_2o_z, ALn => b5_voSc3_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b12_2_St6KCa_jHv[11]_net_1\);
    
    \genblk9.b7_nYJ_BFM[138]\ : SLE
      port map(D => \b7_nYJ_BFM[137]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[138]\);
    
    \genblk9.b3_PfG[75]\ : SLE
      port map(D => \b3_PfG_6[75]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[75]\);
    
    \genblk9.b3_PfG_RNO[59]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[60]\, C => 
        \b7_vFW_PlM[58]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[59]\);
    
    \genblk9.b3_PfG_RNO[67]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[68]\, C => 
        \b7_vFW_PlM[66]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[67]\);
    
    \genblk9.b7_nYJ_BFM[6]\ : SLE
      port map(D => \b7_nYJ_BFM[5]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[6]\);
    
    \genblk9.b7_nYJ_BFM[29]\ : SLE
      port map(D => \b7_nYJ_BFM[28]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[29]\);
    
    \genblk9.b3_PfG_RNO[81]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[82]\, C => 
        \b7_vFW_PlM[80]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[81]\);
    
    \genblk9.b3_PfG[130]\ : SLE
      port map(D => \b3_PfG_6[130]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[130]\);
    
    \genblk9.b3_PfG_RNO[80]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[81]\, C => 
        \b7_vFW_PlM[79]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[80]\);
    
    \genblk9.b9_v_mzCDYXs[5]\ : SLE
      port map(D => \b9_v_mzCDYXs_s[5]\, CLK => 
        IICE_comm2iice(11), EN => b9_v_mzCDYXs13, ALn => 
        b5_voSc3_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \b9_v_mzCDYXs[5]\);
    
    \genblk9.b3_PfG_RNO[47]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[48]\, C => 
        \b7_vFW_PlM[46]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[47]\);
    
    \genblk9.b3_PfG_RNO[100]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[101]\, C => 
        \b7_vFW_PlM[99]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[100]\);
    
    samplerStatus : b19_nczQ_DYg_YFaRM_oUoP_28s_1s_x_0
      port map(b8_FZFFLXYE(11) => \b8_FZFFLXYE[11]_net_1\, 
        b8_FZFFLXYE(10) => \b8_FZFFLXYE[10]_net_1\, 
        b8_FZFFLXYE(9) => \b8_FZFFLXYE[9]_net_1\, b8_FZFFLXYE(8)
         => \b8_FZFFLXYE[8]_net_1\, b8_FZFFLXYE(7) => 
        \b8_FZFFLXYE[7]_net_1\, b8_FZFFLXYE(6) => 
        \b8_FZFFLXYE[6]_net_1\, b8_FZFFLXYE(5) => 
        \b8_FZFFLXYE[5]_net_1\, b8_FZFFLXYE(4) => 
        \b8_FZFFLXYE[4]_net_1\, b8_FZFFLXYE(3) => 
        \b8_FZFFLXYE[3]_net_1\, b8_FZFFLXYE(2) => 
        \b8_FZFFLXYE[2]_net_1\, b8_FZFFLXYE(1) => 
        \b8_FZFFLXYE[1]_net_1\, b8_FZFFLXYE(0) => 
        \b8_FZFFLXYE[0]_net_1\, b12_PSyi_KyDbLbb(11) => 
        \b12_PSyi_KyDbLbb[11]_net_1\, b12_PSyi_KyDbLbb(10) => 
        \b12_PSyi_KyDbLbb[10]_net_1\, b12_PSyi_KyDbLbb(9) => 
        \b12_PSyi_KyDbLbb[9]_net_1\, b12_PSyi_KyDbLbb(8) => 
        \b12_PSyi_KyDbLbb[8]_net_1\, b12_PSyi_KyDbLbb(7) => 
        \b12_PSyi_KyDbLbb[7]_net_1\, b12_PSyi_KyDbLbb(6) => 
        \b12_PSyi_KyDbLbb[6]_net_1\, b12_PSyi_KyDbLbb(5) => 
        \b12_PSyi_KyDbLbb[5]_net_1\, b12_PSyi_KyDbLbb(4) => 
        \b12_PSyi_KyDbLbb[4]_net_1\, b12_PSyi_KyDbLbb(3) => 
        \b12_PSyi_KyDbLbb[3]_net_1\, b12_PSyi_KyDbLbb(2) => 
        \b12_PSyi_KyDbLbb[2]_net_1\, b12_PSyi_KyDbLbb(1) => 
        \b12_PSyi_KyDbLbb[1]_net_1\, b12_PSyi_KyDbLbb(0) => 
        \b12_PSyi_KyDbLbb[0]_net_1\, IICE_comm2iice_5 => 
        IICE_comm2iice(11), IICE_comm2iice_3 => IICE_comm2iice(9), 
        IICE_comm2iice_0 => IICE_comm2iice(6), IICE_comm2iice_4
         => IICE_comm2iice(10), b7_yYh03wy5 => b7_yYh03wy5, 
        b8_jAA_KlCO => \b8_jAA_KlCO\, ttdo => ttdo);
    
    \genblk9.b3_PfG_RNO[3]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[4]\, C => 
        \b7_vFW_PlM[2]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[3]\);
    
    \genblk9.b3_PfG[39]\ : SLE
      port map(D => \b3_PfG_6[39]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[39]\);
    
    \genblk9.b7_nYJ_BFM[46]\ : SLE
      port map(D => \b7_nYJ_BFM[45]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[46]\);
    
    \genblk9.b3_PfG[65]\ : SLE
      port map(D => \b3_PfG_6[65]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[65]\);
    
    \genblk9.b7_nYJ_BFM[160]\ : SLE
      port map(D => \b7_nYJ_BFM[159]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[160]\);
    
    \genblk9.b7_nYJ_BFM[140]\ : SLE
      port map(D => \b7_nYJ_BFM[139]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[140]\);
    
    \genblk9.b3_PfG[13]\ : SLE
      port map(D => \b3_PfG_6[13]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[13]\);
    
    \genblk9.b3_PfG_RNO[54]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[55]\, C => 
        \b7_vFW_PlM[53]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[54]\);
    
    \b12_2_St6KCa_jHv[9]\ : SLE
      port map(D => \b12_2_St6KCa_jHv_s[9]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b4_2o_z, ALn => b5_voSc3_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b12_2_St6KCa_jHv[9]_net_1\);
    
    \genblk9.b7_nYJ_BFM[156]\ : SLE
      port map(D => \b7_nYJ_BFM[155]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[156]\);
    
    \genblk9.b3_PfG[57]\ : SLE
      port map(D => \b3_PfG_6[57]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[57]\);
    
    \genblk9.b3_PfG[98]\ : SLE
      port map(D => \b3_PfG_6[98]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[98]\);
    
    \genblk9.b3_PfG_RNO[33]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[34]\, C => 
        \b7_vFW_PlM[32]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[33]\);
    
    b12_2_St6KCa_jHv_s_900 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \b12_2_St6KCa_jHv[0]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => 
        OPEN, Y => OPEN, FCO => b12_2_St6KCa_jHv_s_900_FCO);
    
    \genblk9.b3_PfG[149]\ : SLE
      port map(D => \b3_PfG_6[149]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[149]\);
    
    \genblk9.b3_PfG[24]\ : SLE
      port map(D => \b3_PfG_6[24]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[24]\);
    
    \genblk9.b7_nYJ_BFM[28]\ : SLE
      port map(D => \b7_nYJ_BFM[27]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[28]\);
    
    \genblk9.b7_nYJ_BFM[70]\ : SLE
      port map(D => \b7_nYJ_BFM[69]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[70]\);
    
    \genblk9.b3_PfG_RNO[16]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[17]\, C => 
        \b7_vFW_PlM[15]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[16]\);
    
    \genblk9.b3_PfG[153]\ : SLE
      port map(D => \b3_PfG_6[153]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[153]\);
    
    \genblk9.b11_nFG0rDY_9e2_2_0_a2\ : CFG3
      generic map(INIT => x"80")

      port map(A => IICE_comm2iice(6), B => b7_yYh03wy5, C => 
        IICE_comm2iice(10), Y => b11_nFG0rDY_9e2_2);
    
    \genblk9.b3_PfG_RNO[95]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[96]\, C => 
        \b7_vFW_PlM[94]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[95]\);
    
    \genblk9.b3_PfG_RNO[162]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[163]\, C => 
        \b7_vFW_PlM[161]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[162]\);
    
    \genblk9.b7_nYJ_BFM[60]\ : SLE
      port map(D => \b7_nYJ_BFM[59]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[60]\);
    
    \genblk9.b3_PfG[150]\ : SLE
      port map(D => \b3_PfG_6[150]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[150]\);
    
    \b12_2_St6KCa_jHv[8]\ : SLE
      port map(D => \b12_2_St6KCa_jHv_s[8]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b4_2o_z, ALn => b5_voSc3_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b12_2_St6KCa_jHv[8]_net_1\);
    
    \genblk9.b3_PfG[52]\ : SLE
      port map(D => \b3_PfG_6[52]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[52]\);
    
    \genblk9.b7_nYJ_BFM[13]\ : SLE
      port map(D => \b7_nYJ_BFM[12]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[13]\);
    
    \genblk9.b3_PfG[33]\ : SLE
      port map(D => \b3_PfG_6[33]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[33]\);
    
    \genblk9.b3_PfG[114]\ : SLE
      port map(D => \b3_PfG_6[114]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[114]\);
    
    \genblk9.b9_v_mzCDYXs[9]\ : SLE
      port map(D => \b9_v_mzCDYXs_s[9]\, CLK => 
        IICE_comm2iice(11), EN => b9_v_mzCDYXs13, ALn => 
        b5_voSc3_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \b9_v_mzCDYXs[9]\);
    
    \genblk9.b3_PfG[21]\ : SLE
      port map(D => \b3_PfG_6[21]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[21]\);
    
    \genblk9.b3_PfG_RNO[2]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[3]\, C => 
        \b7_vFW_PlM[1]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[2]\);
    
    \genblk9.b3_PfG_RNO[71]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[72]\, C => 
        \b7_vFW_PlM[70]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[71]\);
    
    \genblk9.b3_PfG_RNO[70]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[71]\, C => 
        \b7_vFW_PlM[69]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[70]\);
    
    \b12_PSyi_KyDbLbb[0]\ : SLE
      port map(D => \b12_2_St6KCa_jHv[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \b12_PSyi_KyDbLbb_0_sqmuxa\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \b12_PSyi_KyDbLbb[0]_net_1\);
    
    \genblk9.b3_PfG_RNO[168]\ : CFG3
      generic map(INIT => x"C8")

      port map(A => \b7_nYJ_BFM[174]\, B => \b7_vFW_PlM[167]\, C
         => b11_nFG0rDY_9e2, Y => \b3_PfG_6[168]\);
    
    \genblk9.b3_PfG_RNO[8]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[9]\, C => 
        \b7_vFW_PlM[7]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[8]\);
    
    \genblk9.b7_nYJ_BFM[90]\ : SLE
      port map(D => \b7_nYJ_BFM[89]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[90]\);
    
    \genblk9.b7_nYJ_BFM[52]\ : SLE
      port map(D => \b7_nYJ_BFM[51]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[52]\);
    
    \genblk9.b3_PfG_RNO[167]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[168]\, C => 
        \b7_vFW_PlM[166]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[167]\);
    
    \genblk9.b3_PfG[59]\ : SLE
      port map(D => \b3_PfG_6[59]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[59]\);
    
    \genblk9.b7_nYJ_BFM[32]\ : SLE
      port map(D => \b7_nYJ_BFM[31]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[32]\);
    
    \genblk9.b3_PfG[84]\ : SLE
      port map(D => \b3_PfG_6[84]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[84]\);
    
    \genblk9.b3_PfG_RNO[37]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[38]\, C => 
        \b7_vFW_PlM[36]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[37]\);
    
    \genblk9.b3_PfG[48]\ : SLE
      port map(D => \b3_PfG_6[48]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[48]\);
    
    \genblk9.b3_PfG[97]\ : SLE
      port map(D => \b3_PfG_6[97]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[97]\);
    
    \genblk9.b3_PfG_RNO[88]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[89]\, C => 
        \b7_vFW_PlM[87]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[88]\);
    
    \genblk9.b3_PfG[147]\ : SLE
      port map(D => \b3_PfG_6[147]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[147]\);
    
    \genblk9.b7_nYJ_BFM[14]\ : SLE
      port map(D => \b7_nYJ_BFM[13]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[14]\);
    
    \genblk9.b3_PfG_RNO[142]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[143]\, C => 
        \b7_vFW_PlM[141]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[142]\);
    
    \genblk9.b7_nYJ_BFM[169]\ : SLE
      port map(D => \b7_nYJ_BFM[168]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[169]\);
    
    \genblk9.b7_nYJ_BFM[149]\ : SLE
      port map(D => \b7_nYJ_BFM[148]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[149]\);
    
    \genblk9.b7_nYJ_BFM[7]\ : SLE
      port map(D => \b7_nYJ_BFM[6]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[7]\);
    
    \genblk9.b7_nYJ_BFM[47]\ : SLE
      port map(D => \b7_nYJ_BFM[46]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[47]\);
    
    \genblk9.b3_PfG[118]\ : SLE
      port map(D => \b3_PfG_6[118]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[118]\);
    
    \genblk9.b7_nYJ_BFM[85]\ : SLE
      port map(D => \b7_nYJ_BFM[84]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[85]\);
    
    \genblk9.b7_nYJ_BFM[0]\ : SLE
      port map(D => \b7_nYJ_BFM[174]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[0]\);
    
    \genblk9.b3_PfG[134]\ : SLE
      port map(D => \b3_PfG_6[134]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[134]\);
    
    \genblk9.b3_PfG_RNO[15]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[16]\, C => 
        \b7_vFW_PlM[14]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[15]\);
    
    \genblk9.b9_v_mzCDYXs[10]\ : SLE
      port map(D => \b9_v_mzCDYXs_s[10]\, CLK => 
        IICE_comm2iice(11), EN => b9_v_mzCDYXs13, ALn => 
        b5_voSc3_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \b9_v_mzCDYXs[10]\);
    
    \genblk9.b3_PfG[125]\ : SLE
      port map(D => \b3_PfG_6[125]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[125]\);
    
    b12_PSyi_KyDbLbb_0_sqmuxa : CFG4
      generic map(INIT => x"0008")

      port map(A => b13_wRBtT_ME83hHx, B => b4_2o_z, C => 
        \b9_PSyil9s_2\, D => b5_voSc3, Y => 
        \b12_PSyi_KyDbLbb_0_sqmuxa\);
    
    \genblk9.b3_PfG_RNO[122]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[123]\, C => 
        \b7_vFW_PlM[121]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[122]\);
    
    \genblk9.b3_PfG[81]\ : SLE
      port map(D => \b3_PfG_6[81]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[81]\);
    
    b8_jAA_KlCO_0_sqmuxa_1 : CFG4
      generic map(INIT => x"7FFF")

      port map(A => \b12_2_St6KCa_jHv[3]_net_1\, B => 
        \b12_2_St6KCa_jHv[2]_net_1\, C => 
        \b12_2_St6KCa_jHv[0]_net_1\, D => b4_2o_z, Y => 
        \b8_jAA_KlCO_0_sqmuxa_1\);
    
    \genblk9.b3_PfG_RNO[148]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[149]\, C => 
        \b7_vFW_PlM[147]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[148]\);
    
    \genblk9.b3_PfG_RNO[51]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[52]\, C => 
        \b7_vFW_PlM[50]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[51]\);
    
    \genblk9.b7_nYJ_BFM[165]\ : SLE
      port map(D => \b7_nYJ_BFM[164]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[165]\);
    
    \genblk9.b7_nYJ_BFM[145]\ : SLE
      port map(D => \b7_nYJ_BFM[144]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[145]\);
    
    \genblk9.b3_PfG_RNO[99]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[100]\, C => 
        \b7_vFW_PlM[98]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[99]\);
    
    \genblk9.b3_PfG[26]\ : SLE
      port map(D => \b3_PfG_6[26]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[26]\);
    
    \genblk9.b3_PfG_RNO[50]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[51]\, C => 
        \b7_vFW_PlM[49]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[50]\);
    
    \genblk9.b3_PfG_RNO[136]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[137]\, C => 
        \b7_vFW_PlM[135]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[136]\);
    
    \genblk9.b3_PfG_RNO[147]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[148]\, C => 
        \b7_vFW_PlM[146]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[147]\);
    
    \genblk9.b3_PfG[105]\ : SLE
      port map(D => \b3_PfG_6[105]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[105]\);
    
    \genblk9.b7_nYJ_BFM[73]\ : SLE
      port map(D => \b7_nYJ_BFM[72]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[73]\);
    
    \b12_2_St6KCa_jHv_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \b12_2_St6KCa_jHv[9]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \b12_2_St6KCa_jHv_cry[8]_net_1\, S => 
        \b12_2_St6KCa_jHv_s[9]\, Y => OPEN, FCO => 
        \b12_2_St6KCa_jHv_cry[9]_net_1\);
    
    \genblk9.b7_nYJ_BFM[163]\ : SLE
      port map(D => \b7_nYJ_BFM[162]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[163]\);
    
    \genblk9.b7_nYJ_BFM[143]\ : SLE
      port map(D => \b7_nYJ_BFM[142]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[143]\);
    
    \genblk9.b3_PfG_RNO[155]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[156]\, C => 
        \b7_vFW_PlM[154]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[155]\);
    
    \genblk9.b7_nYJ_BFM[5]\ : SLE
      port map(D => \b7_nYJ_BFM[4]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[5]\);
    
    \genblk9.b9_v_mzCDYXs_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \b9_v_mzCDYXs[0]\, Y => \b9_v_mzCDYXs_s[0]\);
    
    \genblk9.b3_PfG[53]\ : SLE
      port map(D => \b3_PfG_6[53]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[53]\);
    
    \genblk9.b3_PfG[92]\ : SLE
      port map(D => \b3_PfG_6[92]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[92]\);
    
    \genblk9.b3_PfG[167]\ : SLE
      port map(D => \b3_PfG_6[167]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[167]\);
    
    \genblk9.b7_nYJ_BFM[63]\ : SLE
      port map(D => \b7_nYJ_BFM[62]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[63]\);
    
    \genblk9.b3_PfG_RNO[106]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[107]\, C => 
        \b7_vFW_PlM[105]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[106]\);
    
    \genblk9.b3_PfG_RNO[128]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[129]\, C => 
        \b7_vFW_PlM[127]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[128]\);
    
    \genblk9.b3_PfG[138]\ : SLE
      port map(D => \b3_PfG_6[138]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[138]\);
    
    \genblk9.b7_nYJ_BFM[81]\ : SLE
      port map(D => \b7_nYJ_BFM[80]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[81]\);
    
    \genblk9.b3_PfG_RNO[94]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[95]\, C => 
        \b7_vFW_PlM[93]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[94]\);
    
    \genblk9.b7_nYJ_BFM[164]\ : SLE
      port map(D => \b7_nYJ_BFM[163]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[164]\);
    
    \genblk9.b7_nYJ_BFM[2]\ : SLE
      port map(D => \b7_nYJ_BFM[1]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[2]\);
    
    \genblk9.b7_nYJ_BFM[144]\ : SLE
      port map(D => \b7_nYJ_BFM[143]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[144]\);
    
    \genblk9.b3_PfG_RNO[127]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[128]\, C => 
        \b7_vFW_PlM[126]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[127]\);
    
    \genblk9.b3_PfG[99]\ : SLE
      port map(D => \b3_PfG_6[99]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[99]\);
    
    \genblk9.b3_PfG_RNO[151]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[152]\, C => 
        \b7_vFW_PlM[150]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[151]\);
    
    \genblk9.b7_nYJ_BFM[59]\ : SLE
      port map(D => \b7_nYJ_BFM[58]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[59]\);
    
    \genblk9.b9_v_mzCDYXs_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \b9_v_mzCDYXs[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => \b9_v_mzCDYXs_cry[9]\, 
        S => \b9_v_mzCDYXs_s[10]\, Y => OPEN, FCO => 
        \b9_v_mzCDYXs_cry[10]\);
    
    \genblk9.b3_PfG[47]\ : SLE
      port map(D => \b3_PfG_6[47]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[47]\);
    
    \genblk9.b3_PfG[154]\ : SLE
      port map(D => \b3_PfG_6[154]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[154]\);
    
    \genblk9.b7_nYJ_BFM[39]\ : SLE
      port map(D => \b7_nYJ_BFM[38]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[39]\);
    
    \genblk9.b3_PfG_RNO[78]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[79]\, C => 
        \b7_vFW_PlM[77]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[78]\);
    
    \genblk9.b3_PfG[142]\ : SLE
      port map(D => \b3_PfG_6[142]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[142]\);
    
    \genblk9.b3_PfG[70]\ : SLE
      port map(D => \b3_PfG_6[70]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[70]\);
    
    \genblk9.b7_nYJ_BFM[74]\ : SLE
      port map(D => \b7_nYJ_BFM[73]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[74]\);
    
    \genblk9.b3_PfG_RNO[154]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[155]\, C => 
        \b7_vFW_PlM[153]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[154]\);
    
    \genblk9.b3_PfG[123]\ : SLE
      port map(D => \b3_PfG_6[123]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[123]\);
    
    \genblk9.b3_PfG[15]\ : SLE
      port map(D => \b3_PfG_6[15]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[15]\);
    
    \genblk9.b3_PfG_RNO[26]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[27]\, C => 
        \b7_vFW_PlM[25]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[26]\);
    
    \genblk9.b3_PfG_RNO[112]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[113]\, C => 
        \b7_vFW_PlM[111]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[112]\);
    
    \genblk9.b7_nYJ_BFM[93]\ : SLE
      port map(D => \b7_nYJ_BFM[92]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[93]\);
    
    \genblk9.b7_nYJ_BFM[127]\ : SLE
      port map(D => \b7_nYJ_BFM[126]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[127]\);
    
    \b12_PSyi_KyDbLbb[3]\ : SLE
      port map(D => \b12_2_St6KCa_jHv[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \b12_PSyi_KyDbLbb_0_sqmuxa\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \b12_PSyi_KyDbLbb[3]_net_1\);
    
    \genblk9.b7_nYJ_BFM[64]\ : SLE
      port map(D => \b7_nYJ_BFM[63]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[64]\);
    
    \genblk9.b3_PfG[103]\ : SLE
      port map(D => \b3_PfG_6[103]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[103]\);
    
    b8_jAA_KlCO_0_sqmuxa : CFG4
      generic map(INIT => x"0080")

      port map(A => \b12_2_St6KCa_jHv[1]_net_1\, B => 
        \b8_jAA_KlCO_0_sqmuxa_8\, C => \b8_jAA_KlCO_0_sqmuxa_7\, 
        D => \b8_jAA_KlCO_0_sqmuxa_1\, Y => 
        \b8_jAA_KlCO_0_sqmuxa\);
    
    \genblk9.b3_PfG[60]\ : SLE
      port map(D => \b3_PfG_6[60]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[60]\);
    
    \genblk9.b3_PfG[120]\ : SLE
      port map(D => \b3_PfG_6[120]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[120]\);
    
    \genblk9.b3_PfG_RNO[159]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[160]\, C => 
        \b7_vFW_PlM[158]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[159]\);
    
    \genblk9.b7_nYJ_BFM[16]\ : SLE
      port map(D => \b7_nYJ_BFM[15]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[16]\);
    
    \genblk9.b7_nYJ_BFM[58]\ : SLE
      port map(D => \b7_nYJ_BFM[57]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[58]\);
    
    \genblk9.b3_PfG_RNO[153]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[154]\, C => 
        \b7_vFW_PlM[152]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[153]\);
    
    \genblk9.b3_PfG[86]\ : SLE
      port map(D => \b3_PfG_6[86]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[86]\);
    
    \genblk9.b7_nYJ_BFM[162]\ : SLE
      port map(D => \b7_nYJ_BFM[161]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[162]\);
    
    \genblk9.b9_v_mzCDYXs[8]\ : SLE
      port map(D => \b9_v_mzCDYXs_s[8]\, CLK => 
        IICE_comm2iice(11), EN => b9_v_mzCDYXs13, ALn => 
        b5_voSc3_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \b9_v_mzCDYXs[8]\);
    
    \genblk9.b3_PfG_RNO[160]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[161]\, C => 
        \b7_vFW_PlM[159]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[160]\);
    
    \genblk9.b7_nYJ_BFM[142]\ : SLE
      port map(D => \b7_nYJ_BFM[141]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[142]\);
    
    \genblk9.b7_nYJ_BFM[20]\ : SLE
      port map(D => \b7_nYJ_BFM[19]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[20]\);
    
    \genblk9.b3_PfG_RNO[19]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[20]\, C => 
        \b7_vFW_PlM[18]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[19]\);
    
    \genblk9.b3_PfG[4]\ : SLE
      port map(D => \b3_PfG_6[4]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[4]\);
    
    \genblk9.b7_nYJ_BFM[38]\ : SLE
      port map(D => \b7_nYJ_BFM[37]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[38]\);
    
    \genblk9.b7_nYJ_BFM[100]\ : SLE
      port map(D => \b7_nYJ_BFM[99]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[100]\);
    
    \genblk9.b3_PfG[100]\ : SLE
      port map(D => \b3_PfG_6[100]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[100]\);
    
    \genblk9.b3_PfG_RNO[118]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[119]\, C => 
        \b7_vFW_PlM[117]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[118]\);
    
    \genblk9.b3_PfG[158]\ : SLE
      port map(D => \b3_PfG_6[158]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[158]\);
    
    \genblk9.b9_v_mzCDYXs_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \b9_v_mzCDYXs[9]\, C => 
        GND_net_1, D => GND_net_1, FCI => \b9_v_mzCDYXs_cry[8]\, 
        S => \b9_v_mzCDYXs_s[9]\, Y => OPEN, FCO => 
        \b9_v_mzCDYXs_cry[9]\);
    
    \genblk9.b9_v_mzCDYXs13_0_a2\ : CFG3
      generic map(INIT => x"80")

      port map(A => b9_OFWNT9_ab, B => \b7_nYJ_BFM[0]\, C => 
        IICE_comm2iice(10), Y => b9_v_mzCDYXs13);
    
    \genblk9.b3_PfG_RNO[117]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[118]\, C => 
        \b7_vFW_PlM[116]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[117]\);
    
    \genblk9.b3_PfG_RNO[66]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[67]\, C => 
        \b7_vFW_PlM[65]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[66]\);
    
    \genblk9.b3_PfG[42]\ : SLE
      port map(D => \b3_PfG_6[42]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[42]\);
    
    \genblk9.b7_nYJ_BFM[94]\ : SLE
      port map(D => \b7_nYJ_BFM[93]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[94]\);
    
    \genblk9.b3_PfG[162]\ : SLE
      port map(D => \b3_PfG_6[162]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[162]\);
    
    \b12_2_St6KCa_jHv_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \b12_2_St6KCa_jHv[6]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \b12_2_St6KCa_jHv_cry[5]_net_1\, S => 
        \b12_2_St6KCa_jHv_s[6]\, Y => OPEN, FCO => 
        \b12_2_St6KCa_jHv_cry[6]_net_1\);
    
    \genblk9.b7_nYJ_BFM[117]\ : SLE
      port map(D => \b7_nYJ_BFM[116]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[117]\);
    
    b8_jAA_KlCO : SLE
      port map(D => VCC_net_1, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \b8_jAA_KlCO_0_sqmuxa\, ALn => b5_voSc3_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b8_jAA_KlCO\);
    
    \genblk9.b3_PfG_RNO[46]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[47]\, C => 
        \b7_vFW_PlM[45]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[46]\);
    
    \genblk9.b3_PfG[93]\ : SLE
      port map(D => \b3_PfG_6[93]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[93]\);
    
    \genblk9.b3_PfG[35]\ : SLE
      port map(D => \b3_PfG_6[35]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[35]\);
    
    \genblk9.b3_PfG_RNO[14]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[15]\, C => 
        \b7_vFW_PlM[13]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[14]\);
    
    b3_SoW : b13_vFW_xNywD_EdR_174s_12s_4096s_0s_x_0
      port map(b11_OFWNT9L_8tZ(167) => \b11_OFWNT9L_8tZ[167]\, 
        b11_OFWNT9L_8tZ(166) => \b11_OFWNT9L_8tZ[166]\, 
        b11_OFWNT9L_8tZ(165) => \b11_OFWNT9L_8tZ[165]\, 
        b11_OFWNT9L_8tZ(164) => \b11_OFWNT9L_8tZ[164]\, 
        b11_OFWNT9L_8tZ(163) => \b11_OFWNT9L_8tZ[163]\, 
        b11_OFWNT9L_8tZ(162) => \b11_OFWNT9L_8tZ[162]\, 
        b11_OFWNT9L_8tZ(161) => \b11_OFWNT9L_8tZ[161]\, 
        b11_OFWNT9L_8tZ(160) => \b11_OFWNT9L_8tZ[160]\, 
        b11_OFWNT9L_8tZ(159) => \b11_OFWNT9L_8tZ[159]\, 
        b11_OFWNT9L_8tZ(158) => \b11_OFWNT9L_8tZ[158]\, 
        b11_OFWNT9L_8tZ(157) => \b11_OFWNT9L_8tZ[157]\, 
        b11_OFWNT9L_8tZ(156) => \b11_OFWNT9L_8tZ[156]\, 
        b11_OFWNT9L_8tZ(155) => \b11_OFWNT9L_8tZ[155]\, 
        b11_OFWNT9L_8tZ(154) => \b11_OFWNT9L_8tZ[154]\, 
        b11_OFWNT9L_8tZ(153) => \b11_OFWNT9L_8tZ[153]\, 
        b11_OFWNT9L_8tZ(152) => \b11_OFWNT9L_8tZ[152]\, 
        b11_OFWNT9L_8tZ(151) => \b11_OFWNT9L_8tZ[151]\, 
        b11_OFWNT9L_8tZ(150) => \b11_OFWNT9L_8tZ[150]\, 
        b11_OFWNT9L_8tZ(149) => \b11_OFWNT9L_8tZ[149]\, 
        b11_OFWNT9L_8tZ(148) => \b11_OFWNT9L_8tZ[148]\, 
        b11_OFWNT9L_8tZ(147) => \b11_OFWNT9L_8tZ[147]\, 
        b11_OFWNT9L_8tZ(146) => \b11_OFWNT9L_8tZ[146]\, 
        b11_OFWNT9L_8tZ(145) => \b11_OFWNT9L_8tZ[145]\, 
        b11_OFWNT9L_8tZ(144) => \b11_OFWNT9L_8tZ[144]\, 
        b11_OFWNT9L_8tZ(143) => \b11_OFWNT9L_8tZ[143]\, 
        b11_OFWNT9L_8tZ(142) => \b11_OFWNT9L_8tZ[142]\, 
        b11_OFWNT9L_8tZ(141) => \b11_OFWNT9L_8tZ[141]\, 
        b11_OFWNT9L_8tZ(140) => \b11_OFWNT9L_8tZ[140]\, 
        b11_OFWNT9L_8tZ(139) => \b11_OFWNT9L_8tZ[139]\, 
        b11_OFWNT9L_8tZ(138) => \b11_OFWNT9L_8tZ[138]\, 
        b11_OFWNT9L_8tZ(137) => \b11_OFWNT9L_8tZ[137]\, 
        b11_OFWNT9L_8tZ(136) => \b11_OFWNT9L_8tZ[136]\, 
        b11_OFWNT9L_8tZ(135) => \b11_OFWNT9L_8tZ[135]\, 
        b11_OFWNT9L_8tZ(134) => \b11_OFWNT9L_8tZ[134]\, 
        b11_OFWNT9L_8tZ(133) => \b11_OFWNT9L_8tZ[133]\, 
        b11_OFWNT9L_8tZ(132) => \b11_OFWNT9L_8tZ[132]\, 
        b11_OFWNT9L_8tZ(131) => \b11_OFWNT9L_8tZ[131]\, 
        b11_OFWNT9L_8tZ(130) => \b11_OFWNT9L_8tZ[130]\, 
        b11_OFWNT9L_8tZ(129) => \b11_OFWNT9L_8tZ[129]\, 
        b11_OFWNT9L_8tZ(128) => \b11_OFWNT9L_8tZ[128]\, 
        b11_OFWNT9L_8tZ(127) => \b11_OFWNT9L_8tZ[127]\, 
        b11_OFWNT9L_8tZ(126) => \b11_OFWNT9L_8tZ[126]\, 
        b11_OFWNT9L_8tZ(125) => \b11_OFWNT9L_8tZ[125]\, 
        b11_OFWNT9L_8tZ(124) => \b11_OFWNT9L_8tZ[124]\, 
        b11_OFWNT9L_8tZ(123) => \b11_OFWNT9L_8tZ[123]\, 
        b11_OFWNT9L_8tZ(122) => \b11_OFWNT9L_8tZ[122]\, 
        b11_OFWNT9L_8tZ(121) => \b11_OFWNT9L_8tZ[121]\, 
        b11_OFWNT9L_8tZ(120) => \b11_OFWNT9L_8tZ[120]\, 
        b11_OFWNT9L_8tZ(119) => \b11_OFWNT9L_8tZ[119]\, 
        b11_OFWNT9L_8tZ(118) => \b11_OFWNT9L_8tZ[118]\, 
        b11_OFWNT9L_8tZ(117) => \b11_OFWNT9L_8tZ[117]\, 
        b11_OFWNT9L_8tZ(116) => \b11_OFWNT9L_8tZ[116]\, 
        b11_OFWNT9L_8tZ(115) => \b11_OFWNT9L_8tZ[115]\, 
        b11_OFWNT9L_8tZ(114) => \b11_OFWNT9L_8tZ[114]\, 
        b11_OFWNT9L_8tZ(113) => \b11_OFWNT9L_8tZ[113]\, 
        b11_OFWNT9L_8tZ(112) => \b11_OFWNT9L_8tZ[112]\, 
        b11_OFWNT9L_8tZ(111) => \b11_OFWNT9L_8tZ[111]\, 
        b11_OFWNT9L_8tZ(110) => \b11_OFWNT9L_8tZ[110]\, 
        b11_OFWNT9L_8tZ(109) => \b11_OFWNT9L_8tZ[109]\, 
        b11_OFWNT9L_8tZ(108) => \b11_OFWNT9L_8tZ[108]\, 
        b11_OFWNT9L_8tZ(107) => \b11_OFWNT9L_8tZ[107]\, 
        b11_OFWNT9L_8tZ(106) => \b11_OFWNT9L_8tZ[106]\, 
        b11_OFWNT9L_8tZ(105) => \b11_OFWNT9L_8tZ[105]\, 
        b11_OFWNT9L_8tZ(104) => \b11_OFWNT9L_8tZ[104]\, 
        b11_OFWNT9L_8tZ(103) => \b11_OFWNT9L_8tZ[103]\, 
        b11_OFWNT9L_8tZ(102) => \b11_OFWNT9L_8tZ[102]\, 
        b11_OFWNT9L_8tZ(101) => \b11_OFWNT9L_8tZ[101]\, 
        b11_OFWNT9L_8tZ(100) => \b11_OFWNT9L_8tZ[100]\, 
        b11_OFWNT9L_8tZ(99) => \b11_OFWNT9L_8tZ[99]\, 
        b11_OFWNT9L_8tZ(98) => \b11_OFWNT9L_8tZ[98]\, 
        b11_OFWNT9L_8tZ(97) => \b11_OFWNT9L_8tZ[97]\, 
        b11_OFWNT9L_8tZ(96) => \b11_OFWNT9L_8tZ[96]\, 
        b11_OFWNT9L_8tZ(95) => \b11_OFWNT9L_8tZ[95]\, 
        b11_OFWNT9L_8tZ(94) => \b11_OFWNT9L_8tZ[94]\, 
        b11_OFWNT9L_8tZ(93) => \b11_OFWNT9L_8tZ[93]\, 
        b11_OFWNT9L_8tZ(92) => \b11_OFWNT9L_8tZ[92]\, 
        b11_OFWNT9L_8tZ(91) => \b11_OFWNT9L_8tZ[91]\, 
        b11_OFWNT9L_8tZ(90) => \b11_OFWNT9L_8tZ[90]\, 
        b11_OFWNT9L_8tZ(89) => \b11_OFWNT9L_8tZ[89]\, 
        b11_OFWNT9L_8tZ(88) => \b11_OFWNT9L_8tZ[88]\, 
        b11_OFWNT9L_8tZ(87) => \b11_OFWNT9L_8tZ[87]\, 
        b11_OFWNT9L_8tZ(86) => \b11_OFWNT9L_8tZ[86]\, 
        b11_OFWNT9L_8tZ(85) => \b11_OFWNT9L_8tZ[85]\, 
        b11_OFWNT9L_8tZ(84) => \b11_OFWNT9L_8tZ[84]\, 
        b11_OFWNT9L_8tZ(83) => \b11_OFWNT9L_8tZ[83]\, 
        b11_OFWNT9L_8tZ(82) => \b11_OFWNT9L_8tZ[82]\, 
        b11_OFWNT9L_8tZ(81) => \b11_OFWNT9L_8tZ[81]\, 
        b11_OFWNT9L_8tZ(80) => \b11_OFWNT9L_8tZ[80]\, 
        b11_OFWNT9L_8tZ(79) => \b11_OFWNT9L_8tZ[79]\, 
        b11_OFWNT9L_8tZ(78) => \b11_OFWNT9L_8tZ[78]\, 
        b11_OFWNT9L_8tZ(77) => \b11_OFWNT9L_8tZ[77]\, 
        b11_OFWNT9L_8tZ(76) => \b11_OFWNT9L_8tZ[76]\, 
        b11_OFWNT9L_8tZ(75) => \b11_OFWNT9L_8tZ[75]\, 
        b11_OFWNT9L_8tZ(74) => \b11_OFWNT9L_8tZ[74]\, 
        b11_OFWNT9L_8tZ(73) => \b11_OFWNT9L_8tZ[73]\, 
        b11_OFWNT9L_8tZ(72) => \b11_OFWNT9L_8tZ[72]\, 
        b11_OFWNT9L_8tZ(71) => \b11_OFWNT9L_8tZ[71]\, 
        b11_OFWNT9L_8tZ(70) => \b11_OFWNT9L_8tZ[70]\, 
        b11_OFWNT9L_8tZ(69) => \b11_OFWNT9L_8tZ[69]\, 
        b11_OFWNT9L_8tZ(68) => \b11_OFWNT9L_8tZ[68]\, 
        b11_OFWNT9L_8tZ(67) => \b11_OFWNT9L_8tZ[67]\, 
        b11_OFWNT9L_8tZ(66) => \b11_OFWNT9L_8tZ[66]\, 
        b11_OFWNT9L_8tZ(65) => \b11_OFWNT9L_8tZ[65]\, 
        b11_OFWNT9L_8tZ(64) => \b11_OFWNT9L_8tZ[64]\, 
        b11_OFWNT9L_8tZ(63) => \b11_OFWNT9L_8tZ[63]\, 
        b11_OFWNT9L_8tZ(62) => \b11_OFWNT9L_8tZ[62]\, 
        b11_OFWNT9L_8tZ(61) => \b11_OFWNT9L_8tZ[61]\, 
        b11_OFWNT9L_8tZ(60) => \b11_OFWNT9L_8tZ[60]\, 
        b11_OFWNT9L_8tZ(59) => \b11_OFWNT9L_8tZ[59]\, 
        b11_OFWNT9L_8tZ(58) => \b11_OFWNT9L_8tZ[58]\, 
        b11_OFWNT9L_8tZ(57) => \b11_OFWNT9L_8tZ[57]\, 
        b11_OFWNT9L_8tZ(56) => \b11_OFWNT9L_8tZ[56]\, 
        b11_OFWNT9L_8tZ(55) => \b11_OFWNT9L_8tZ[55]\, 
        b11_OFWNT9L_8tZ(54) => \b11_OFWNT9L_8tZ[54]\, 
        b11_OFWNT9L_8tZ(53) => \b11_OFWNT9L_8tZ[53]\, 
        b11_OFWNT9L_8tZ(52) => \b11_OFWNT9L_8tZ[52]\, 
        b11_OFWNT9L_8tZ(51) => \b11_OFWNT9L_8tZ[51]\, 
        b11_OFWNT9L_8tZ(50) => \b11_OFWNT9L_8tZ[50]\, 
        b11_OFWNT9L_8tZ(49) => \b11_OFWNT9L_8tZ[49]\, 
        b11_OFWNT9L_8tZ(48) => \b11_OFWNT9L_8tZ[48]\, 
        b11_OFWNT9L_8tZ(47) => \b11_OFWNT9L_8tZ[47]\, 
        b11_OFWNT9L_8tZ(46) => \b11_OFWNT9L_8tZ[46]\, 
        b11_OFWNT9L_8tZ(45) => \b11_OFWNT9L_8tZ[45]\, 
        b11_OFWNT9L_8tZ(44) => \b11_OFWNT9L_8tZ[44]\, 
        b11_OFWNT9L_8tZ(43) => \b11_OFWNT9L_8tZ[43]\, 
        b11_OFWNT9L_8tZ(42) => \b11_OFWNT9L_8tZ[42]\, 
        b11_OFWNT9L_8tZ(41) => \b11_OFWNT9L_8tZ[41]\, 
        b11_OFWNT9L_8tZ(40) => \b11_OFWNT9L_8tZ[40]\, 
        b11_OFWNT9L_8tZ(39) => \b11_OFWNT9L_8tZ[39]\, 
        b11_OFWNT9L_8tZ(38) => \b11_OFWNT9L_8tZ[38]\, 
        b11_OFWNT9L_8tZ(37) => \b11_OFWNT9L_8tZ[37]\, 
        b11_OFWNT9L_8tZ(36) => \b11_OFWNT9L_8tZ[36]\, 
        b11_OFWNT9L_8tZ(35) => \b11_OFWNT9L_8tZ[35]\, 
        b11_OFWNT9L_8tZ(34) => \b11_OFWNT9L_8tZ[34]\, 
        b11_OFWNT9L_8tZ(33) => \b11_OFWNT9L_8tZ[33]\, 
        b11_OFWNT9L_8tZ(32) => \b11_OFWNT9L_8tZ[32]\, 
        b11_OFWNT9L_8tZ(31) => \b11_OFWNT9L_8tZ[31]\, 
        b11_OFWNT9L_8tZ(30) => \b11_OFWNT9L_8tZ[30]\, 
        b11_OFWNT9L_8tZ(29) => \b11_OFWNT9L_8tZ[29]\, 
        b11_OFWNT9L_8tZ(28) => \b11_OFWNT9L_8tZ[28]\, 
        b11_OFWNT9L_8tZ(27) => \b11_OFWNT9L_8tZ[27]\, 
        b11_OFWNT9L_8tZ(26) => \b11_OFWNT9L_8tZ[26]\, 
        b11_OFWNT9L_8tZ(25) => \b11_OFWNT9L_8tZ[25]\, 
        b11_OFWNT9L_8tZ(24) => \b11_OFWNT9L_8tZ[24]\, 
        b11_OFWNT9L_8tZ(23) => \b11_OFWNT9L_8tZ[23]\, 
        b11_OFWNT9L_8tZ(22) => \b11_OFWNT9L_8tZ[22]\, 
        b11_OFWNT9L_8tZ(21) => \b11_OFWNT9L_8tZ[21]\, 
        b11_OFWNT9L_8tZ(20) => \b11_OFWNT9L_8tZ[20]\, 
        b11_OFWNT9L_8tZ(19) => \b11_OFWNT9L_8tZ[19]\, 
        b11_OFWNT9L_8tZ(18) => \b11_OFWNT9L_8tZ[18]\, 
        b11_OFWNT9L_8tZ(17) => \b11_OFWNT9L_8tZ[17]\, 
        b11_OFWNT9L_8tZ(16) => \b11_OFWNT9L_8tZ[16]\, 
        b11_OFWNT9L_8tZ(15) => \b11_OFWNT9L_8tZ[15]\, 
        b11_OFWNT9L_8tZ(14) => \b11_OFWNT9L_8tZ[14]\, 
        b11_OFWNT9L_8tZ(13) => \b11_OFWNT9L_8tZ[13]\, 
        b11_OFWNT9L_8tZ(12) => \b11_OFWNT9L_8tZ[12]\, 
        b11_OFWNT9L_8tZ(11) => \b11_OFWNT9L_8tZ[11]\, 
        b11_OFWNT9L_8tZ(10) => \b11_OFWNT9L_8tZ[10]\, 
        b11_OFWNT9L_8tZ(9) => \b11_OFWNT9L_8tZ[9]\, 
        b11_OFWNT9L_8tZ(8) => \b11_OFWNT9L_8tZ[8]\, 
        b11_OFWNT9L_8tZ(7) => \b11_OFWNT9L_8tZ[7]\, 
        b11_OFWNT9L_8tZ(6) => \b11_OFWNT9L_8tZ[6]\, 
        b11_OFWNT9L_8tZ(5) => \b11_OFWNT9L_8tZ[5]\, 
        b11_OFWNT9L_8tZ(4) => \b11_OFWNT9L_8tZ[4]\, 
        b11_OFWNT9L_8tZ(3) => \b11_OFWNT9L_8tZ[3]\, 
        b11_OFWNT9L_8tZ(2) => \b11_OFWNT9L_8tZ[2]\, 
        b11_OFWNT9L_8tZ(1) => \b11_OFWNT9L_8tZ[1]\, 
        b11_OFWNT9L_8tZ(0) => \b11_OFWNT9L_8tZ[0]\, 
        b7_vFW_PlM(167) => \b7_vFW_PlM[167]\, b7_vFW_PlM(166) => 
        \b7_vFW_PlM[166]\, b7_vFW_PlM(165) => \b7_vFW_PlM[165]\, 
        b7_vFW_PlM(164) => \b7_vFW_PlM[164]\, b7_vFW_PlM(163) => 
        \b7_vFW_PlM[163]\, b7_vFW_PlM(162) => \b7_vFW_PlM[162]\, 
        b7_vFW_PlM(161) => \b7_vFW_PlM[161]\, b7_vFW_PlM(160) => 
        \b7_vFW_PlM[160]\, b7_vFW_PlM(159) => \b7_vFW_PlM[159]\, 
        b7_vFW_PlM(158) => \b7_vFW_PlM[158]\, b7_vFW_PlM(157) => 
        \b7_vFW_PlM[157]\, b7_vFW_PlM(156) => \b7_vFW_PlM[156]\, 
        b7_vFW_PlM(155) => \b7_vFW_PlM[155]\, b7_vFW_PlM(154) => 
        \b7_vFW_PlM[154]\, b7_vFW_PlM(153) => \b7_vFW_PlM[153]\, 
        b7_vFW_PlM(152) => \b7_vFW_PlM[152]\, b7_vFW_PlM(151) => 
        \b7_vFW_PlM[151]\, b7_vFW_PlM(150) => \b7_vFW_PlM[150]\, 
        b7_vFW_PlM(149) => \b7_vFW_PlM[149]\, b7_vFW_PlM(148) => 
        \b7_vFW_PlM[148]\, b7_vFW_PlM(147) => \b7_vFW_PlM[147]\, 
        b7_vFW_PlM(146) => \b7_vFW_PlM[146]\, b7_vFW_PlM(145) => 
        \b7_vFW_PlM[145]\, b7_vFW_PlM(144) => \b7_vFW_PlM[144]\, 
        b7_vFW_PlM(143) => \b7_vFW_PlM[143]\, b7_vFW_PlM(142) => 
        \b7_vFW_PlM[142]\, b7_vFW_PlM(141) => \b7_vFW_PlM[141]\, 
        b7_vFW_PlM(140) => \b7_vFW_PlM[140]\, b7_vFW_PlM(139) => 
        \b7_vFW_PlM[139]\, b7_vFW_PlM(138) => \b7_vFW_PlM[138]\, 
        b7_vFW_PlM(137) => \b7_vFW_PlM[137]\, b7_vFW_PlM(136) => 
        \b7_vFW_PlM[136]\, b7_vFW_PlM(135) => \b7_vFW_PlM[135]\, 
        b7_vFW_PlM(134) => \b7_vFW_PlM[134]\, b7_vFW_PlM(133) => 
        \b7_vFW_PlM[133]\, b7_vFW_PlM(132) => \b7_vFW_PlM[132]\, 
        b7_vFW_PlM(131) => \b7_vFW_PlM[131]\, b7_vFW_PlM(130) => 
        \b7_vFW_PlM[130]\, b7_vFW_PlM(129) => \b7_vFW_PlM[129]\, 
        b7_vFW_PlM(128) => \b7_vFW_PlM[128]\, b7_vFW_PlM(127) => 
        \b7_vFW_PlM[127]\, b7_vFW_PlM(126) => \b7_vFW_PlM[126]\, 
        b7_vFW_PlM(125) => \b7_vFW_PlM[125]\, b7_vFW_PlM(124) => 
        \b7_vFW_PlM[124]\, b7_vFW_PlM(123) => \b7_vFW_PlM[123]\, 
        b7_vFW_PlM(122) => \b7_vFW_PlM[122]\, b7_vFW_PlM(121) => 
        \b7_vFW_PlM[121]\, b7_vFW_PlM(120) => \b7_vFW_PlM[120]\, 
        b7_vFW_PlM(119) => \b7_vFW_PlM[119]\, b7_vFW_PlM(118) => 
        \b7_vFW_PlM[118]\, b7_vFW_PlM(117) => \b7_vFW_PlM[117]\, 
        b7_vFW_PlM(116) => \b7_vFW_PlM[116]\, b7_vFW_PlM(115) => 
        \b7_vFW_PlM[115]\, b7_vFW_PlM(114) => \b7_vFW_PlM[114]\, 
        b7_vFW_PlM(113) => \b7_vFW_PlM[113]\, b7_vFW_PlM(112) => 
        \b7_vFW_PlM[112]\, b7_vFW_PlM(111) => \b7_vFW_PlM[111]\, 
        b7_vFW_PlM(110) => \b7_vFW_PlM[110]\, b7_vFW_PlM(109) => 
        \b7_vFW_PlM[109]\, b7_vFW_PlM(108) => \b7_vFW_PlM[108]\, 
        b7_vFW_PlM(107) => \b7_vFW_PlM[107]\, b7_vFW_PlM(106) => 
        \b7_vFW_PlM[106]\, b7_vFW_PlM(105) => \b7_vFW_PlM[105]\, 
        b7_vFW_PlM(104) => \b7_vFW_PlM[104]\, b7_vFW_PlM(103) => 
        \b7_vFW_PlM[103]\, b7_vFW_PlM(102) => \b7_vFW_PlM[102]\, 
        b7_vFW_PlM(101) => \b7_vFW_PlM[101]\, b7_vFW_PlM(100) => 
        \b7_vFW_PlM[100]\, b7_vFW_PlM(99) => \b7_vFW_PlM[99]\, 
        b7_vFW_PlM(98) => \b7_vFW_PlM[98]\, b7_vFW_PlM(97) => 
        \b7_vFW_PlM[97]\, b7_vFW_PlM(96) => \b7_vFW_PlM[96]\, 
        b7_vFW_PlM(95) => \b7_vFW_PlM[95]\, b7_vFW_PlM(94) => 
        \b7_vFW_PlM[94]\, b7_vFW_PlM(93) => \b7_vFW_PlM[93]\, 
        b7_vFW_PlM(92) => \b7_vFW_PlM[92]\, b7_vFW_PlM(91) => 
        \b7_vFW_PlM[91]\, b7_vFW_PlM(90) => \b7_vFW_PlM[90]\, 
        b7_vFW_PlM(89) => \b7_vFW_PlM[89]\, b7_vFW_PlM(88) => 
        \b7_vFW_PlM[88]\, b7_vFW_PlM(87) => \b7_vFW_PlM[87]\, 
        b7_vFW_PlM(86) => \b7_vFW_PlM[86]\, b7_vFW_PlM(85) => 
        \b7_vFW_PlM[85]\, b7_vFW_PlM(84) => \b7_vFW_PlM[84]\, 
        b7_vFW_PlM(83) => \b7_vFW_PlM[83]\, b7_vFW_PlM(82) => 
        \b7_vFW_PlM[82]\, b7_vFW_PlM(81) => \b7_vFW_PlM[81]\, 
        b7_vFW_PlM(80) => \b7_vFW_PlM[80]\, b7_vFW_PlM(79) => 
        \b7_vFW_PlM[79]\, b7_vFW_PlM(78) => \b7_vFW_PlM[78]\, 
        b7_vFW_PlM(77) => \b7_vFW_PlM[77]\, b7_vFW_PlM(76) => 
        \b7_vFW_PlM[76]\, b7_vFW_PlM(75) => \b7_vFW_PlM[75]\, 
        b7_vFW_PlM(74) => \b7_vFW_PlM[74]\, b7_vFW_PlM(73) => 
        \b7_vFW_PlM[73]\, b7_vFW_PlM(72) => \b7_vFW_PlM[72]\, 
        b7_vFW_PlM(71) => \b7_vFW_PlM[71]\, b7_vFW_PlM(70) => 
        \b7_vFW_PlM[70]\, b7_vFW_PlM(69) => \b7_vFW_PlM[69]\, 
        b7_vFW_PlM(68) => \b7_vFW_PlM[68]\, b7_vFW_PlM(67) => 
        \b7_vFW_PlM[67]\, b7_vFW_PlM(66) => \b7_vFW_PlM[66]\, 
        b7_vFW_PlM(65) => \b7_vFW_PlM[65]\, b7_vFW_PlM(64) => 
        \b7_vFW_PlM[64]\, b7_vFW_PlM(63) => \b7_vFW_PlM[63]\, 
        b7_vFW_PlM(62) => \b7_vFW_PlM[62]\, b7_vFW_PlM(61) => 
        \b7_vFW_PlM[61]\, b7_vFW_PlM(60) => \b7_vFW_PlM[60]\, 
        b7_vFW_PlM(59) => \b7_vFW_PlM[59]\, b7_vFW_PlM(58) => 
        \b7_vFW_PlM[58]\, b7_vFW_PlM(57) => \b7_vFW_PlM[57]\, 
        b7_vFW_PlM(56) => \b7_vFW_PlM[56]\, b7_vFW_PlM(55) => 
        \b7_vFW_PlM[55]\, b7_vFW_PlM(54) => \b7_vFW_PlM[54]\, 
        b7_vFW_PlM(53) => \b7_vFW_PlM[53]\, b7_vFW_PlM(52) => 
        \b7_vFW_PlM[52]\, b7_vFW_PlM(51) => \b7_vFW_PlM[51]\, 
        b7_vFW_PlM(50) => \b7_vFW_PlM[50]\, b7_vFW_PlM(49) => 
        \b7_vFW_PlM[49]\, b7_vFW_PlM(48) => \b7_vFW_PlM[48]\, 
        b7_vFW_PlM(47) => \b7_vFW_PlM[47]\, b7_vFW_PlM(46) => 
        \b7_vFW_PlM[46]\, b7_vFW_PlM(45) => \b7_vFW_PlM[45]\, 
        b7_vFW_PlM(44) => \b7_vFW_PlM[44]\, b7_vFW_PlM(43) => 
        \b7_vFW_PlM[43]\, b7_vFW_PlM(42) => \b7_vFW_PlM[42]\, 
        b7_vFW_PlM(41) => \b7_vFW_PlM[41]\, b7_vFW_PlM(40) => 
        \b7_vFW_PlM[40]\, b7_vFW_PlM(39) => \b7_vFW_PlM[39]\, 
        b7_vFW_PlM(38) => \b7_vFW_PlM[38]\, b7_vFW_PlM(37) => 
        \b7_vFW_PlM[37]\, b7_vFW_PlM(36) => \b7_vFW_PlM[36]\, 
        b7_vFW_PlM(35) => \b7_vFW_PlM[35]\, b7_vFW_PlM(34) => 
        \b7_vFW_PlM[34]\, b7_vFW_PlM(33) => \b7_vFW_PlM[33]\, 
        b7_vFW_PlM(32) => \b7_vFW_PlM[32]\, b7_vFW_PlM(31) => 
        \b7_vFW_PlM[31]\, b7_vFW_PlM(30) => \b7_vFW_PlM[30]\, 
        b7_vFW_PlM(29) => \b7_vFW_PlM[29]\, b7_vFW_PlM(28) => 
        \b7_vFW_PlM[28]\, b7_vFW_PlM(27) => \b7_vFW_PlM[27]\, 
        b7_vFW_PlM(26) => \b7_vFW_PlM[26]\, b7_vFW_PlM(25) => 
        \b7_vFW_PlM[25]\, b7_vFW_PlM(24) => \b7_vFW_PlM[24]\, 
        b7_vFW_PlM(23) => \b7_vFW_PlM[23]\, b7_vFW_PlM(22) => 
        \b7_vFW_PlM[22]\, b7_vFW_PlM(21) => \b7_vFW_PlM[21]\, 
        b7_vFW_PlM(20) => \b7_vFW_PlM[20]\, b7_vFW_PlM(19) => 
        \b7_vFW_PlM[19]\, b7_vFW_PlM(18) => \b7_vFW_PlM[18]\, 
        b7_vFW_PlM(17) => \b7_vFW_PlM[17]\, b7_vFW_PlM(16) => 
        \b7_vFW_PlM[16]\, b7_vFW_PlM(15) => \b7_vFW_PlM[15]\, 
        b7_vFW_PlM(14) => \b7_vFW_PlM[14]\, b7_vFW_PlM(13) => 
        \b7_vFW_PlM[13]\, b7_vFW_PlM(12) => \b7_vFW_PlM[12]\, 
        b7_vFW_PlM(11) => \b7_vFW_PlM[11]\, b7_vFW_PlM(10) => 
        \b7_vFW_PlM[10]\, b7_vFW_PlM(9) => \b7_vFW_PlM[9]\, 
        b7_vFW_PlM(8) => \b7_vFW_PlM[8]\, b7_vFW_PlM(7) => 
        \b7_vFW_PlM[7]\, b7_vFW_PlM(6) => \b7_vFW_PlM[6]\, 
        b7_vFW_PlM(5) => \b7_vFW_PlM[5]\, b7_vFW_PlM(4) => 
        \b7_vFW_PlM[4]\, b7_vFW_PlM(3) => \b7_vFW_PlM[3]\, 
        b7_vFW_PlM(2) => \b7_vFW_PlM[2]\, b7_vFW_PlM(1) => 
        \b7_vFW_PlM[1]\, b7_vFW_PlM(0) => \b7_vFW_PlM[0]\, 
        b12_2_St6KCa_jHv(11) => \b12_2_St6KCa_jHv[11]_net_1\, 
        b12_2_St6KCa_jHv(10) => \b12_2_St6KCa_jHv[10]_net_1\, 
        b12_2_St6KCa_jHv(9) => \b12_2_St6KCa_jHv[9]_net_1\, 
        b12_2_St6KCa_jHv(8) => \b12_2_St6KCa_jHv[8]_net_1\, 
        b12_2_St6KCa_jHv(7) => \b12_2_St6KCa_jHv[7]_net_1\, 
        b12_2_St6KCa_jHv(6) => \b12_2_St6KCa_jHv[6]_net_1\, 
        b12_2_St6KCa_jHv(5) => \b12_2_St6KCa_jHv[5]_net_1\, 
        b12_2_St6KCa_jHv(4) => \b12_2_St6KCa_jHv[4]_net_1\, 
        b12_2_St6KCa_jHv(3) => \b12_2_St6KCa_jHv[3]_net_1\, 
        b12_2_St6KCa_jHv(2) => \b12_2_St6KCa_jHv[2]_net_1\, 
        b12_2_St6KCa_jHv(1) => \b12_2_St6KCa_jHv[1]_net_1\, 
        b12_2_St6KCa_jHv(0) => \b12_2_St6KCa_jHv[0]_net_1\, 
        b9_v_mzCDYXs(11) => \b9_v_mzCDYXs[11]\, b9_v_mzCDYXs(10)
         => \b9_v_mzCDYXs[10]\, b9_v_mzCDYXs(9) => 
        \b9_v_mzCDYXs[9]\, b9_v_mzCDYXs(8) => \b9_v_mzCDYXs[8]\, 
        b9_v_mzCDYXs(7) => \b9_v_mzCDYXs[7]\, b9_v_mzCDYXs(6) => 
        \b9_v_mzCDYXs[6]\, b9_v_mzCDYXs(5) => \b9_v_mzCDYXs[5]\, 
        b9_v_mzCDYXs(4) => \b9_v_mzCDYXs[4]\, b9_v_mzCDYXs(3) => 
        \b9_v_mzCDYXs[3]\, b9_v_mzCDYXs(2) => \b9_v_mzCDYXs[2]\, 
        b9_v_mzCDYXs(1) => \b9_v_mzCDYXs[1]\, b9_v_mzCDYXs(0) => 
        \b9_v_mzCDYXs[0]\, IICE_comm2iice_0 => IICE_comm2iice(11), 
        b4_2o_z => b4_2o_z, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0);
    
    \genblk9.b3_PfG[49]\ : SLE
      port map(D => \b3_PfG_6[49]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[49]\);
    
    \genblk9.b3_PfG_RNO[5]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[6]\, C => 
        \b7_vFW_PlM[4]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[5]\);
    
    \b12_PSyi_KyDbLbb[10]\ : SLE
      port map(D => \b12_2_St6KCa_jHv[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \b12_PSyi_KyDbLbb_0_sqmuxa\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \b12_PSyi_KyDbLbb[10]_net_1\);
    
    \genblk9.b3_PfG_RNO[58]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[59]\, C => 
        \b7_vFW_PlM[57]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[58]\);
    
    \genblk9.b7_nYJ_BFM[45]\ : SLE
      port map(D => \b7_nYJ_BFM[44]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[45]\);
    
    \b12_2_St6KCa_jHv_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \b12_2_St6KCa_jHv[10]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \b12_2_St6KCa_jHv_cry[9]_net_1\, S => 
        \b12_2_St6KCa_jHv_s[10]\, Y => OPEN, FCO => 
        \b12_2_St6KCa_jHv_cry[10]_net_1\);
    
    \genblk9.b9_v_mzCDYXs[11]\ : SLE
      port map(D => \b9_v_mzCDYXs_s[11]\, CLK => 
        IICE_comm2iice(11), EN => b9_v_mzCDYXs13, ALn => 
        b5_voSc3_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \b9_v_mzCDYXs[11]\);
    
    virOut : b19_nczQ_DYg_YFaRM_oUoP_32s_1s_x_0
      port map(IICE_comm2iice_5 => IICE_comm2iice(11), 
        IICE_comm2iice_3 => IICE_comm2iice(9), IICE_comm2iice_0
         => IICE_comm2iice(6), IICE_comm2iice_4 => 
        IICE_comm2iice(10), N_1261_i => N_1261_i, ttdo => ttdo, 
        b7_yYh03wy5 => b7_yYh03wy5, b7_yYh03wy4 => b7_yYh03wy4);
    
    \genblk9.b3_PfG[28]\ : SLE
      port map(D => \b3_PfG_6[28]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[28]\);
    
    \genblk9.b3_PfG[119]\ : SLE
      port map(D => \b3_PfG_6[119]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[119]\);
    
    \genblk9.b3_PfG_RNO[140]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[141]\, C => 
        \b7_vFW_PlM[139]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[140]\);
    
    \genblk9.b3_PfG[3]\ : SLE
      port map(D => \b3_PfG_6[3]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[3]\);
    
    b6_SoWyQD : b11_SoWyP0zEFKY_Z2_x_0
      port map(mdiclink_reg(167) => mdiclink_reg(167), 
        mdiclink_reg(166) => mdiclink_reg(166), mdiclink_reg(165)
         => mdiclink_reg(165), mdiclink_reg(164) => 
        mdiclink_reg(164), mdiclink_reg(163) => mdiclink_reg(163), 
        mdiclink_reg(162) => mdiclink_reg(162), mdiclink_reg(161)
         => mdiclink_reg(161), mdiclink_reg(160) => 
        mdiclink_reg(160), mdiclink_reg(159) => mdiclink_reg(159), 
        mdiclink_reg(158) => mdiclink_reg(158), mdiclink_reg(157)
         => mdiclink_reg(157), mdiclink_reg(156) => 
        mdiclink_reg(156), mdiclink_reg(155) => mdiclink_reg(155), 
        mdiclink_reg(154) => mdiclink_reg(154), mdiclink_reg(153)
         => mdiclink_reg(153), mdiclink_reg(152) => 
        mdiclink_reg(152), mdiclink_reg(151) => mdiclink_reg(151), 
        mdiclink_reg(150) => mdiclink_reg(150), mdiclink_reg(149)
         => mdiclink_reg(149), mdiclink_reg(148) => 
        mdiclink_reg(148), mdiclink_reg(147) => mdiclink_reg(147), 
        mdiclink_reg(146) => mdiclink_reg(146), mdiclink_reg(145)
         => mdiclink_reg(145), mdiclink_reg(144) => 
        mdiclink_reg(144), mdiclink_reg(143) => mdiclink_reg(143), 
        mdiclink_reg(142) => mdiclink_reg(142), mdiclink_reg(141)
         => mdiclink_reg(141), mdiclink_reg(140) => 
        mdiclink_reg(140), mdiclink_reg(139) => mdiclink_reg(139), 
        mdiclink_reg(138) => mdiclink_reg(138), mdiclink_reg(137)
         => mdiclink_reg(137), mdiclink_reg(136) => 
        mdiclink_reg(136), mdiclink_reg(135) => mdiclink_reg(135), 
        mdiclink_reg(134) => mdiclink_reg(134), mdiclink_reg(133)
         => mdiclink_reg(133), mdiclink_reg(132) => 
        mdiclink_reg(132), mdiclink_reg(131) => mdiclink_reg(131), 
        mdiclink_reg(130) => mdiclink_reg(130), mdiclink_reg(129)
         => mdiclink_reg(129), mdiclink_reg(128) => 
        mdiclink_reg(128), mdiclink_reg(127) => mdiclink_reg(127), 
        mdiclink_reg(126) => mdiclink_reg(126), mdiclink_reg(125)
         => mdiclink_reg(125), mdiclink_reg(124) => 
        mdiclink_reg(124), mdiclink_reg(123) => mdiclink_reg(123), 
        mdiclink_reg(122) => mdiclink_reg(122), mdiclink_reg(121)
         => mdiclink_reg(121), mdiclink_reg(120) => 
        mdiclink_reg(120), mdiclink_reg(119) => mdiclink_reg(119), 
        mdiclink_reg(118) => mdiclink_reg(118), mdiclink_reg(117)
         => mdiclink_reg(117), mdiclink_reg(116) => 
        mdiclink_reg(116), mdiclink_reg(115) => mdiclink_reg(115), 
        mdiclink_reg(114) => mdiclink_reg(114), mdiclink_reg(113)
         => mdiclink_reg(113), mdiclink_reg(112) => 
        mdiclink_reg(112), mdiclink_reg(111) => mdiclink_reg(111), 
        mdiclink_reg(110) => mdiclink_reg(110), mdiclink_reg(109)
         => mdiclink_reg(109), mdiclink_reg(108) => 
        mdiclink_reg(108), mdiclink_reg(107) => mdiclink_reg(107), 
        mdiclink_reg(106) => mdiclink_reg(106), mdiclink_reg(105)
         => mdiclink_reg(105), mdiclink_reg(104) => 
        mdiclink_reg(104), mdiclink_reg(103) => mdiclink_reg(103), 
        mdiclink_reg(102) => mdiclink_reg(102), mdiclink_reg(101)
         => mdiclink_reg(101), mdiclink_reg(100) => 
        mdiclink_reg(100), mdiclink_reg(99) => mdiclink_reg(99), 
        mdiclink_reg(98) => mdiclink_reg(98), mdiclink_reg(97)
         => mdiclink_reg(97), mdiclink_reg(96) => 
        mdiclink_reg(96), mdiclink_reg(95) => mdiclink_reg(95), 
        mdiclink_reg(94) => mdiclink_reg(94), mdiclink_reg(93)
         => mdiclink_reg(93), mdiclink_reg(92) => 
        mdiclink_reg(92), mdiclink_reg(91) => mdiclink_reg(91), 
        mdiclink_reg(90) => mdiclink_reg(90), mdiclink_reg(89)
         => mdiclink_reg(89), mdiclink_reg(88) => 
        mdiclink_reg(88), mdiclink_reg(87) => mdiclink_reg(87), 
        mdiclink_reg(86) => mdiclink_reg(86), mdiclink_reg(85)
         => mdiclink_reg(85), mdiclink_reg(84) => 
        mdiclink_reg(84), mdiclink_reg(83) => mdiclink_reg(83), 
        mdiclink_reg(82) => mdiclink_reg(82), mdiclink_reg(81)
         => mdiclink_reg(81), mdiclink_reg(80) => 
        mdiclink_reg(80), mdiclink_reg(79) => mdiclink_reg(79), 
        mdiclink_reg(78) => mdiclink_reg(78), mdiclink_reg(77)
         => mdiclink_reg(77), mdiclink_reg(76) => 
        mdiclink_reg(76), mdiclink_reg(75) => mdiclink_reg(75), 
        mdiclink_reg(74) => mdiclink_reg(74), mdiclink_reg(73)
         => mdiclink_reg(73), mdiclink_reg(72) => 
        mdiclink_reg(72), mdiclink_reg(71) => mdiclink_reg(71), 
        mdiclink_reg(70) => mdiclink_reg(70), mdiclink_reg(69)
         => mdiclink_reg(69), mdiclink_reg(68) => 
        mdiclink_reg(68), mdiclink_reg(67) => mdiclink_reg(67), 
        mdiclink_reg(66) => mdiclink_reg(66), mdiclink_reg(65)
         => mdiclink_reg(65), mdiclink_reg(64) => 
        mdiclink_reg(64), mdiclink_reg(63) => mdiclink_reg(63), 
        mdiclink_reg(62) => mdiclink_reg(62), mdiclink_reg(61)
         => mdiclink_reg(61), mdiclink_reg(60) => 
        mdiclink_reg(60), mdiclink_reg(59) => mdiclink_reg(59), 
        mdiclink_reg(58) => mdiclink_reg(58), mdiclink_reg(57)
         => mdiclink_reg(57), mdiclink_reg(56) => 
        mdiclink_reg(56), mdiclink_reg(55) => mdiclink_reg(55), 
        mdiclink_reg(54) => mdiclink_reg(54), mdiclink_reg(53)
         => mdiclink_reg(53), mdiclink_reg(52) => 
        mdiclink_reg(52), mdiclink_reg(51) => mdiclink_reg(51), 
        mdiclink_reg(50) => mdiclink_reg(50), mdiclink_reg(49)
         => mdiclink_reg(49), mdiclink_reg(48) => 
        mdiclink_reg(48), mdiclink_reg(47) => mdiclink_reg(47), 
        mdiclink_reg(46) => mdiclink_reg(46), mdiclink_reg(45)
         => mdiclink_reg(45), mdiclink_reg(44) => 
        mdiclink_reg(44), mdiclink_reg(43) => mdiclink_reg(43), 
        mdiclink_reg(42) => mdiclink_reg(42), mdiclink_reg(41)
         => mdiclink_reg(41), mdiclink_reg(40) => 
        mdiclink_reg(40), mdiclink_reg(39) => mdiclink_reg(39), 
        mdiclink_reg(38) => mdiclink_reg(38), mdiclink_reg(37)
         => mdiclink_reg(37), mdiclink_reg(36) => 
        mdiclink_reg(36), mdiclink_reg(35) => mdiclink_reg(35), 
        mdiclink_reg(34) => mdiclink_reg(34), mdiclink_reg(33)
         => mdiclink_reg(33), mdiclink_reg(32) => 
        mdiclink_reg(32), mdiclink_reg(31) => mdiclink_reg(31), 
        mdiclink_reg(30) => mdiclink_reg(30), mdiclink_reg(29)
         => mdiclink_reg(29), mdiclink_reg(28) => 
        mdiclink_reg(28), mdiclink_reg(27) => mdiclink_reg(27), 
        mdiclink_reg(26) => mdiclink_reg(26), mdiclink_reg(25)
         => mdiclink_reg(25), mdiclink_reg(24) => 
        mdiclink_reg(24), mdiclink_reg(23) => mdiclink_reg(23), 
        mdiclink_reg(22) => mdiclink_reg(22), mdiclink_reg(21)
         => mdiclink_reg(21), mdiclink_reg(20) => 
        mdiclink_reg(20), mdiclink_reg(19) => mdiclink_reg(19), 
        mdiclink_reg(18) => mdiclink_reg(18), mdiclink_reg(17)
         => mdiclink_reg(17), mdiclink_reg(16) => 
        mdiclink_reg(16), mdiclink_reg(15) => mdiclink_reg(15), 
        mdiclink_reg(14) => mdiclink_reg(14), mdiclink_reg(13)
         => mdiclink_reg(13), mdiclink_reg(12) => 
        mdiclink_reg(12), mdiclink_reg(11) => mdiclink_reg(11), 
        mdiclink_reg(10) => mdiclink_reg(10), mdiclink_reg(9) => 
        mdiclink_reg(9), mdiclink_reg(8) => mdiclink_reg(8), 
        mdiclink_reg(7) => mdiclink_reg(7), mdiclink_reg(6) => 
        mdiclink_reg(6), mdiclink_reg(5) => mdiclink_reg(5), 
        mdiclink_reg(4) => mdiclink_reg(4), mdiclink_reg(3) => 
        mdiclink_reg(3), mdiclink_reg(2) => mdiclink_reg(2), 
        mdiclink_reg(1) => mdiclink_reg(1), mdiclink_reg(0) => 
        mdiclink_reg(0), b11_OFWNT9L_8tZ(167) => 
        \b11_OFWNT9L_8tZ[167]\, b11_OFWNT9L_8tZ(166) => 
        \b11_OFWNT9L_8tZ[166]\, b11_OFWNT9L_8tZ(165) => 
        \b11_OFWNT9L_8tZ[165]\, b11_OFWNT9L_8tZ(164) => 
        \b11_OFWNT9L_8tZ[164]\, b11_OFWNT9L_8tZ(163) => 
        \b11_OFWNT9L_8tZ[163]\, b11_OFWNT9L_8tZ(162) => 
        \b11_OFWNT9L_8tZ[162]\, b11_OFWNT9L_8tZ(161) => 
        \b11_OFWNT9L_8tZ[161]\, b11_OFWNT9L_8tZ(160) => 
        \b11_OFWNT9L_8tZ[160]\, b11_OFWNT9L_8tZ(159) => 
        \b11_OFWNT9L_8tZ[159]\, b11_OFWNT9L_8tZ(158) => 
        \b11_OFWNT9L_8tZ[158]\, b11_OFWNT9L_8tZ(157) => 
        \b11_OFWNT9L_8tZ[157]\, b11_OFWNT9L_8tZ(156) => 
        \b11_OFWNT9L_8tZ[156]\, b11_OFWNT9L_8tZ(155) => 
        \b11_OFWNT9L_8tZ[155]\, b11_OFWNT9L_8tZ(154) => 
        \b11_OFWNT9L_8tZ[154]\, b11_OFWNT9L_8tZ(153) => 
        \b11_OFWNT9L_8tZ[153]\, b11_OFWNT9L_8tZ(152) => 
        \b11_OFWNT9L_8tZ[152]\, b11_OFWNT9L_8tZ(151) => 
        \b11_OFWNT9L_8tZ[151]\, b11_OFWNT9L_8tZ(150) => 
        \b11_OFWNT9L_8tZ[150]\, b11_OFWNT9L_8tZ(149) => 
        \b11_OFWNT9L_8tZ[149]\, b11_OFWNT9L_8tZ(148) => 
        \b11_OFWNT9L_8tZ[148]\, b11_OFWNT9L_8tZ(147) => 
        \b11_OFWNT9L_8tZ[147]\, b11_OFWNT9L_8tZ(146) => 
        \b11_OFWNT9L_8tZ[146]\, b11_OFWNT9L_8tZ(145) => 
        \b11_OFWNT9L_8tZ[145]\, b11_OFWNT9L_8tZ(144) => 
        \b11_OFWNT9L_8tZ[144]\, b11_OFWNT9L_8tZ(143) => 
        \b11_OFWNT9L_8tZ[143]\, b11_OFWNT9L_8tZ(142) => 
        \b11_OFWNT9L_8tZ[142]\, b11_OFWNT9L_8tZ(141) => 
        \b11_OFWNT9L_8tZ[141]\, b11_OFWNT9L_8tZ(140) => 
        \b11_OFWNT9L_8tZ[140]\, b11_OFWNT9L_8tZ(139) => 
        \b11_OFWNT9L_8tZ[139]\, b11_OFWNT9L_8tZ(138) => 
        \b11_OFWNT9L_8tZ[138]\, b11_OFWNT9L_8tZ(137) => 
        \b11_OFWNT9L_8tZ[137]\, b11_OFWNT9L_8tZ(136) => 
        \b11_OFWNT9L_8tZ[136]\, b11_OFWNT9L_8tZ(135) => 
        \b11_OFWNT9L_8tZ[135]\, b11_OFWNT9L_8tZ(134) => 
        \b11_OFWNT9L_8tZ[134]\, b11_OFWNT9L_8tZ(133) => 
        \b11_OFWNT9L_8tZ[133]\, b11_OFWNT9L_8tZ(132) => 
        \b11_OFWNT9L_8tZ[132]\, b11_OFWNT9L_8tZ(131) => 
        \b11_OFWNT9L_8tZ[131]\, b11_OFWNT9L_8tZ(130) => 
        \b11_OFWNT9L_8tZ[130]\, b11_OFWNT9L_8tZ(129) => 
        \b11_OFWNT9L_8tZ[129]\, b11_OFWNT9L_8tZ(128) => 
        \b11_OFWNT9L_8tZ[128]\, b11_OFWNT9L_8tZ(127) => 
        \b11_OFWNT9L_8tZ[127]\, b11_OFWNT9L_8tZ(126) => 
        \b11_OFWNT9L_8tZ[126]\, b11_OFWNT9L_8tZ(125) => 
        \b11_OFWNT9L_8tZ[125]\, b11_OFWNT9L_8tZ(124) => 
        \b11_OFWNT9L_8tZ[124]\, b11_OFWNT9L_8tZ(123) => 
        \b11_OFWNT9L_8tZ[123]\, b11_OFWNT9L_8tZ(122) => 
        \b11_OFWNT9L_8tZ[122]\, b11_OFWNT9L_8tZ(121) => 
        \b11_OFWNT9L_8tZ[121]\, b11_OFWNT9L_8tZ(120) => 
        \b11_OFWNT9L_8tZ[120]\, b11_OFWNT9L_8tZ(119) => 
        \b11_OFWNT9L_8tZ[119]\, b11_OFWNT9L_8tZ(118) => 
        \b11_OFWNT9L_8tZ[118]\, b11_OFWNT9L_8tZ(117) => 
        \b11_OFWNT9L_8tZ[117]\, b11_OFWNT9L_8tZ(116) => 
        \b11_OFWNT9L_8tZ[116]\, b11_OFWNT9L_8tZ(115) => 
        \b11_OFWNT9L_8tZ[115]\, b11_OFWNT9L_8tZ(114) => 
        \b11_OFWNT9L_8tZ[114]\, b11_OFWNT9L_8tZ(113) => 
        \b11_OFWNT9L_8tZ[113]\, b11_OFWNT9L_8tZ(112) => 
        \b11_OFWNT9L_8tZ[112]\, b11_OFWNT9L_8tZ(111) => 
        \b11_OFWNT9L_8tZ[111]\, b11_OFWNT9L_8tZ(110) => 
        \b11_OFWNT9L_8tZ[110]\, b11_OFWNT9L_8tZ(109) => 
        \b11_OFWNT9L_8tZ[109]\, b11_OFWNT9L_8tZ(108) => 
        \b11_OFWNT9L_8tZ[108]\, b11_OFWNT9L_8tZ(107) => 
        \b11_OFWNT9L_8tZ[107]\, b11_OFWNT9L_8tZ(106) => 
        \b11_OFWNT9L_8tZ[106]\, b11_OFWNT9L_8tZ(105) => 
        \b11_OFWNT9L_8tZ[105]\, b11_OFWNT9L_8tZ(104) => 
        \b11_OFWNT9L_8tZ[104]\, b11_OFWNT9L_8tZ(103) => 
        \b11_OFWNT9L_8tZ[103]\, b11_OFWNT9L_8tZ(102) => 
        \b11_OFWNT9L_8tZ[102]\, b11_OFWNT9L_8tZ(101) => 
        \b11_OFWNT9L_8tZ[101]\, b11_OFWNT9L_8tZ(100) => 
        \b11_OFWNT9L_8tZ[100]\, b11_OFWNT9L_8tZ(99) => 
        \b11_OFWNT9L_8tZ[99]\, b11_OFWNT9L_8tZ(98) => 
        \b11_OFWNT9L_8tZ[98]\, b11_OFWNT9L_8tZ(97) => 
        \b11_OFWNT9L_8tZ[97]\, b11_OFWNT9L_8tZ(96) => 
        \b11_OFWNT9L_8tZ[96]\, b11_OFWNT9L_8tZ(95) => 
        \b11_OFWNT9L_8tZ[95]\, b11_OFWNT9L_8tZ(94) => 
        \b11_OFWNT9L_8tZ[94]\, b11_OFWNT9L_8tZ(93) => 
        \b11_OFWNT9L_8tZ[93]\, b11_OFWNT9L_8tZ(92) => 
        \b11_OFWNT9L_8tZ[92]\, b11_OFWNT9L_8tZ(91) => 
        \b11_OFWNT9L_8tZ[91]\, b11_OFWNT9L_8tZ(90) => 
        \b11_OFWNT9L_8tZ[90]\, b11_OFWNT9L_8tZ(89) => 
        \b11_OFWNT9L_8tZ[89]\, b11_OFWNT9L_8tZ(88) => 
        \b11_OFWNT9L_8tZ[88]\, b11_OFWNT9L_8tZ(87) => 
        \b11_OFWNT9L_8tZ[87]\, b11_OFWNT9L_8tZ(86) => 
        \b11_OFWNT9L_8tZ[86]\, b11_OFWNT9L_8tZ(85) => 
        \b11_OFWNT9L_8tZ[85]\, b11_OFWNT9L_8tZ(84) => 
        \b11_OFWNT9L_8tZ[84]\, b11_OFWNT9L_8tZ(83) => 
        \b11_OFWNT9L_8tZ[83]\, b11_OFWNT9L_8tZ(82) => 
        \b11_OFWNT9L_8tZ[82]\, b11_OFWNT9L_8tZ(81) => 
        \b11_OFWNT9L_8tZ[81]\, b11_OFWNT9L_8tZ(80) => 
        \b11_OFWNT9L_8tZ[80]\, b11_OFWNT9L_8tZ(79) => 
        \b11_OFWNT9L_8tZ[79]\, b11_OFWNT9L_8tZ(78) => 
        \b11_OFWNT9L_8tZ[78]\, b11_OFWNT9L_8tZ(77) => 
        \b11_OFWNT9L_8tZ[77]\, b11_OFWNT9L_8tZ(76) => 
        \b11_OFWNT9L_8tZ[76]\, b11_OFWNT9L_8tZ(75) => 
        \b11_OFWNT9L_8tZ[75]\, b11_OFWNT9L_8tZ(74) => 
        \b11_OFWNT9L_8tZ[74]\, b11_OFWNT9L_8tZ(73) => 
        \b11_OFWNT9L_8tZ[73]\, b11_OFWNT9L_8tZ(72) => 
        \b11_OFWNT9L_8tZ[72]\, b11_OFWNT9L_8tZ(71) => 
        \b11_OFWNT9L_8tZ[71]\, b11_OFWNT9L_8tZ(70) => 
        \b11_OFWNT9L_8tZ[70]\, b11_OFWNT9L_8tZ(69) => 
        \b11_OFWNT9L_8tZ[69]\, b11_OFWNT9L_8tZ(68) => 
        \b11_OFWNT9L_8tZ[68]\, b11_OFWNT9L_8tZ(67) => 
        \b11_OFWNT9L_8tZ[67]\, b11_OFWNT9L_8tZ(66) => 
        \b11_OFWNT9L_8tZ[66]\, b11_OFWNT9L_8tZ(65) => 
        \b11_OFWNT9L_8tZ[65]\, b11_OFWNT9L_8tZ(64) => 
        \b11_OFWNT9L_8tZ[64]\, b11_OFWNT9L_8tZ(63) => 
        \b11_OFWNT9L_8tZ[63]\, b11_OFWNT9L_8tZ(62) => 
        \b11_OFWNT9L_8tZ[62]\, b11_OFWNT9L_8tZ(61) => 
        \b11_OFWNT9L_8tZ[61]\, b11_OFWNT9L_8tZ(60) => 
        \b11_OFWNT9L_8tZ[60]\, b11_OFWNT9L_8tZ(59) => 
        \b11_OFWNT9L_8tZ[59]\, b11_OFWNT9L_8tZ(58) => 
        \b11_OFWNT9L_8tZ[58]\, b11_OFWNT9L_8tZ(57) => 
        \b11_OFWNT9L_8tZ[57]\, b11_OFWNT9L_8tZ(56) => 
        \b11_OFWNT9L_8tZ[56]\, b11_OFWNT9L_8tZ(55) => 
        \b11_OFWNT9L_8tZ[55]\, b11_OFWNT9L_8tZ(54) => 
        \b11_OFWNT9L_8tZ[54]\, b11_OFWNT9L_8tZ(53) => 
        \b11_OFWNT9L_8tZ[53]\, b11_OFWNT9L_8tZ(52) => 
        \b11_OFWNT9L_8tZ[52]\, b11_OFWNT9L_8tZ(51) => 
        \b11_OFWNT9L_8tZ[51]\, b11_OFWNT9L_8tZ(50) => 
        \b11_OFWNT9L_8tZ[50]\, b11_OFWNT9L_8tZ(49) => 
        \b11_OFWNT9L_8tZ[49]\, b11_OFWNT9L_8tZ(48) => 
        \b11_OFWNT9L_8tZ[48]\, b11_OFWNT9L_8tZ(47) => 
        \b11_OFWNT9L_8tZ[47]\, b11_OFWNT9L_8tZ(46) => 
        \b11_OFWNT9L_8tZ[46]\, b11_OFWNT9L_8tZ(45) => 
        \b11_OFWNT9L_8tZ[45]\, b11_OFWNT9L_8tZ(44) => 
        \b11_OFWNT9L_8tZ[44]\, b11_OFWNT9L_8tZ(43) => 
        \b11_OFWNT9L_8tZ[43]\, b11_OFWNT9L_8tZ(42) => 
        \b11_OFWNT9L_8tZ[42]\, b11_OFWNT9L_8tZ(41) => 
        \b11_OFWNT9L_8tZ[41]\, b11_OFWNT9L_8tZ(40) => 
        \b11_OFWNT9L_8tZ[40]\, b11_OFWNT9L_8tZ(39) => 
        \b11_OFWNT9L_8tZ[39]\, b11_OFWNT9L_8tZ(38) => 
        \b11_OFWNT9L_8tZ[38]\, b11_OFWNT9L_8tZ(37) => 
        \b11_OFWNT9L_8tZ[37]\, b11_OFWNT9L_8tZ(36) => 
        \b11_OFWNT9L_8tZ[36]\, b11_OFWNT9L_8tZ(35) => 
        \b11_OFWNT9L_8tZ[35]\, b11_OFWNT9L_8tZ(34) => 
        \b11_OFWNT9L_8tZ[34]\, b11_OFWNT9L_8tZ(33) => 
        \b11_OFWNT9L_8tZ[33]\, b11_OFWNT9L_8tZ(32) => 
        \b11_OFWNT9L_8tZ[32]\, b11_OFWNT9L_8tZ(31) => 
        \b11_OFWNT9L_8tZ[31]\, b11_OFWNT9L_8tZ(30) => 
        \b11_OFWNT9L_8tZ[30]\, b11_OFWNT9L_8tZ(29) => 
        \b11_OFWNT9L_8tZ[29]\, b11_OFWNT9L_8tZ(28) => 
        \b11_OFWNT9L_8tZ[28]\, b11_OFWNT9L_8tZ(27) => 
        \b11_OFWNT9L_8tZ[27]\, b11_OFWNT9L_8tZ(26) => 
        \b11_OFWNT9L_8tZ[26]\, b11_OFWNT9L_8tZ(25) => 
        \b11_OFWNT9L_8tZ[25]\, b11_OFWNT9L_8tZ(24) => 
        \b11_OFWNT9L_8tZ[24]\, b11_OFWNT9L_8tZ(23) => 
        \b11_OFWNT9L_8tZ[23]\, b11_OFWNT9L_8tZ(22) => 
        \b11_OFWNT9L_8tZ[22]\, b11_OFWNT9L_8tZ(21) => 
        \b11_OFWNT9L_8tZ[21]\, b11_OFWNT9L_8tZ(20) => 
        \b11_OFWNT9L_8tZ[20]\, b11_OFWNT9L_8tZ(19) => 
        \b11_OFWNT9L_8tZ[19]\, b11_OFWNT9L_8tZ(18) => 
        \b11_OFWNT9L_8tZ[18]\, b11_OFWNT9L_8tZ(17) => 
        \b11_OFWNT9L_8tZ[17]\, b11_OFWNT9L_8tZ(16) => 
        \b11_OFWNT9L_8tZ[16]\, b11_OFWNT9L_8tZ(15) => 
        \b11_OFWNT9L_8tZ[15]\, b11_OFWNT9L_8tZ(14) => 
        \b11_OFWNT9L_8tZ[14]\, b11_OFWNT9L_8tZ(13) => 
        \b11_OFWNT9L_8tZ[13]\, b11_OFWNT9L_8tZ(12) => 
        \b11_OFWNT9L_8tZ[12]\, b11_OFWNT9L_8tZ(11) => 
        \b11_OFWNT9L_8tZ[11]\, b11_OFWNT9L_8tZ(10) => 
        \b11_OFWNT9L_8tZ[10]\, b11_OFWNT9L_8tZ(9) => 
        \b11_OFWNT9L_8tZ[9]\, b11_OFWNT9L_8tZ(8) => 
        \b11_OFWNT9L_8tZ[8]\, b11_OFWNT9L_8tZ(7) => 
        \b11_OFWNT9L_8tZ[7]\, b11_OFWNT9L_8tZ(6) => 
        \b11_OFWNT9L_8tZ[6]\, b11_OFWNT9L_8tZ(5) => 
        \b11_OFWNT9L_8tZ[5]\, b11_OFWNT9L_8tZ(4) => 
        \b11_OFWNT9L_8tZ[4]\, b11_OFWNT9L_8tZ(3) => 
        \b11_OFWNT9L_8tZ[3]\, b11_OFWNT9L_8tZ(2) => 
        \b11_OFWNT9L_8tZ[2]\, b11_OFWNT9L_8tZ(1) => 
        \b11_OFWNT9L_8tZ[1]\, b11_OFWNT9L_8tZ(0) => 
        \b11_OFWNT9L_8tZ[0]\, N_145_i => N_145_i, b4_2o_z => 
        b4_2o_z, CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0);
    
    \genblk9.b7_nYJ_BFM[168]\ : SLE
      port map(D => \b7_nYJ_BFM[167]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[168]\);
    
    \genblk9.b3_PfG_RNO[82]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[83]\, C => 
        \b7_vFW_PlM[81]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[82]\);
    
    \genblk9.b7_nYJ_BFM[148]\ : SLE
      port map(D => \b7_nYJ_BFM[147]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[148]\);
    
    \genblk9.b3_PfG_RNO[25]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[26]\, C => 
        \b7_vFW_PlM[24]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[25]\);
    
    \genblk9.b7_nYJ_BFM[76]\ : SLE
      port map(D => \b7_nYJ_BFM[75]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[76]\);
    
    \genblk9.b7_nYJ_BFM[121]\ : SLE
      port map(D => \b7_nYJ_BFM[120]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[121]\);
    
    \b12_PSyi_KyDbLbb[5]\ : SLE
      port map(D => \b12_2_St6KCa_jHv[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \b12_PSyi_KyDbLbb_0_sqmuxa\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \b12_PSyi_KyDbLbb[5]_net_1\);
    
    \genblk9.b7_nYJ_BFM[137]\ : SLE
      port map(D => \b7_nYJ_BFM[136]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[137]\);
    
    \genblk9.b3_PfG_RNO[91]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[92]\, C => 
        \b7_vFW_PlM[90]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[91]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \genblk9.b3_PfG_RNO[90]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[91]\, C => 
        \b7_vFW_PlM[89]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[90]\);
    
    \genblk9.b7_nYJ_BFM[66]\ : SLE
      port map(D => \b7_nYJ_BFM[65]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[66]\);
    
    \genblk9.b3_PfG_RNO[120]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[121]\, C => 
        \b7_vFW_PlM[119]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[120]\);
    
    \genblk9.b9_v_mzCDYXs_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \b9_v_mzCDYXs[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => \b9_v_mzCDYXs_cry[5]\, 
        S => \b9_v_mzCDYXs_s[6]\, Y => OPEN, FCO => 
        \b9_v_mzCDYXs_cry[6]\);
    
    \genblk9.b3_PfG[141]\ : SLE
      port map(D => \b3_PfG_6[141]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[141]\);
    
    \genblk9.b7_nYJ_BFM[41]\ : SLE
      port map(D => \b7_nYJ_BFM[40]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[41]\);
    
    \genblk9.b7_nYJ_BFM[171]\ : SLE
      port map(D => \b7_nYJ_BFM[170]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[171]\);
    
    \genblk9.b9_v_mzCDYXs_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \b9_v_mzCDYXs[8]\, C => 
        GND_net_1, D => GND_net_1, FCI => \b9_v_mzCDYXs_cry[7]\, 
        S => \b9_v_mzCDYXs_s[8]\, Y => OPEN, FCO => 
        \b9_v_mzCDYXs_cry[8]\);
    
    \genblk9.b7_nYJ_BFM[82]\ : SLE
      port map(D => \b7_nYJ_BFM[81]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[82]\);
    
    \b12_PSyi_KyDbLbb[8]\ : SLE
      port map(D => \b12_2_St6KCa_jHv[8]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \b12_PSyi_KyDbLbb_0_sqmuxa\, 
        ALn => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \b12_PSyi_KyDbLbb[8]_net_1\);
    
    \genblk9.b7_nYJ_BFM[150]\ : SLE
      port map(D => \b7_nYJ_BFM[149]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[150]\);
    
    \genblk9.b3_PfG[43]\ : SLE
      port map(D => \b3_PfG_6[43]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[43]\);
    
    \genblk9.b3_PfG_RNO[65]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[66]\, C => 
        \b7_vFW_PlM[64]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[65]\);
    
    \genblk9.b7_nYJ_BFM[17]\ : SLE
      port map(D => \b7_nYJ_BFM[16]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[17]\);
    
    \genblk9.b7_nYJ_BFM[109]\ : SLE
      port map(D => \b7_nYJ_BFM[108]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[109]\);
    
    \genblk9.b3_PfG[139]\ : SLE
      port map(D => \b3_PfG_6[139]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[139]\);
    
    \genblk9.b3_PfG_RNO[45]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[46]\, C => 
        \b7_vFW_PlM[44]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[45]\);
    
    \genblk9.b3_PfG[55]\ : SLE
      port map(D => \b3_PfG_6[55]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[55]\);
    
    \genblk9.b9_v_mzCDYXs_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \b9_v_mzCDYXs[3]\, C => 
        GND_net_1, D => GND_net_1, FCI => \b9_v_mzCDYXs_cry[2]\, 
        S => \b9_v_mzCDYXs_s[3]\, Y => OPEN, FCO => 
        \b9_v_mzCDYXs_cry[3]\);
    
    \genblk9.b7_nYJ_BFM[111]\ : SLE
      port map(D => \b7_nYJ_BFM[110]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[111]\);
    
    \genblk9.b3_PfG[8]\ : SLE
      port map(D => \b3_PfG_6[8]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[8]\);
    
    \genblk9.b7_nYJ_BFM[23]\ : SLE
      port map(D => \b7_nYJ_BFM[22]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[23]\);
    
    \genblk9.b3_PfG[124]\ : SLE
      port map(D => \b3_PfG_6[124]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[124]\);
    
    \genblk9.b7_nYJ_BFM[126]\ : SLE
      port map(D => \b7_nYJ_BFM[125]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[126]\);
    
    \genblk9.b7_nYJ_BFM[96]\ : SLE
      port map(D => \b7_nYJ_BFM[95]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[96]\);
    
    \genblk9.b3_PfG_RNO[36]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[37]\, C => 
        \b7_vFW_PlM[35]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[36]\);
    
    \genblk9.b3_PfG[88]\ : SLE
      port map(D => \b3_PfG_6[88]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[88]\);
    
    \genblk9.b3_PfG[146]\ : SLE
      port map(D => \b3_PfG_6[146]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[146]\);
    
    \genblk9.b9_v_mzCDYXs[6]\ : SLE
      port map(D => \b9_v_mzCDYXs_s[6]\, CLK => 
        IICE_comm2iice(11), EN => b9_v_mzCDYXs13, ALn => 
        b5_voSc3_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \b9_v_mzCDYXs[6]\);
    
    \genblk9.b3_PfG[27]\ : SLE
      port map(D => \b3_PfG_6[27]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[27]\);
    
    \genblk9.b3_PfG[104]\ : SLE
      port map(D => \b3_PfG_6[104]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[104]\);
    
    \genblk9.b3_PfG[117]\ : SLE
      port map(D => \b3_PfG_6[117]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[117]\);
    
    \genblk9.b3_PfG[161]\ : SLE
      port map(D => \b3_PfG_6[161]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[161]\);
    
    \genblk9.b9_v_mzCDYXs_s[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \b9_v_mzCDYXs[11]\, C => 
        GND_net_1, D => GND_net_1, FCI => \b9_v_mzCDYXs_cry[10]\, 
        S => \b9_v_mzCDYXs_s[11]\, Y => OPEN, FCO => OPEN);
    
    \genblk9.b7_nYJ_BFM[105]\ : SLE
      port map(D => \b7_nYJ_BFM[104]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[105]\);
    
    \genblk9.b3_PfG_RNO[83]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[84]\, C => 
        \b7_vFW_PlM[82]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[83]\);
    
    \genblk9.b3_PfG_RNO[72]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[73]\, C => 
        \b7_vFW_PlM[71]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[72]\);
    
    \genblk9.b7_nYJ_BFM[103]\ : SLE
      port map(D => \b7_nYJ_BFM[102]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[103]\);
    
    \genblk9.b3_PfG_RNO[110]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[111]\, C => 
        \b7_vFW_PlM[109]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[110]\);
    
    \genblk9.b7_nYJ_BFM[8]\ : SLE
      port map(D => \b7_nYJ_BFM[7]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[8]\);
    
    \genblk9.b7_nYJ_BFM[24]\ : SLE
      port map(D => \b7_nYJ_BFM[23]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[24]\);
    
    \genblk9.b3_PfG[74]\ : SLE
      port map(D => \b3_PfG_6[74]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[74]\);
    
    \genblk9.b3_PfG_RNO[11]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[12]\, C => 
        \b7_vFW_PlM[10]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[11]\);
    
    \genblk9.b7_nYJ_BFM[116]\ : SLE
      port map(D => \b7_nYJ_BFM[115]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[116]\);
    
    \genblk9.b3_PfG_RNO[10]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[11]\, C => 
        \b7_vFW_PlM[9]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[10]\);
    
    \genblk9.b3_PfG[128]\ : SLE
      port map(D => \b3_PfG_6[128]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[128]\);
    
    \genblk9.b3_PfG_RNO[29]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[30]\, C => 
        \b7_vFW_PlM[28]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[29]\);
    
    \genblk9.b3_PfG_RNO[166]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[167]\, C => 
        \b7_vFW_PlM[165]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[166]\);
    
    \genblk9.b7_nYJ_BFM[104]\ : SLE
      port map(D => \b7_nYJ_BFM[103]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[104]\);
    
    \genblk9.b3_PfG[159]\ : SLE
      port map(D => \b3_PfG_6[159]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[159]\);
    
    \genblk9.b3_PfG[10]\ : SLE
      port map(D => \b3_PfG_6[10]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[10]\);
    
    \b12_2_St6KCa_jHv[7]\ : SLE
      port map(D => \b12_2_St6KCa_jHv_s[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b4_2o_z, ALn => b5_voSc3_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b12_2_St6KCa_jHv[7]_net_1\);
    
    \genblk9.b7_nYJ_BFM[131]\ : SLE
      port map(D => \b7_nYJ_BFM[130]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[131]\);
    
    \genblk9.b3_PfG[166]\ : SLE
      port map(D => \b3_PfG_6[166]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[166]\);
    
    \genblk9.b3_PfG[64]\ : SLE
      port map(D => \b3_PfG_6[64]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[64]\);
    
    \genblk9.b3_PfG[108]\ : SLE
      port map(D => \b3_PfG_6[108]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[108]\);
    
    \b12_2_St6KCa_jHv_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \b12_2_St6KCa_jHv[7]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \b12_2_St6KCa_jHv_cry[6]_net_1\, S => 
        \b12_2_St6KCa_jHv_s[7]\, Y => OPEN, FCO => 
        \b12_2_St6KCa_jHv_cry[7]_net_1\);
    
    \b8_FZFFLXYE[1]\ : SLE
      port map(D => \b12_2_St6KCa_jHv[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b4_2o_z, ALn => b5_voSc3_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b8_FZFFLXYE[1]_net_1\);
    
    \genblk9.b7_nYJ_BFM[89]\ : SLE
      port map(D => \b7_nYJ_BFM[88]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[89]\);
    
    \genblk9.b7_nYJ_BFM[77]\ : SLE
      port map(D => \b7_nYJ_BFM[76]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[77]\);
    
    \genblk9.b7_nYJ_BFM[50]\ : SLE
      port map(D => \b7_nYJ_BFM[49]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[50]\);
    
    \genblk9.b3_PfG[22]\ : SLE
      port map(D => \b3_PfG_6[22]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[22]\);
    
    \genblk9.b3_PfG_RNO[24]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[25]\, C => 
        \b7_vFW_PlM[23]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[24]\);
    
    \genblk9.b3_PfG[137]\ : SLE
      port map(D => \b3_PfG_6[137]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[137]\);
    
    \genblk9.b3_PfG_RNO[98]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[99]\, C => 
        \b7_vFW_PlM[97]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[98]\);
    
    \genblk9.b7_nYJ_BFM[30]\ : SLE
      port map(D => \b7_nYJ_BFM[29]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[30]\);
    
    \genblk9.b7_nYJ_BFM[67]\ : SLE
      port map(D => \b7_nYJ_BFM[66]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[67]\);
    
    \genblk9.b7_nYJ_BFM[159]\ : SLE
      port map(D => \b7_nYJ_BFM[158]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[159]\);
    
    \genblk9.b3_PfG[95]\ : SLE
      port map(D => \b3_PfG_6[95]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[95]\);
    
    \genblk9.b3_PfG[71]\ : SLE
      port map(D => \b3_PfG_6[71]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[71]\);
    
    \genblk9.b3_PfG[1]\ : SLE
      port map(D => \b3_PfG_6[1]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[1]\);
    
    \genblk9.b3_PfG[29]\ : SLE
      port map(D => \b3_PfG_6[29]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[29]\);
    
    \genblk9.b3_PfG_RNO[69]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[70]\, C => 
        \b7_vFW_PlM[68]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[69]\);
    
    \genblk9.b3_PfG[87]\ : SLE
      port map(D => \b3_PfG_6[87]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[87]\);
    
    b7_yYh03wy4_0_a2 : CFG4
      generic map(INIT => x"1000")

      port map(A => IICE_comm2iice(5), B => IICE_comm2iice(4), C
         => IICE_comm2iice(2), D => \b7_yYh03wy4_0_a2_0_2\, Y => 
        b7_yYh03wy4);
    
    \genblk9.b7_nYJ_BFM[102]\ : SLE
      port map(D => \b7_nYJ_BFM[101]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[102]\);
    
    \genblk9.b3_PfG_RNO[49]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[50]\, C => 
        \b7_vFW_PlM[48]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[49]\);
    
    \genblk9.b3_PfG_RNO[35]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[36]\, C => 
        \b7_vFW_PlM[34]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[35]\);
    
    \genblk9.b3_PfG_RNO[52]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[53]\, C => 
        \b7_vFW_PlM[51]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[52]\);
    
    \genblk9.b3_PfG[112]\ : SLE
      port map(D => \b3_PfG_6[112]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[112]\);
    
    \genblk9.b3_PfG_RNO[87]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[88]\, C => 
        \b7_vFW_PlM[86]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[87]\);
    
    \b8_FZFFLXYE[9]\ : SLE
      port map(D => \b12_2_St6KCa_jHv[9]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b4_2o_z, ALn => b5_voSc3_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b8_FZFFLXYE[9]_net_1\);
    
    \b8_FZFFLXYE[5]\ : SLE
      port map(D => \b12_2_St6KCa_jHv[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b4_2o_z, ALn => b5_voSc3_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b8_FZFFLXYE[5]_net_1\);
    
    \genblk9.b3_PfG_RNO[73]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[74]\, C => 
        \b7_vFW_PlM[72]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[73]\);
    
    \genblk9.b3_PfG[61]\ : SLE
      port map(D => \b3_PfG_6[61]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[61]\);
    
    \genblk9.b7_nYJ_BFM[136]\ : SLE
      port map(D => \b7_nYJ_BFM[135]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[136]\);
    
    \genblk9.b9_v_mzCDYXs_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \b9_v_mzCDYXs[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => \b9_v_mzCDYXs_cry[6]\, 
        S => \b9_v_mzCDYXs_s[7]\, Y => OPEN, FCO => 
        \b9_v_mzCDYXs_cry[7]\);
    
    \genblk9.b7_nYJ_BFM[88]\ : SLE
      port map(D => \b7_nYJ_BFM[87]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[88]\);
    
    \genblk9.b3_PfG[30]\ : SLE
      port map(D => \b3_PfG_6[30]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[30]\);
    
    \genblk9.b3_PfG_RNO[146]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[147]\, C => 
        \b7_vFW_PlM[145]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[146]\);
    
    \genblk9.b3_PfG_RNO[64]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[65]\, C => 
        \b7_vFW_PlM[63]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[64]\);
    
    \genblk9.b7_nYJ_BFM[155]\ : SLE
      port map(D => \b7_nYJ_BFM[154]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[155]\);
    
    \genblk9.b7_nYJ_BFM[97]\ : SLE
      port map(D => \b7_nYJ_BFM[96]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[97]\);
    
    \genblk9.b7_nYJ_BFM[42]\ : SLE
      port map(D => \b7_nYJ_BFM[41]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[42]\);
    
    \genblk9.b3_PfG_RNO[44]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[45]\, C => 
        \b7_vFW_PlM[43]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[44]\);
    
    \genblk9.b7_nYJ_BFM[153]\ : SLE
      port map(D => \b7_nYJ_BFM[152]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[153]\);
    
    \genblk9.b3_PfG_RNO[152]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[153]\, C => 
        \b7_vFW_PlM[151]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[152]\);
    
    \b12_2_St6KCa_jHv_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \b12_2_St6KCa_jHv[2]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \b12_2_St6KCa_jHv_cry[1]_net_1\, S => 
        \b12_2_St6KCa_jHv_s[2]\, Y => OPEN, FCO => 
        \b12_2_St6KCa_jHv_cry[2]_net_1\);
    
    \genblk9.b7_nYJ_BFM[15]\ : SLE
      port map(D => \b7_nYJ_BFM[14]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[15]\);
    
    \genblk9.b3_PfG[157]\ : SLE
      port map(D => \b3_PfG_6[157]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[157]\);
    
    \genblk9.b3_PfG_RNO[126]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[127]\, C => 
        \b7_vFW_PlM[125]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[126]\);
    
    \genblk9.b3_PfG[82]\ : SLE
      port map(D => \b3_PfG_6[82]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[82]\);
    
    \genblk9.b7_nYJ_BFM[154]\ : SLE
      port map(D => \b7_nYJ_BFM[153]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[154]\);
    
    \genblk9.b7_nYJ_BFM[26]\ : SLE
      port map(D => \b7_nYJ_BFM[25]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[26]\);
    
    \genblk9.b9_v_mzCDYXs_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \b9_v_mzCDYXs[1]\, C => 
        GND_net_1, D => GND_net_1, FCI => b9_v_mzCDYXs_s_901_FCO, 
        S => \b9_v_mzCDYXs_s[1]\, Y => OPEN, FCO => 
        \b9_v_mzCDYXs_cry[1]\);
    
    \genblk9.b3_PfG[132]\ : SLE
      port map(D => \b3_PfG_6[132]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[132]\);
    
    \genblk9.b3_PfG_6[0]\ : CFG3
      generic map(INIT => x"02")

      port map(A => \b3_PfG[1]\, B => b11_nFG0rDY_9e2, C => 
        \b7_nYJ_BFM[174]\, Y => \b3_PfG_6[0]\);
    
    \genblk9.b3_PfG_RNO[18]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[19]\, C => 
        \b7_vFW_PlM[17]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[18]\);
    
    \genblk9.b3_PfG[23]\ : SLE
      port map(D => \b3_PfG_6[23]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[23]\);
    
    \genblk9.b3_PfG[89]\ : SLE
      port map(D => \b3_PfG_6[89]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[89]\);
    
    \genblk9.b3_PfG[76]\ : SLE
      port map(D => \b3_PfG_6[76]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[76]\);
    
    \genblk9.b3_PfG[45]\ : SLE
      port map(D => \b3_PfG_6[45]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[45]\);
    
    \genblk9.b3_PfG_RNO[158]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[159]\, C => 
        \b7_vFW_PlM[157]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[158]\);
    
    \genblk9.b7_nYJ_BFM[108]\ : SLE
      port map(D => \b7_nYJ_BFM[107]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[108]\);
    
    \genblk9.b3_PfG_RNO[157]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[158]\, C => 
        \b7_vFW_PlM[156]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[157]\);
    
    \genblk9.b3_PfG_RNO[53]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[54]\, C => 
        \b7_vFW_PlM[52]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[53]\);
    
    \genblk9.b3_PfG_RNO[77]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[78]\, C => 
        \b7_vFW_PlM[76]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[77]\);
    
    \genblk9.b3_PfG[66]\ : SLE
      port map(D => \b3_PfG_6[66]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[66]\);
    
    \genblk9.b7_nYJ_BFM[53]\ : SLE
      port map(D => \b7_nYJ_BFM[52]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[53]\);
    
    \genblk9.b7_nYJ_BFM[11]\ : SLE
      port map(D => \b7_nYJ_BFM[10]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[11]\);
    
    b8_jAA_KlCO_0_sqmuxa_8 : CFG4
      generic map(INIT => x"8000")

      port map(A => \b12_2_St6KCa_jHv[7]_net_1\, B => 
        \b12_2_St6KCa_jHv[6]_net_1\, C => 
        \b12_2_St6KCa_jHv[5]_net_1\, D => 
        \b12_2_St6KCa_jHv[4]_net_1\, Y => 
        \b8_jAA_KlCO_0_sqmuxa_8\);
    
    \genblk9.b7_nYJ_BFM[9]\ : SLE
      port map(D => \b7_nYJ_BFM[8]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[9]\);
    
    \b8_FZFFLXYE[10]\ : SLE
      port map(D => \b12_2_St6KCa_jHv[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b4_2o_z, ALn => b5_voSc3_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b8_FZFFLXYE[10]_net_1\);
    
    \b12_2_St6KCa_jHv[2]\ : SLE
      port map(D => \b12_2_St6KCa_jHv_s[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b4_2o_z, ALn => b5_voSc3_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b12_2_St6KCa_jHv[2]_net_1\);
    
    \genblk9.b7_nYJ_BFM[152]\ : SLE
      port map(D => \b7_nYJ_BFM[151]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[152]\);
    
    \genblk9.b3_PfG_RNO[135]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[136]\, C => 
        \b7_vFW_PlM[134]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[135]\);
    
    \b12_2_St6KCa_jHv_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \b12_2_St6KCa_jHv[5]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \b12_2_St6KCa_jHv_cry[4]_net_1\, S => 
        \b12_2_St6KCa_jHv_s[5]\, Y => OPEN, FCO => 
        \b12_2_St6KCa_jHv_cry[5]_net_1\);
    
    \genblk9.b7_nYJ_BFM[33]\ : SLE
      port map(D => \b7_nYJ_BFM[32]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[33]\);
    
    \genblk9.b3_PfG[50]\ : SLE
      port map(D => \b3_PfG_6[50]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[50]\);
    
    \genblk9.b3_PfG_RNO[39]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[40]\, C => 
        \b7_vFW_PlM[38]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[39]\);
    
    \genblk9.b3_PfG_RNO[116]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[117]\, C => 
        \b7_vFW_PlM[115]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[116]\);
    
    \genblk9.b3_PfG[0]\ : SLE
      port map(D => \b3_PfG_6[0]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => b10_OFWNT9_Y2x);
    
    \genblk9.b3_PfG_RNO[21]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[22]\, C => 
        \b7_vFW_PlM[20]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[21]\);
    
    \genblk9.b3_PfG_RNO[20]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[21]\, C => 
        \b7_vFW_PlM[19]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[20]\);
    
    \genblk9.b3_PfG[129]\ : SLE
      port map(D => \b3_PfG_6[129]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[129]\);
    
    \genblk9.b7_nYJ_BFM[49]\ : SLE
      port map(D => \b7_nYJ_BFM[48]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[49]\);
    
    \genblk9.b3_PfG_RNO[105]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[106]\, C => 
        \b7_vFW_PlM[104]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[105]\);
    
    \genblk9.b7_nYJ_BFM[75]\ : SLE
      port map(D => \b7_nYJ_BFM[74]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[75]\);
    
    \genblk9.b3_PfG_RNO[131]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[132]\, C => 
        \b7_vFW_PlM[130]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[131]\);
    
    \genblk9.b3_PfG[152]\ : SLE
      port map(D => \b3_PfG_6[152]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[152]\);
    
    \b12_2_St6KCa_jHv_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \b12_2_St6KCa_jHv[4]_net_1\, 
        C => GND_net_1, D => GND_net_1, FCI => 
        \b12_2_St6KCa_jHv_cry[3]_net_1\, S => 
        \b12_2_St6KCa_jHv_s[4]\, Y => OPEN, FCO => 
        \b12_2_St6KCa_jHv_cry[4]_net_1\);
    
    \genblk9.b3_PfG[111]\ : SLE
      port map(D => \b3_PfG_6[111]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[111]\);
    
    b7_yYh03wy5_0_a2 : CFG4
      generic map(INIT => x"2000")

      port map(A => IICE_comm2iice(5), B => IICE_comm2iice(4), C
         => IICE_comm2iice(2), D => \b7_yYh03wy4_0_a2_0_2\, Y => 
        b7_yYh03wy5);
    
    \genblk9.b3_PfG_RNO[34]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[35]\, C => 
        \b7_vFW_PlM[33]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[34]\);
    
    \genblk9.b7_nYJ_BFM[54]\ : SLE
      port map(D => \b7_nYJ_BFM[53]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[54]\);
    
    \genblk9.b7_nYJ_BFM[65]\ : SLE
      port map(D => \b7_nYJ_BFM[64]\, CLK => IICE_comm2iice(11), 
        EN => \N_15_i\, ALn => b5_voSc3_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b7_nYJ_BFM[65]\);
    
    \genblk9.b3_PfG[109]\ : SLE
      port map(D => \b3_PfG_6[109]\, CLK => IICE_comm2iice(11), 
        EN => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[109]\);
    
    \genblk9.b3_PfG[83]\ : SLE
      port map(D => \b3_PfG_6[83]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[83]\);
    
    \b12_2_St6KCa_jHv[1]\ : SLE
      port map(D => \b12_2_St6KCa_jHv_s[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b4_2o_z, ALn => b5_voSc3_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b12_2_St6KCa_jHv[1]_net_1\);
    
    \genblk9.b3_PfG_RNO[134]\ : CFG4
      generic map(INIT => x"F0E4")

      port map(A => b11_nFG0rDY_9e2, B => \b3_PfG[135]\, C => 
        \b7_vFW_PlM[133]\, D => \b7_nYJ_BFM[174]\, Y => 
        \b3_PfG_6[134]\);
    
    \genblk9.b3_PfG[7]\ : SLE
      port map(D => \b3_PfG_6[7]\, CLK => IICE_comm2iice(11), EN
         => un1_b7_nYJ_BFM8, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b3_PfG[7]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b3_uKr_x is

    port( b13_nvmFL_fx2rbuQ : in    std_logic_vector(6 downto 1);
          b11_uRrc_9urXBb   : in    std_logic;
          b3_PLy            : in    std_logic;
          b3_PLF            : out   std_logic;
          b7_PLy_PlM        : out   std_logic;
          b7_nUTQ_9u        : out   std_logic;
          b7_PSyi_9u        : out   std_logic;
          b9_OFWNT9_ab      : out   std_logic;
          b9_PbTt39_ab      : out   std_logic;
          b9_PKFoLX_ab      : out   std_logic;
          b9_vbTtJX_ab      : out   std_logic;
          b8_ubTt3_YG       : out   std_logic;
          b9_ibScJX_ab      : out   std_logic;
          b7_yYh0_9u        : out   std_logic;
          b8_nUTQ_XlK       : in    std_logic;
          b8_PSyi_XlK       : in    std_logic;
          b10_OFWNT9_Y2x    : in    std_logic;
          b10_PbTt39_Y2x    : in    std_logic;
          b10_PKFoLX_Y2x    : in    std_logic;
          b10_vbTtJX_Y2x    : in    std_logic;
          b9_ubTt3_Mxf      : in    std_logic;
          b10_ibScJX_Y2x    : in    std_logic;
          b8_yYh0_XlK       : in    std_logic
        );

end b3_uKr_x;

architecture DEF_ARCH of b3_uKr_x is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \b3_PLy\, GND_net_1, VCC_net_1, N_29, N_30, N_50, 
        b9_ibScJX_ab_0_a2_0_0, \b9_ibScJX_ab_0_a2_0\, 
        \b9_OFWNT9_ab_0_a2_0_m1_e_2_1\, 
        \b7_PSyi_9u_0_a2_m1_0_a2_0\, \b9_PKFoLX_ab_0_a2_m1_e_0\, 
        \b3_PLF_u_0_a2_0_0\, b3_PLF_u_0_1, \b3_PLF_u_0_N_4L5_1\, 
        b3_PLF_5_i_m2_0_0_y0, b3_PLF_5_i_m2_0_0_co0 : std_logic;

begin 

    \b3_PLy\ <= b3_PLy;
    b7_PLy_PlM <= \b3_PLy\;

    b9_vbTtJX_ab_0_a2 : CFG4
      generic map(INIT => x"2000")

      port map(A => b13_nvmFL_fx2rbuQ(3), B => 
        b13_nvmFL_fx2rbuQ(2), C => b13_nvmFL_fx2rbuQ(1), D => 
        N_50, Y => b9_vbTtJX_ab);
    
    b7_yYh0_9u_0_a2 : CFG4
      generic map(INIT => x"8000")

      port map(A => b13_nvmFL_fx2rbuQ(6), B => 
        b13_nvmFL_fx2rbuQ(5), C => b13_nvmFL_fx2rbuQ(4), D => 
        b11_uRrc_9urXBb, Y => b7_yYh0_9u);
    
    b3_PLF_u_0 : CFG4
      generic map(INIT => x"8A0A")

      port map(A => b11_uRrc_9urXBb, B => \b3_PLF_u_0_a2_0_0\, C
         => b3_PLF_u_0_1, D => b8_yYh0_XlK, Y => b3_PLF);
    
    b9_OFWNT9_ab_0_a2_0_m1_e_2_1 : CFG3
      generic map(INIT => x"04")

      port map(A => b13_nvmFL_fx2rbuQ(4), B => 
        b13_nvmFL_fx2rbuQ(2), C => b13_nvmFL_fx2rbuQ(1), Y => 
        \b9_OFWNT9_ab_0_a2_0_m1_e_2_1\);
    
    b8_ubTt3_YG_0_a2 : CFG4
      generic map(INIT => x"8000")

      port map(A => b9_ibScJX_ab_0_a2_0_0, B => 
        b13_nvmFL_fx2rbuQ(3), C => b11_uRrc_9urXBb, D => 
        \b9_OFWNT9_ab_0_a2_0_m1_e_2_1\, Y => b8_ubTt3_YG);
    
    b7_nUTQ_9u_0_a2 : CFG4
      generic map(INIT => x"0100")

      port map(A => b13_nvmFL_fx2rbuQ(3), B => 
        b13_nvmFL_fx2rbuQ(2), C => b13_nvmFL_fx2rbuQ(1), D => 
        N_50, Y => b7_nUTQ_9u);
    
    b9_OFWNT9_ab_0_a2_m1_e : CFG4
      generic map(INIT => x"2000")

      port map(A => b9_ibScJX_ab_0_a2_0_0, B => 
        b13_nvmFL_fx2rbuQ(3), C => b11_uRrc_9urXBb, D => 
        \b9_OFWNT9_ab_0_a2_0_m1_e_2_1\, Y => b9_OFWNT9_ab);
    
    b9_ibScJX_ab_0_a2_0 : CFG3
      generic map(INIT => x"02")

      port map(A => b13_nvmFL_fx2rbuQ(4), B => 
        b13_nvmFL_fx2rbuQ(3), C => b13_nvmFL_fx2rbuQ(2), Y => 
        \b9_ibScJX_ab_0_a2_0\);
    
    b3_PLF_u_0_N_4L5_1 : CFG3
      generic map(INIT => x"10")

      port map(A => b13_nvmFL_fx2rbuQ(4), B => 
        b13_nvmFL_fx2rbuQ(2), C => N_29, Y => 
        \b3_PLF_u_0_N_4L5_1\);
    
    b3_PLF_u_0_a2_0_0 : CFG3
      generic map(INIT => x"80")

      port map(A => b13_nvmFL_fx2rbuQ(6), B => 
        b13_nvmFL_fx2rbuQ(5), C => b13_nvmFL_fx2rbuQ(4), Y => 
        \b3_PLF_u_0_a2_0_0\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_PLF_2_i_m2 : CFG3
      generic map(INIT => x"B8")

      port map(A => b9_ubTt3_Mxf, B => b13_nvmFL_fx2rbuQ(3), C
         => b10_OFWNT9_Y2x, Y => N_30);
    
    b9_ibScJX_ab_0_a2_0_0_0 : CFG2
      generic map(INIT => x"1")

      port map(A => b13_nvmFL_fx2rbuQ(5), B => 
        b13_nvmFL_fx2rbuQ(6), Y => b9_ibScJX_ab_0_a2_0_0);
    
    b3_PLF_u_0_N_4L5 : CFG4
      generic map(INIT => x"13FF")

      port map(A => \b9_OFWNT9_ab_0_a2_0_m1_e_2_1\, B => 
        \b3_PLF_u_0_N_4L5_1\, C => N_30, D => 
        b9_ibScJX_ab_0_a2_0_0, Y => b3_PLF_u_0_1);
    
    b9_PKFoLX_ab_0_a2_m1_e : CFG4
      generic map(INIT => x"4000")

      port map(A => b13_nvmFL_fx2rbuQ(2), B => 
        b13_nvmFL_fx2rbuQ(3), C => b11_uRrc_9urXBb, D => 
        \b9_PKFoLX_ab_0_a2_m1_e_0\, Y => b9_PKFoLX_ab);
    
    b9_ibScJX_ab_0_a2 : CFG4
      generic map(INIT => x"4000")

      port map(A => b13_nvmFL_fx2rbuQ(1), B => b11_uRrc_9urXBb, C
         => b9_ibScJX_ab_0_a2_0_0, D => \b9_ibScJX_ab_0_a2_0\, Y
         => b9_ibScJX_ab);
    
    b7_PSyi_9u_0_a2_m1_0_a2 : CFG4
      generic map(INIT => x"2000")

      port map(A => b9_ibScJX_ab_0_a2_0_0, B => 
        b13_nvmFL_fx2rbuQ(4), C => b11_uRrc_9urXBb, D => 
        \b7_PSyi_9u_0_a2_m1_0_a2_0\, Y => b7_PSyi_9u);
    
    b9_PbTt39_ab_0_a2 : CFG4
      generic map(INIT => x"4000")

      port map(A => b13_nvmFL_fx2rbuQ(3), B => 
        b13_nvmFL_fx2rbuQ(2), C => b13_nvmFL_fx2rbuQ(1), D => 
        N_50, Y => b9_PbTt39_ab);
    
    b3_PLF_5_i_m2_0_0_wmux_0 : ARI1
      generic map(INIT => x"0F588")

      port map(A => b3_PLF_5_i_m2_0_0_y0, B => 
        b13_nvmFL_fx2rbuQ(3), C => b10_PKFoLX_Y2x, D => 
        b10_vbTtJX_Y2x, FCI => b3_PLF_5_i_m2_0_0_co0, S => OPEN, 
        Y => N_29, FCO => OPEN);
    
    b3_PLF_5_i_m2_0_0_wmux : ARI1
      generic map(INIT => x"0FA44")

      port map(A => b13_nvmFL_fx2rbuQ(1), B => 
        b13_nvmFL_fx2rbuQ(3), C => b8_nUTQ_XlK, D => b8_PSyi_XlK, 
        FCI => VCC_net_1, S => OPEN, Y => b3_PLF_5_i_m2_0_0_y0, 
        FCO => b3_PLF_5_i_m2_0_0_co0);
    
    b7_PSyi_9u_0_a2_m1_0_a2_0 : CFG3
      generic map(INIT => x"10")

      port map(A => b13_nvmFL_fx2rbuQ(3), B => 
        b13_nvmFL_fx2rbuQ(2), C => b13_nvmFL_fx2rbuQ(1), Y => 
        \b7_PSyi_9u_0_a2_m1_0_a2_0\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b9_PKFoLX_ab_0_a2_m1_e_0 : CFG3
      generic map(INIT => x"10")

      port map(A => b13_nvmFL_fx2rbuQ(4), B => 
        b13_nvmFL_fx2rbuQ(1), C => b9_ibScJX_ab_0_a2_0_0, Y => 
        \b9_PKFoLX_ab_0_a2_m1_e_0\);
    
    b3_PLF_u_0_a2_2 : CFG3
      generic map(INIT => x"20")

      port map(A => b11_uRrc_9urXBb, B => b13_nvmFL_fx2rbuQ(4), C
         => b9_ibScJX_ab_0_a2_0_0, Y => N_50);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b5_nvmFL_504s_x_0 is

    port( b4_nUAi          : out   std_logic_vector(502 downto 0);
          IICE_comm2iice_4 : in    std_logic;
          IICE_comm2iice_0 : in    std_logic;
          IICE_comm2iice_3 : in    std_logic;
          b7_PSyi_9u       : in    std_logic;
          b12_PSyi_XlK_qHv : out   std_logic
        );

end b5_nvmFL_504s_x_0;

architecture DEF_ARCH of b5_nvmFL_504s_x_0 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \b4_nUAi[6]\, VCC_net_1, \b4_nUAi[5]\, \b6_OKctIF4\, 
        GND_net_1, \b4_nUAi[4]\, \b4_nUAi[3]\, \b4_nUAi[2]\, 
        \b4_nUAi[1]\, \b4_nUAi[0]\, \b4_nUAi[21]\, \b4_nUAi[20]\, 
        \b4_nUAi[19]\, \b4_nUAi[18]\, \b4_nUAi[17]\, 
        \b4_nUAi[16]\, \b4_nUAi[15]\, \b4_nUAi[14]\, 
        \b4_nUAi[13]\, \b4_nUAi[12]\, \b4_nUAi[11]\, 
        \b4_nUAi[10]\, \b4_nUAi[9]\, \b4_nUAi[8]\, \b4_nUAi[7]\, 
        \b4_nUAi[36]\, \b4_nUAi[35]\, \b4_nUAi[34]\, 
        \b4_nUAi[33]\, \b4_nUAi[32]\, \b4_nUAi[31]\, 
        \b4_nUAi[30]\, \b4_nUAi[29]\, \b4_nUAi[28]\, 
        \b4_nUAi[27]\, \b4_nUAi[26]\, \b4_nUAi[25]\, 
        \b4_nUAi[24]\, \b4_nUAi[23]\, \b4_nUAi[22]\, 
        \b4_nUAi[51]\, \b4_nUAi[50]\, \b4_nUAi[49]\, 
        \b4_nUAi[48]\, \b4_nUAi[47]\, \b4_nUAi[46]\, 
        \b4_nUAi[45]\, \b4_nUAi[44]\, \b4_nUAi[43]\, 
        \b4_nUAi[42]\, \b4_nUAi[41]\, \b4_nUAi[40]\, 
        \b4_nUAi[39]\, \b4_nUAi[38]\, \b4_nUAi[37]\, 
        \b4_nUAi[66]\, \b4_nUAi[65]\, \b4_nUAi[64]\, 
        \b4_nUAi[63]\, \b4_nUAi[62]\, \b4_nUAi[61]\, 
        \b4_nUAi[60]\, \b4_nUAi[59]\, \b4_nUAi[58]\, 
        \b4_nUAi[57]\, \b4_nUAi[56]\, \b4_nUAi[55]\, 
        \b4_nUAi[54]\, \b4_nUAi[53]\, \b4_nUAi[52]\, 
        \b4_nUAi[81]\, \b4_nUAi[80]\, \b4_nUAi[79]\, 
        \b4_nUAi[78]\, \b4_nUAi[77]\, \b4_nUAi[76]\, 
        \b4_nUAi[75]\, \b4_nUAi[74]\, \b4_nUAi[73]\, 
        \b4_nUAi[72]\, \b4_nUAi[71]\, \b4_nUAi[70]\, 
        \b4_nUAi[69]\, \b4_nUAi[68]\, \b4_nUAi[67]\, 
        \b4_nUAi[96]\, \b4_nUAi[95]\, \b4_nUAi[94]\, 
        \b4_nUAi[93]\, \b4_nUAi[92]\, \b4_nUAi[91]\, 
        \b4_nUAi[90]\, \b4_nUAi[89]\, \b4_nUAi[88]\, 
        \b4_nUAi[87]\, \b4_nUAi[86]\, \b4_nUAi[85]\, 
        \b4_nUAi[84]\, \b4_nUAi[83]\, \b4_nUAi[82]\, 
        \b4_nUAi[111]\, \b4_nUAi[110]\, \b4_nUAi[109]\, 
        \b4_nUAi[108]\, \b4_nUAi[107]\, \b4_nUAi[106]\, 
        \b4_nUAi[105]\, \b4_nUAi[104]\, \b4_nUAi[103]\, 
        \b4_nUAi[102]\, \b4_nUAi[101]\, \b4_nUAi[100]\, 
        \b4_nUAi[99]\, \b4_nUAi[98]\, \b4_nUAi[97]\, 
        \b4_nUAi[126]\, \b4_nUAi[125]\, \b4_nUAi[124]\, 
        \b4_nUAi[123]\, \b4_nUAi[122]\, \b4_nUAi[121]\, 
        \b4_nUAi[120]\, \b4_nUAi[119]\, \b4_nUAi[118]\, 
        \b4_nUAi[117]\, \b4_nUAi[116]\, \b4_nUAi[115]\, 
        \b4_nUAi[114]\, \b4_nUAi[113]\, \b4_nUAi[112]\, 
        \b4_nUAi[141]\, \b4_nUAi[140]\, \b4_nUAi[139]\, 
        \b4_nUAi[138]\, \b4_nUAi[137]\, \b4_nUAi[136]\, 
        \b4_nUAi[135]\, \b4_nUAi[134]\, \b4_nUAi[133]\, 
        \b4_nUAi[132]\, \b4_nUAi[131]\, \b4_nUAi[130]\, 
        \b4_nUAi[129]\, \b4_nUAi[128]\, \b4_nUAi[127]\, 
        \b4_nUAi[156]\, \b4_nUAi[155]\, \b4_nUAi[154]\, 
        \b4_nUAi[153]\, \b4_nUAi[152]\, \b4_nUAi[151]\, 
        \b4_nUAi[150]\, \b4_nUAi[149]\, \b4_nUAi[148]\, 
        \b4_nUAi[147]\, \b4_nUAi[146]\, \b4_nUAi[145]\, 
        \b4_nUAi[144]\, \b4_nUAi[143]\, \b4_nUAi[142]\, 
        \b4_nUAi[171]\, \b4_nUAi[170]\, \b4_nUAi[169]\, 
        \b4_nUAi[168]\, \b4_nUAi[167]\, \b4_nUAi[166]\, 
        \b4_nUAi[165]\, \b4_nUAi[164]\, \b4_nUAi[163]\, 
        \b4_nUAi[162]\, \b4_nUAi[161]\, \b4_nUAi[160]\, 
        \b4_nUAi[159]\, \b4_nUAi[158]\, \b4_nUAi[157]\, 
        \b4_nUAi[186]\, \b4_nUAi[185]\, \b4_nUAi[184]\, 
        \b4_nUAi[183]\, \b4_nUAi[182]\, \b4_nUAi[181]\, 
        \b4_nUAi[180]\, \b4_nUAi[179]\, \b4_nUAi[178]\, 
        \b4_nUAi[177]\, \b4_nUAi[176]\, \b4_nUAi[175]\, 
        \b4_nUAi[174]\, \b4_nUAi[173]\, \b4_nUAi[172]\, 
        \b4_nUAi[201]\, \b4_nUAi[200]\, \b4_nUAi[199]\, 
        \b4_nUAi[198]\, \b4_nUAi[197]\, \b4_nUAi[196]\, 
        \b4_nUAi[195]\, \b4_nUAi[194]\, \b4_nUAi[193]\, 
        \b4_nUAi[192]\, \b4_nUAi[191]\, \b4_nUAi[190]\, 
        \b4_nUAi[189]\, \b4_nUAi[188]\, \b4_nUAi[187]\, 
        \b4_nUAi[216]\, \b4_nUAi[215]\, \b4_nUAi[214]\, 
        \b4_nUAi[213]\, \b4_nUAi[212]\, \b4_nUAi[211]\, 
        \b4_nUAi[210]\, \b4_nUAi[209]\, \b4_nUAi[208]\, 
        \b4_nUAi[207]\, \b4_nUAi[206]\, \b4_nUAi[205]\, 
        \b4_nUAi[204]\, \b4_nUAi[203]\, \b4_nUAi[202]\, 
        \b4_nUAi[231]\, \b4_nUAi[230]\, \b4_nUAi[229]\, 
        \b4_nUAi[228]\, \b4_nUAi[227]\, \b4_nUAi[226]\, 
        \b4_nUAi[225]\, \b4_nUAi[224]\, \b4_nUAi[223]\, 
        \b4_nUAi[222]\, \b4_nUAi[221]\, \b4_nUAi[220]\, 
        \b4_nUAi[219]\, \b4_nUAi[218]\, \b4_nUAi[217]\, 
        \b4_nUAi[246]\, \b4_nUAi[245]\, \b4_nUAi[244]\, 
        \b4_nUAi[243]\, \b4_nUAi[242]\, \b4_nUAi[241]\, 
        \b4_nUAi[240]\, \b4_nUAi[239]\, \b4_nUAi[238]\, 
        \b4_nUAi[237]\, \b4_nUAi[236]\, \b4_nUAi[235]\, 
        \b4_nUAi[234]\, \b4_nUAi[233]\, \b4_nUAi[232]\, 
        \b4_nUAi[261]\, \b4_nUAi[260]\, \b4_nUAi[259]\, 
        \b4_nUAi[258]\, \b4_nUAi[257]\, \b4_nUAi[256]\, 
        \b4_nUAi[255]\, \b4_nUAi[254]\, \b4_nUAi[253]\, 
        \b4_nUAi[252]\, \b4_nUAi[251]\, \b4_nUAi[250]\, 
        \b4_nUAi[249]\, \b4_nUAi[248]\, \b4_nUAi[247]\, 
        \b4_nUAi[276]\, \b4_nUAi[275]\, \b4_nUAi[274]\, 
        \b4_nUAi[273]\, \b4_nUAi[272]\, \b4_nUAi[271]\, 
        \b4_nUAi[270]\, \b4_nUAi[269]\, \b4_nUAi[268]\, 
        \b4_nUAi[267]\, \b4_nUAi[266]\, \b4_nUAi[265]\, 
        \b4_nUAi[264]\, \b4_nUAi[263]\, \b4_nUAi[262]\, 
        \b4_nUAi[291]\, \b4_nUAi[290]\, \b4_nUAi[289]\, 
        \b4_nUAi[288]\, \b4_nUAi[287]\, \b4_nUAi[286]\, 
        \b4_nUAi[285]\, \b4_nUAi[284]\, \b4_nUAi[283]\, 
        \b4_nUAi[282]\, \b4_nUAi[281]\, \b4_nUAi[280]\, 
        \b4_nUAi[279]\, \b4_nUAi[278]\, \b4_nUAi[277]\, 
        \b4_nUAi[306]\, \b4_nUAi[305]\, \b4_nUAi[304]\, 
        \b4_nUAi[303]\, \b4_nUAi[302]\, \b4_nUAi[301]\, 
        \b4_nUAi[300]\, \b4_nUAi[299]\, \b4_nUAi[298]\, 
        \b4_nUAi[297]\, \b4_nUAi[296]\, \b4_nUAi[295]\, 
        \b4_nUAi[294]\, \b4_nUAi[293]\, \b4_nUAi[292]\, 
        \b4_nUAi[321]\, \b4_nUAi[320]\, \b4_nUAi[319]\, 
        \b4_nUAi[318]\, \b4_nUAi[317]\, \b4_nUAi[316]\, 
        \b4_nUAi[315]\, \b4_nUAi[314]\, \b4_nUAi[313]\, 
        \b4_nUAi[312]\, \b4_nUAi[311]\, \b4_nUAi[310]\, 
        \b4_nUAi[309]\, \b4_nUAi[308]\, \b4_nUAi[307]\, 
        \b4_nUAi[336]\, \b4_nUAi[335]\, \b4_nUAi[334]\, 
        \b4_nUAi[333]\, \b4_nUAi[332]\, \b4_nUAi[331]\, 
        \b4_nUAi[330]\, \b4_nUAi[329]\, \b4_nUAi[328]\, 
        \b4_nUAi[327]\, \b4_nUAi[326]\, \b4_nUAi[325]\, 
        \b4_nUAi[324]\, \b4_nUAi[323]\, \b4_nUAi[322]\, 
        \b4_nUAi[351]\, \b4_nUAi[350]\, \b4_nUAi[349]\, 
        \b4_nUAi[348]\, \b4_nUAi[347]\, \b4_nUAi[346]\, 
        \b4_nUAi[345]\, \b4_nUAi[344]\, \b4_nUAi[343]\, 
        \b4_nUAi[342]\, \b4_nUAi[341]\, \b4_nUAi[340]\, 
        \b4_nUAi[339]\, \b4_nUAi[338]\, \b4_nUAi[337]\, 
        \b4_nUAi[366]\, \b4_nUAi[365]\, \b4_nUAi[364]\, 
        \b4_nUAi[363]\, \b4_nUAi[362]\, \b4_nUAi[361]\, 
        \b4_nUAi[360]\, \b4_nUAi[359]\, \b4_nUAi[358]\, 
        \b4_nUAi[357]\, \b4_nUAi[356]\, \b4_nUAi[355]\, 
        \b4_nUAi[354]\, \b4_nUAi[353]\, \b4_nUAi[352]\, 
        \b4_nUAi[381]\, \b4_nUAi[380]\, \b4_nUAi[379]\, 
        \b4_nUAi[378]\, \b4_nUAi[377]\, \b4_nUAi[376]\, 
        \b4_nUAi[375]\, \b4_nUAi[374]\, \b4_nUAi[373]\, 
        \b4_nUAi[372]\, \b4_nUAi[371]\, \b4_nUAi[370]\, 
        \b4_nUAi[369]\, \b4_nUAi[368]\, \b4_nUAi[367]\, 
        \b4_nUAi[396]\, \b4_nUAi[395]\, \b4_nUAi[394]\, 
        \b4_nUAi[393]\, \b4_nUAi[392]\, \b4_nUAi[391]\, 
        \b4_nUAi[390]\, \b4_nUAi[389]\, \b4_nUAi[388]\, 
        \b4_nUAi[387]\, \b4_nUAi[386]\, \b4_nUAi[385]\, 
        \b4_nUAi[384]\, \b4_nUAi[383]\, \b4_nUAi[382]\, 
        \b4_nUAi[411]\, \b4_nUAi[410]\, \b4_nUAi[409]\, 
        \b4_nUAi[408]\, \b4_nUAi[407]\, \b4_nUAi[406]\, 
        \b4_nUAi[405]\, \b4_nUAi[404]\, \b4_nUAi[403]\, 
        \b4_nUAi[402]\, \b4_nUAi[401]\, \b4_nUAi[400]\, 
        \b4_nUAi[399]\, \b4_nUAi[398]\, \b4_nUAi[397]\, 
        \b4_nUAi[426]\, \b4_nUAi[425]\, \b4_nUAi[424]\, 
        \b4_nUAi[423]\, \b4_nUAi[422]\, \b4_nUAi[421]\, 
        \b4_nUAi[420]\, \b4_nUAi[419]\, \b4_nUAi[418]\, 
        \b4_nUAi[417]\, \b4_nUAi[416]\, \b4_nUAi[415]\, 
        \b4_nUAi[414]\, \b4_nUAi[413]\, \b4_nUAi[412]\, 
        \b4_nUAi[441]\, \b4_nUAi[440]\, \b4_nUAi[439]\, 
        \b4_nUAi[438]\, \b4_nUAi[437]\, \b4_nUAi[436]\, 
        \b4_nUAi[435]\, \b4_nUAi[434]\, \b4_nUAi[433]\, 
        \b4_nUAi[432]\, \b4_nUAi[431]\, \b4_nUAi[430]\, 
        \b4_nUAi[429]\, \b4_nUAi[428]\, \b4_nUAi[427]\, 
        \b4_nUAi[456]\, \b4_nUAi[455]\, \b4_nUAi[454]\, 
        \b4_nUAi[453]\, \b4_nUAi[452]\, \b4_nUAi[451]\, 
        \b4_nUAi[450]\, \b4_nUAi[449]\, \b4_nUAi[448]\, 
        \b4_nUAi[447]\, \b4_nUAi[446]\, \b4_nUAi[445]\, 
        \b4_nUAi[444]\, \b4_nUAi[443]\, \b4_nUAi[442]\, 
        \b4_nUAi[471]\, \b4_nUAi[470]\, \b4_nUAi[469]\, 
        \b4_nUAi[468]\, \b4_nUAi[467]\, \b4_nUAi[466]\, 
        \b4_nUAi[465]\, \b4_nUAi[464]\, \b4_nUAi[463]\, 
        \b4_nUAi[462]\, \b4_nUAi[461]\, \b4_nUAi[460]\, 
        \b4_nUAi[459]\, \b4_nUAi[458]\, \b4_nUAi[457]\, 
        \b4_nUAi[486]\, \b4_nUAi[485]\, \b4_nUAi[484]\, 
        \b4_nUAi[483]\, \b4_nUAi[482]\, \b4_nUAi[481]\, 
        \b4_nUAi[480]\, \b4_nUAi[479]\, \b4_nUAi[478]\, 
        \b4_nUAi[477]\, \b4_nUAi[476]\, \b4_nUAi[475]\, 
        \b4_nUAi[474]\, \b4_nUAi[473]\, \b4_nUAi[472]\, 
        \b4_nUAi[501]\, \b4_nUAi[500]\, \b4_nUAi[499]\, 
        \b4_nUAi[498]\, \b4_nUAi[497]\, \b4_nUAi[496]\, 
        \b4_nUAi[495]\, \b4_nUAi[494]\, \b4_nUAi[493]\, 
        \b4_nUAi[492]\, \b4_nUAi[491]\, \b4_nUAi[490]\, 
        \b4_nUAi[489]\, \b4_nUAi[488]\, \b4_nUAi[487]\, 
        \b4_nUAi[502]\ : std_logic;

begin 

    b4_nUAi(502) <= \b4_nUAi[502]\;
    b4_nUAi(501) <= \b4_nUAi[501]\;
    b4_nUAi(500) <= \b4_nUAi[500]\;
    b4_nUAi(499) <= \b4_nUAi[499]\;
    b4_nUAi(498) <= \b4_nUAi[498]\;
    b4_nUAi(497) <= \b4_nUAi[497]\;
    b4_nUAi(496) <= \b4_nUAi[496]\;
    b4_nUAi(495) <= \b4_nUAi[495]\;
    b4_nUAi(494) <= \b4_nUAi[494]\;
    b4_nUAi(493) <= \b4_nUAi[493]\;
    b4_nUAi(492) <= \b4_nUAi[492]\;
    b4_nUAi(491) <= \b4_nUAi[491]\;
    b4_nUAi(490) <= \b4_nUAi[490]\;
    b4_nUAi(489) <= \b4_nUAi[489]\;
    b4_nUAi(488) <= \b4_nUAi[488]\;
    b4_nUAi(487) <= \b4_nUAi[487]\;
    b4_nUAi(486) <= \b4_nUAi[486]\;
    b4_nUAi(485) <= \b4_nUAi[485]\;
    b4_nUAi(484) <= \b4_nUAi[484]\;
    b4_nUAi(483) <= \b4_nUAi[483]\;
    b4_nUAi(482) <= \b4_nUAi[482]\;
    b4_nUAi(481) <= \b4_nUAi[481]\;
    b4_nUAi(480) <= \b4_nUAi[480]\;
    b4_nUAi(479) <= \b4_nUAi[479]\;
    b4_nUAi(478) <= \b4_nUAi[478]\;
    b4_nUAi(477) <= \b4_nUAi[477]\;
    b4_nUAi(476) <= \b4_nUAi[476]\;
    b4_nUAi(475) <= \b4_nUAi[475]\;
    b4_nUAi(474) <= \b4_nUAi[474]\;
    b4_nUAi(473) <= \b4_nUAi[473]\;
    b4_nUAi(472) <= \b4_nUAi[472]\;
    b4_nUAi(471) <= \b4_nUAi[471]\;
    b4_nUAi(470) <= \b4_nUAi[470]\;
    b4_nUAi(469) <= \b4_nUAi[469]\;
    b4_nUAi(468) <= \b4_nUAi[468]\;
    b4_nUAi(467) <= \b4_nUAi[467]\;
    b4_nUAi(466) <= \b4_nUAi[466]\;
    b4_nUAi(465) <= \b4_nUAi[465]\;
    b4_nUAi(464) <= \b4_nUAi[464]\;
    b4_nUAi(463) <= \b4_nUAi[463]\;
    b4_nUAi(462) <= \b4_nUAi[462]\;
    b4_nUAi(461) <= \b4_nUAi[461]\;
    b4_nUAi(460) <= \b4_nUAi[460]\;
    b4_nUAi(459) <= \b4_nUAi[459]\;
    b4_nUAi(458) <= \b4_nUAi[458]\;
    b4_nUAi(457) <= \b4_nUAi[457]\;
    b4_nUAi(456) <= \b4_nUAi[456]\;
    b4_nUAi(455) <= \b4_nUAi[455]\;
    b4_nUAi(454) <= \b4_nUAi[454]\;
    b4_nUAi(453) <= \b4_nUAi[453]\;
    b4_nUAi(452) <= \b4_nUAi[452]\;
    b4_nUAi(451) <= \b4_nUAi[451]\;
    b4_nUAi(450) <= \b4_nUAi[450]\;
    b4_nUAi(449) <= \b4_nUAi[449]\;
    b4_nUAi(448) <= \b4_nUAi[448]\;
    b4_nUAi(447) <= \b4_nUAi[447]\;
    b4_nUAi(446) <= \b4_nUAi[446]\;
    b4_nUAi(445) <= \b4_nUAi[445]\;
    b4_nUAi(444) <= \b4_nUAi[444]\;
    b4_nUAi(443) <= \b4_nUAi[443]\;
    b4_nUAi(442) <= \b4_nUAi[442]\;
    b4_nUAi(441) <= \b4_nUAi[441]\;
    b4_nUAi(440) <= \b4_nUAi[440]\;
    b4_nUAi(439) <= \b4_nUAi[439]\;
    b4_nUAi(438) <= \b4_nUAi[438]\;
    b4_nUAi(437) <= \b4_nUAi[437]\;
    b4_nUAi(436) <= \b4_nUAi[436]\;
    b4_nUAi(435) <= \b4_nUAi[435]\;
    b4_nUAi(434) <= \b4_nUAi[434]\;
    b4_nUAi(433) <= \b4_nUAi[433]\;
    b4_nUAi(432) <= \b4_nUAi[432]\;
    b4_nUAi(431) <= \b4_nUAi[431]\;
    b4_nUAi(430) <= \b4_nUAi[430]\;
    b4_nUAi(429) <= \b4_nUAi[429]\;
    b4_nUAi(428) <= \b4_nUAi[428]\;
    b4_nUAi(427) <= \b4_nUAi[427]\;
    b4_nUAi(426) <= \b4_nUAi[426]\;
    b4_nUAi(425) <= \b4_nUAi[425]\;
    b4_nUAi(424) <= \b4_nUAi[424]\;
    b4_nUAi(423) <= \b4_nUAi[423]\;
    b4_nUAi(422) <= \b4_nUAi[422]\;
    b4_nUAi(421) <= \b4_nUAi[421]\;
    b4_nUAi(420) <= \b4_nUAi[420]\;
    b4_nUAi(419) <= \b4_nUAi[419]\;
    b4_nUAi(418) <= \b4_nUAi[418]\;
    b4_nUAi(417) <= \b4_nUAi[417]\;
    b4_nUAi(416) <= \b4_nUAi[416]\;
    b4_nUAi(415) <= \b4_nUAi[415]\;
    b4_nUAi(414) <= \b4_nUAi[414]\;
    b4_nUAi(413) <= \b4_nUAi[413]\;
    b4_nUAi(412) <= \b4_nUAi[412]\;
    b4_nUAi(411) <= \b4_nUAi[411]\;
    b4_nUAi(410) <= \b4_nUAi[410]\;
    b4_nUAi(409) <= \b4_nUAi[409]\;
    b4_nUAi(408) <= \b4_nUAi[408]\;
    b4_nUAi(407) <= \b4_nUAi[407]\;
    b4_nUAi(406) <= \b4_nUAi[406]\;
    b4_nUAi(405) <= \b4_nUAi[405]\;
    b4_nUAi(404) <= \b4_nUAi[404]\;
    b4_nUAi(403) <= \b4_nUAi[403]\;
    b4_nUAi(402) <= \b4_nUAi[402]\;
    b4_nUAi(401) <= \b4_nUAi[401]\;
    b4_nUAi(400) <= \b4_nUAi[400]\;
    b4_nUAi(399) <= \b4_nUAi[399]\;
    b4_nUAi(398) <= \b4_nUAi[398]\;
    b4_nUAi(397) <= \b4_nUAi[397]\;
    b4_nUAi(396) <= \b4_nUAi[396]\;
    b4_nUAi(395) <= \b4_nUAi[395]\;
    b4_nUAi(394) <= \b4_nUAi[394]\;
    b4_nUAi(393) <= \b4_nUAi[393]\;
    b4_nUAi(392) <= \b4_nUAi[392]\;
    b4_nUAi(391) <= \b4_nUAi[391]\;
    b4_nUAi(390) <= \b4_nUAi[390]\;
    b4_nUAi(389) <= \b4_nUAi[389]\;
    b4_nUAi(388) <= \b4_nUAi[388]\;
    b4_nUAi(387) <= \b4_nUAi[387]\;
    b4_nUAi(386) <= \b4_nUAi[386]\;
    b4_nUAi(385) <= \b4_nUAi[385]\;
    b4_nUAi(384) <= \b4_nUAi[384]\;
    b4_nUAi(383) <= \b4_nUAi[383]\;
    b4_nUAi(382) <= \b4_nUAi[382]\;
    b4_nUAi(381) <= \b4_nUAi[381]\;
    b4_nUAi(380) <= \b4_nUAi[380]\;
    b4_nUAi(379) <= \b4_nUAi[379]\;
    b4_nUAi(378) <= \b4_nUAi[378]\;
    b4_nUAi(377) <= \b4_nUAi[377]\;
    b4_nUAi(376) <= \b4_nUAi[376]\;
    b4_nUAi(375) <= \b4_nUAi[375]\;
    b4_nUAi(374) <= \b4_nUAi[374]\;
    b4_nUAi(373) <= \b4_nUAi[373]\;
    b4_nUAi(372) <= \b4_nUAi[372]\;
    b4_nUAi(371) <= \b4_nUAi[371]\;
    b4_nUAi(370) <= \b4_nUAi[370]\;
    b4_nUAi(369) <= \b4_nUAi[369]\;
    b4_nUAi(368) <= \b4_nUAi[368]\;
    b4_nUAi(367) <= \b4_nUAi[367]\;
    b4_nUAi(366) <= \b4_nUAi[366]\;
    b4_nUAi(365) <= \b4_nUAi[365]\;
    b4_nUAi(364) <= \b4_nUAi[364]\;
    b4_nUAi(363) <= \b4_nUAi[363]\;
    b4_nUAi(362) <= \b4_nUAi[362]\;
    b4_nUAi(361) <= \b4_nUAi[361]\;
    b4_nUAi(360) <= \b4_nUAi[360]\;
    b4_nUAi(359) <= \b4_nUAi[359]\;
    b4_nUAi(358) <= \b4_nUAi[358]\;
    b4_nUAi(357) <= \b4_nUAi[357]\;
    b4_nUAi(356) <= \b4_nUAi[356]\;
    b4_nUAi(355) <= \b4_nUAi[355]\;
    b4_nUAi(354) <= \b4_nUAi[354]\;
    b4_nUAi(353) <= \b4_nUAi[353]\;
    b4_nUAi(352) <= \b4_nUAi[352]\;
    b4_nUAi(351) <= \b4_nUAi[351]\;
    b4_nUAi(350) <= \b4_nUAi[350]\;
    b4_nUAi(349) <= \b4_nUAi[349]\;
    b4_nUAi(348) <= \b4_nUAi[348]\;
    b4_nUAi(347) <= \b4_nUAi[347]\;
    b4_nUAi(346) <= \b4_nUAi[346]\;
    b4_nUAi(345) <= \b4_nUAi[345]\;
    b4_nUAi(344) <= \b4_nUAi[344]\;
    b4_nUAi(343) <= \b4_nUAi[343]\;
    b4_nUAi(342) <= \b4_nUAi[342]\;
    b4_nUAi(341) <= \b4_nUAi[341]\;
    b4_nUAi(340) <= \b4_nUAi[340]\;
    b4_nUAi(339) <= \b4_nUAi[339]\;
    b4_nUAi(338) <= \b4_nUAi[338]\;
    b4_nUAi(337) <= \b4_nUAi[337]\;
    b4_nUAi(336) <= \b4_nUAi[336]\;
    b4_nUAi(335) <= \b4_nUAi[335]\;
    b4_nUAi(334) <= \b4_nUAi[334]\;
    b4_nUAi(333) <= \b4_nUAi[333]\;
    b4_nUAi(332) <= \b4_nUAi[332]\;
    b4_nUAi(331) <= \b4_nUAi[331]\;
    b4_nUAi(330) <= \b4_nUAi[330]\;
    b4_nUAi(329) <= \b4_nUAi[329]\;
    b4_nUAi(328) <= \b4_nUAi[328]\;
    b4_nUAi(327) <= \b4_nUAi[327]\;
    b4_nUAi(326) <= \b4_nUAi[326]\;
    b4_nUAi(325) <= \b4_nUAi[325]\;
    b4_nUAi(324) <= \b4_nUAi[324]\;
    b4_nUAi(323) <= \b4_nUAi[323]\;
    b4_nUAi(322) <= \b4_nUAi[322]\;
    b4_nUAi(321) <= \b4_nUAi[321]\;
    b4_nUAi(320) <= \b4_nUAi[320]\;
    b4_nUAi(319) <= \b4_nUAi[319]\;
    b4_nUAi(318) <= \b4_nUAi[318]\;
    b4_nUAi(317) <= \b4_nUAi[317]\;
    b4_nUAi(316) <= \b4_nUAi[316]\;
    b4_nUAi(315) <= \b4_nUAi[315]\;
    b4_nUAi(314) <= \b4_nUAi[314]\;
    b4_nUAi(313) <= \b4_nUAi[313]\;
    b4_nUAi(312) <= \b4_nUAi[312]\;
    b4_nUAi(311) <= \b4_nUAi[311]\;
    b4_nUAi(310) <= \b4_nUAi[310]\;
    b4_nUAi(309) <= \b4_nUAi[309]\;
    b4_nUAi(308) <= \b4_nUAi[308]\;
    b4_nUAi(307) <= \b4_nUAi[307]\;
    b4_nUAi(306) <= \b4_nUAi[306]\;
    b4_nUAi(305) <= \b4_nUAi[305]\;
    b4_nUAi(304) <= \b4_nUAi[304]\;
    b4_nUAi(303) <= \b4_nUAi[303]\;
    b4_nUAi(302) <= \b4_nUAi[302]\;
    b4_nUAi(301) <= \b4_nUAi[301]\;
    b4_nUAi(300) <= \b4_nUAi[300]\;
    b4_nUAi(299) <= \b4_nUAi[299]\;
    b4_nUAi(298) <= \b4_nUAi[298]\;
    b4_nUAi(297) <= \b4_nUAi[297]\;
    b4_nUAi(296) <= \b4_nUAi[296]\;
    b4_nUAi(295) <= \b4_nUAi[295]\;
    b4_nUAi(294) <= \b4_nUAi[294]\;
    b4_nUAi(293) <= \b4_nUAi[293]\;
    b4_nUAi(292) <= \b4_nUAi[292]\;
    b4_nUAi(291) <= \b4_nUAi[291]\;
    b4_nUAi(290) <= \b4_nUAi[290]\;
    b4_nUAi(289) <= \b4_nUAi[289]\;
    b4_nUAi(288) <= \b4_nUAi[288]\;
    b4_nUAi(287) <= \b4_nUAi[287]\;
    b4_nUAi(286) <= \b4_nUAi[286]\;
    b4_nUAi(285) <= \b4_nUAi[285]\;
    b4_nUAi(284) <= \b4_nUAi[284]\;
    b4_nUAi(283) <= \b4_nUAi[283]\;
    b4_nUAi(282) <= \b4_nUAi[282]\;
    b4_nUAi(281) <= \b4_nUAi[281]\;
    b4_nUAi(280) <= \b4_nUAi[280]\;
    b4_nUAi(279) <= \b4_nUAi[279]\;
    b4_nUAi(278) <= \b4_nUAi[278]\;
    b4_nUAi(277) <= \b4_nUAi[277]\;
    b4_nUAi(276) <= \b4_nUAi[276]\;
    b4_nUAi(275) <= \b4_nUAi[275]\;
    b4_nUAi(274) <= \b4_nUAi[274]\;
    b4_nUAi(273) <= \b4_nUAi[273]\;
    b4_nUAi(272) <= \b4_nUAi[272]\;
    b4_nUAi(271) <= \b4_nUAi[271]\;
    b4_nUAi(270) <= \b4_nUAi[270]\;
    b4_nUAi(269) <= \b4_nUAi[269]\;
    b4_nUAi(268) <= \b4_nUAi[268]\;
    b4_nUAi(267) <= \b4_nUAi[267]\;
    b4_nUAi(266) <= \b4_nUAi[266]\;
    b4_nUAi(265) <= \b4_nUAi[265]\;
    b4_nUAi(264) <= \b4_nUAi[264]\;
    b4_nUAi(263) <= \b4_nUAi[263]\;
    b4_nUAi(262) <= \b4_nUAi[262]\;
    b4_nUAi(261) <= \b4_nUAi[261]\;
    b4_nUAi(260) <= \b4_nUAi[260]\;
    b4_nUAi(259) <= \b4_nUAi[259]\;
    b4_nUAi(258) <= \b4_nUAi[258]\;
    b4_nUAi(257) <= \b4_nUAi[257]\;
    b4_nUAi(256) <= \b4_nUAi[256]\;
    b4_nUAi(255) <= \b4_nUAi[255]\;
    b4_nUAi(254) <= \b4_nUAi[254]\;
    b4_nUAi(253) <= \b4_nUAi[253]\;
    b4_nUAi(252) <= \b4_nUAi[252]\;
    b4_nUAi(251) <= \b4_nUAi[251]\;
    b4_nUAi(250) <= \b4_nUAi[250]\;
    b4_nUAi(249) <= \b4_nUAi[249]\;
    b4_nUAi(248) <= \b4_nUAi[248]\;
    b4_nUAi(247) <= \b4_nUAi[247]\;
    b4_nUAi(246) <= \b4_nUAi[246]\;
    b4_nUAi(245) <= \b4_nUAi[245]\;
    b4_nUAi(244) <= \b4_nUAi[244]\;
    b4_nUAi(243) <= \b4_nUAi[243]\;
    b4_nUAi(242) <= \b4_nUAi[242]\;
    b4_nUAi(241) <= \b4_nUAi[241]\;
    b4_nUAi(240) <= \b4_nUAi[240]\;
    b4_nUAi(239) <= \b4_nUAi[239]\;
    b4_nUAi(238) <= \b4_nUAi[238]\;
    b4_nUAi(237) <= \b4_nUAi[237]\;
    b4_nUAi(236) <= \b4_nUAi[236]\;
    b4_nUAi(235) <= \b4_nUAi[235]\;
    b4_nUAi(234) <= \b4_nUAi[234]\;
    b4_nUAi(233) <= \b4_nUAi[233]\;
    b4_nUAi(232) <= \b4_nUAi[232]\;
    b4_nUAi(231) <= \b4_nUAi[231]\;
    b4_nUAi(230) <= \b4_nUAi[230]\;
    b4_nUAi(229) <= \b4_nUAi[229]\;
    b4_nUAi(228) <= \b4_nUAi[228]\;
    b4_nUAi(227) <= \b4_nUAi[227]\;
    b4_nUAi(226) <= \b4_nUAi[226]\;
    b4_nUAi(225) <= \b4_nUAi[225]\;
    b4_nUAi(224) <= \b4_nUAi[224]\;
    b4_nUAi(223) <= \b4_nUAi[223]\;
    b4_nUAi(222) <= \b4_nUAi[222]\;
    b4_nUAi(221) <= \b4_nUAi[221]\;
    b4_nUAi(220) <= \b4_nUAi[220]\;
    b4_nUAi(219) <= \b4_nUAi[219]\;
    b4_nUAi(218) <= \b4_nUAi[218]\;
    b4_nUAi(217) <= \b4_nUAi[217]\;
    b4_nUAi(216) <= \b4_nUAi[216]\;
    b4_nUAi(215) <= \b4_nUAi[215]\;
    b4_nUAi(214) <= \b4_nUAi[214]\;
    b4_nUAi(213) <= \b4_nUAi[213]\;
    b4_nUAi(212) <= \b4_nUAi[212]\;
    b4_nUAi(211) <= \b4_nUAi[211]\;
    b4_nUAi(210) <= \b4_nUAi[210]\;
    b4_nUAi(209) <= \b4_nUAi[209]\;
    b4_nUAi(208) <= \b4_nUAi[208]\;
    b4_nUAi(207) <= \b4_nUAi[207]\;
    b4_nUAi(206) <= \b4_nUAi[206]\;
    b4_nUAi(205) <= \b4_nUAi[205]\;
    b4_nUAi(204) <= \b4_nUAi[204]\;
    b4_nUAi(203) <= \b4_nUAi[203]\;
    b4_nUAi(202) <= \b4_nUAi[202]\;
    b4_nUAi(201) <= \b4_nUAi[201]\;
    b4_nUAi(200) <= \b4_nUAi[200]\;
    b4_nUAi(199) <= \b4_nUAi[199]\;
    b4_nUAi(198) <= \b4_nUAi[198]\;
    b4_nUAi(197) <= \b4_nUAi[197]\;
    b4_nUAi(196) <= \b4_nUAi[196]\;
    b4_nUAi(195) <= \b4_nUAi[195]\;
    b4_nUAi(194) <= \b4_nUAi[194]\;
    b4_nUAi(193) <= \b4_nUAi[193]\;
    b4_nUAi(192) <= \b4_nUAi[192]\;
    b4_nUAi(191) <= \b4_nUAi[191]\;
    b4_nUAi(190) <= \b4_nUAi[190]\;
    b4_nUAi(189) <= \b4_nUAi[189]\;
    b4_nUAi(188) <= \b4_nUAi[188]\;
    b4_nUAi(187) <= \b4_nUAi[187]\;
    b4_nUAi(186) <= \b4_nUAi[186]\;
    b4_nUAi(185) <= \b4_nUAi[185]\;
    b4_nUAi(184) <= \b4_nUAi[184]\;
    b4_nUAi(183) <= \b4_nUAi[183]\;
    b4_nUAi(182) <= \b4_nUAi[182]\;
    b4_nUAi(181) <= \b4_nUAi[181]\;
    b4_nUAi(180) <= \b4_nUAi[180]\;
    b4_nUAi(179) <= \b4_nUAi[179]\;
    b4_nUAi(178) <= \b4_nUAi[178]\;
    b4_nUAi(177) <= \b4_nUAi[177]\;
    b4_nUAi(176) <= \b4_nUAi[176]\;
    b4_nUAi(175) <= \b4_nUAi[175]\;
    b4_nUAi(174) <= \b4_nUAi[174]\;
    b4_nUAi(173) <= \b4_nUAi[173]\;
    b4_nUAi(172) <= \b4_nUAi[172]\;
    b4_nUAi(171) <= \b4_nUAi[171]\;
    b4_nUAi(170) <= \b4_nUAi[170]\;
    b4_nUAi(169) <= \b4_nUAi[169]\;
    b4_nUAi(168) <= \b4_nUAi[168]\;
    b4_nUAi(167) <= \b4_nUAi[167]\;
    b4_nUAi(166) <= \b4_nUAi[166]\;
    b4_nUAi(165) <= \b4_nUAi[165]\;
    b4_nUAi(164) <= \b4_nUAi[164]\;
    b4_nUAi(163) <= \b4_nUAi[163]\;
    b4_nUAi(162) <= \b4_nUAi[162]\;
    b4_nUAi(161) <= \b4_nUAi[161]\;
    b4_nUAi(160) <= \b4_nUAi[160]\;
    b4_nUAi(159) <= \b4_nUAi[159]\;
    b4_nUAi(158) <= \b4_nUAi[158]\;
    b4_nUAi(157) <= \b4_nUAi[157]\;
    b4_nUAi(156) <= \b4_nUAi[156]\;
    b4_nUAi(155) <= \b4_nUAi[155]\;
    b4_nUAi(154) <= \b4_nUAi[154]\;
    b4_nUAi(153) <= \b4_nUAi[153]\;
    b4_nUAi(152) <= \b4_nUAi[152]\;
    b4_nUAi(151) <= \b4_nUAi[151]\;
    b4_nUAi(150) <= \b4_nUAi[150]\;
    b4_nUAi(149) <= \b4_nUAi[149]\;
    b4_nUAi(148) <= \b4_nUAi[148]\;
    b4_nUAi(147) <= \b4_nUAi[147]\;
    b4_nUAi(146) <= \b4_nUAi[146]\;
    b4_nUAi(145) <= \b4_nUAi[145]\;
    b4_nUAi(144) <= \b4_nUAi[144]\;
    b4_nUAi(143) <= \b4_nUAi[143]\;
    b4_nUAi(142) <= \b4_nUAi[142]\;
    b4_nUAi(141) <= \b4_nUAi[141]\;
    b4_nUAi(140) <= \b4_nUAi[140]\;
    b4_nUAi(139) <= \b4_nUAi[139]\;
    b4_nUAi(138) <= \b4_nUAi[138]\;
    b4_nUAi(137) <= \b4_nUAi[137]\;
    b4_nUAi(136) <= \b4_nUAi[136]\;
    b4_nUAi(135) <= \b4_nUAi[135]\;
    b4_nUAi(134) <= \b4_nUAi[134]\;
    b4_nUAi(133) <= \b4_nUAi[133]\;
    b4_nUAi(132) <= \b4_nUAi[132]\;
    b4_nUAi(131) <= \b4_nUAi[131]\;
    b4_nUAi(130) <= \b4_nUAi[130]\;
    b4_nUAi(129) <= \b4_nUAi[129]\;
    b4_nUAi(128) <= \b4_nUAi[128]\;
    b4_nUAi(127) <= \b4_nUAi[127]\;
    b4_nUAi(126) <= \b4_nUAi[126]\;
    b4_nUAi(125) <= \b4_nUAi[125]\;
    b4_nUAi(124) <= \b4_nUAi[124]\;
    b4_nUAi(123) <= \b4_nUAi[123]\;
    b4_nUAi(122) <= \b4_nUAi[122]\;
    b4_nUAi(121) <= \b4_nUAi[121]\;
    b4_nUAi(120) <= \b4_nUAi[120]\;
    b4_nUAi(119) <= \b4_nUAi[119]\;
    b4_nUAi(118) <= \b4_nUAi[118]\;
    b4_nUAi(117) <= \b4_nUAi[117]\;
    b4_nUAi(116) <= \b4_nUAi[116]\;
    b4_nUAi(115) <= \b4_nUAi[115]\;
    b4_nUAi(114) <= \b4_nUAi[114]\;
    b4_nUAi(113) <= \b4_nUAi[113]\;
    b4_nUAi(112) <= \b4_nUAi[112]\;
    b4_nUAi(111) <= \b4_nUAi[111]\;
    b4_nUAi(110) <= \b4_nUAi[110]\;
    b4_nUAi(109) <= \b4_nUAi[109]\;
    b4_nUAi(108) <= \b4_nUAi[108]\;
    b4_nUAi(107) <= \b4_nUAi[107]\;
    b4_nUAi(106) <= \b4_nUAi[106]\;
    b4_nUAi(105) <= \b4_nUAi[105]\;
    b4_nUAi(104) <= \b4_nUAi[104]\;
    b4_nUAi(103) <= \b4_nUAi[103]\;
    b4_nUAi(102) <= \b4_nUAi[102]\;
    b4_nUAi(101) <= \b4_nUAi[101]\;
    b4_nUAi(100) <= \b4_nUAi[100]\;
    b4_nUAi(99) <= \b4_nUAi[99]\;
    b4_nUAi(98) <= \b4_nUAi[98]\;
    b4_nUAi(97) <= \b4_nUAi[97]\;
    b4_nUAi(96) <= \b4_nUAi[96]\;
    b4_nUAi(95) <= \b4_nUAi[95]\;
    b4_nUAi(94) <= \b4_nUAi[94]\;
    b4_nUAi(93) <= \b4_nUAi[93]\;
    b4_nUAi(92) <= \b4_nUAi[92]\;
    b4_nUAi(91) <= \b4_nUAi[91]\;
    b4_nUAi(90) <= \b4_nUAi[90]\;
    b4_nUAi(89) <= \b4_nUAi[89]\;
    b4_nUAi(88) <= \b4_nUAi[88]\;
    b4_nUAi(87) <= \b4_nUAi[87]\;
    b4_nUAi(86) <= \b4_nUAi[86]\;
    b4_nUAi(85) <= \b4_nUAi[85]\;
    b4_nUAi(84) <= \b4_nUAi[84]\;
    b4_nUAi(83) <= \b4_nUAi[83]\;
    b4_nUAi(82) <= \b4_nUAi[82]\;
    b4_nUAi(81) <= \b4_nUAi[81]\;
    b4_nUAi(80) <= \b4_nUAi[80]\;
    b4_nUAi(79) <= \b4_nUAi[79]\;
    b4_nUAi(78) <= \b4_nUAi[78]\;
    b4_nUAi(77) <= \b4_nUAi[77]\;
    b4_nUAi(76) <= \b4_nUAi[76]\;
    b4_nUAi(75) <= \b4_nUAi[75]\;
    b4_nUAi(74) <= \b4_nUAi[74]\;
    b4_nUAi(73) <= \b4_nUAi[73]\;
    b4_nUAi(72) <= \b4_nUAi[72]\;
    b4_nUAi(71) <= \b4_nUAi[71]\;
    b4_nUAi(70) <= \b4_nUAi[70]\;
    b4_nUAi(69) <= \b4_nUAi[69]\;
    b4_nUAi(68) <= \b4_nUAi[68]\;
    b4_nUAi(67) <= \b4_nUAi[67]\;
    b4_nUAi(66) <= \b4_nUAi[66]\;
    b4_nUAi(65) <= \b4_nUAi[65]\;
    b4_nUAi(64) <= \b4_nUAi[64]\;
    b4_nUAi(63) <= \b4_nUAi[63]\;
    b4_nUAi(62) <= \b4_nUAi[62]\;
    b4_nUAi(61) <= \b4_nUAi[61]\;
    b4_nUAi(60) <= \b4_nUAi[60]\;
    b4_nUAi(59) <= \b4_nUAi[59]\;
    b4_nUAi(58) <= \b4_nUAi[58]\;
    b4_nUAi(57) <= \b4_nUAi[57]\;
    b4_nUAi(56) <= \b4_nUAi[56]\;
    b4_nUAi(55) <= \b4_nUAi[55]\;
    b4_nUAi(54) <= \b4_nUAi[54]\;
    b4_nUAi(53) <= \b4_nUAi[53]\;
    b4_nUAi(52) <= \b4_nUAi[52]\;
    b4_nUAi(51) <= \b4_nUAi[51]\;
    b4_nUAi(50) <= \b4_nUAi[50]\;
    b4_nUAi(49) <= \b4_nUAi[49]\;
    b4_nUAi(48) <= \b4_nUAi[48]\;
    b4_nUAi(47) <= \b4_nUAi[47]\;
    b4_nUAi(46) <= \b4_nUAi[46]\;
    b4_nUAi(45) <= \b4_nUAi[45]\;
    b4_nUAi(44) <= \b4_nUAi[44]\;
    b4_nUAi(43) <= \b4_nUAi[43]\;
    b4_nUAi(42) <= \b4_nUAi[42]\;
    b4_nUAi(41) <= \b4_nUAi[41]\;
    b4_nUAi(40) <= \b4_nUAi[40]\;
    b4_nUAi(39) <= \b4_nUAi[39]\;
    b4_nUAi(38) <= \b4_nUAi[38]\;
    b4_nUAi(37) <= \b4_nUAi[37]\;
    b4_nUAi(36) <= \b4_nUAi[36]\;
    b4_nUAi(35) <= \b4_nUAi[35]\;
    b4_nUAi(34) <= \b4_nUAi[34]\;
    b4_nUAi(33) <= \b4_nUAi[33]\;
    b4_nUAi(32) <= \b4_nUAi[32]\;
    b4_nUAi(31) <= \b4_nUAi[31]\;
    b4_nUAi(30) <= \b4_nUAi[30]\;
    b4_nUAi(29) <= \b4_nUAi[29]\;
    b4_nUAi(28) <= \b4_nUAi[28]\;
    b4_nUAi(27) <= \b4_nUAi[27]\;
    b4_nUAi(26) <= \b4_nUAi[26]\;
    b4_nUAi(25) <= \b4_nUAi[25]\;
    b4_nUAi(24) <= \b4_nUAi[24]\;
    b4_nUAi(23) <= \b4_nUAi[23]\;
    b4_nUAi(22) <= \b4_nUAi[22]\;
    b4_nUAi(21) <= \b4_nUAi[21]\;
    b4_nUAi(20) <= \b4_nUAi[20]\;
    b4_nUAi(19) <= \b4_nUAi[19]\;
    b4_nUAi(18) <= \b4_nUAi[18]\;
    b4_nUAi(17) <= \b4_nUAi[17]\;
    b4_nUAi(16) <= \b4_nUAi[16]\;
    b4_nUAi(15) <= \b4_nUAi[15]\;
    b4_nUAi(14) <= \b4_nUAi[14]\;
    b4_nUAi(13) <= \b4_nUAi[13]\;
    b4_nUAi(12) <= \b4_nUAi[12]\;
    b4_nUAi(11) <= \b4_nUAi[11]\;
    b4_nUAi(10) <= \b4_nUAi[10]\;
    b4_nUAi(9) <= \b4_nUAi[9]\;
    b4_nUAi(8) <= \b4_nUAi[8]\;
    b4_nUAi(7) <= \b4_nUAi[7]\;
    b4_nUAi(6) <= \b4_nUAi[6]\;
    b4_nUAi(5) <= \b4_nUAi[5]\;
    b4_nUAi(4) <= \b4_nUAi[4]\;
    b4_nUAi(3) <= \b4_nUAi[3]\;
    b4_nUAi(2) <= \b4_nUAi[2]\;
    b4_nUAi(1) <= \b4_nUAi[1]\;
    b4_nUAi(0) <= \b4_nUAi[0]\;

    \b6_OKctIF[169]\ : SLE
      port map(D => \b4_nUAi[333]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[334]\);
    
    \b6_OKctIF[41]\ : SLE
      port map(D => \b4_nUAi[461]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[462]\);
    
    \b6_OKctIF[269]\ : SLE
      port map(D => \b4_nUAi[233]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[234]\);
    
    \b6_OKctIF[147]\ : SLE
      port map(D => \b4_nUAi[355]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[356]\);
    
    \b6_OKctIF[58]\ : SLE
      port map(D => \b4_nUAi[444]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[445]\);
    
    \b6_OKctIF[55]\ : SLE
      port map(D => \b4_nUAi[447]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[448]\);
    
    \b6_OKctIF[352]\ : SLE
      port map(D => \b4_nUAi[150]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[151]\);
    
    \b6_OKctIF[430]\ : SLE
      port map(D => \b4_nUAi[72]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[73]\);
    
    \b6_OKctIF[204]\ : SLE
      port map(D => \b4_nUAi[298]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[299]\);
    
    \b6_OKctIF[374]\ : SLE
      port map(D => \b4_nUAi[128]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[129]\);
    
    \b6_OKctIF[284]\ : SLE
      port map(D => \b4_nUAi[218]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[219]\);
    
    \b6_OKctIF[2]\ : SLE
      port map(D => \b4_nUAi[500]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[501]\);
    
    \b6_OKctIF[260]\ : SLE
      port map(D => \b4_nUAi[242]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[243]\);
    
    \b6_OKctIF[156]\ : SLE
      port map(D => \b4_nUAi[346]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[347]\);
    
    \b6_OKctIF[47]\ : SLE
      port map(D => \b4_nUAi[455]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[456]\);
    
    \b6_OKctIF[212]\ : SLE
      port map(D => \b4_nUAi[290]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[291]\);
    
    \b6_OKctIF[165]\ : SLE
      port map(D => \b4_nUAi[337]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[338]\);
    
    \b6_OKctIF[477]\ : SLE
      port map(D => \b4_nUAi[25]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[26]\);
    
    \b6_OKctIF[472]\ : SLE
      port map(D => \b4_nUAi[30]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[31]\);
    
    \b6_OKctIF[46]\ : SLE
      port map(D => \b4_nUAi[456]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[457]\);
    
    \b6_OKctIF[43]\ : SLE
      port map(D => \b4_nUAi[459]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[460]\);
    
    \b6_OKctIF[208]\ : SLE
      port map(D => \b4_nUAi[294]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[295]\);
    
    \b6_OKctIF[288]\ : SLE
      port map(D => \b4_nUAi[214]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[215]\);
    
    \b6_OKctIF[405]\ : SLE
      port map(D => \b4_nUAi[97]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[98]\);
    
    \b6_OKctIF[246]\ : SLE
      port map(D => \b4_nUAi[256]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[257]\);
    
    \b6_OKctIF[485]\ : SLE
      port map(D => \b4_nUAi[17]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[18]\);
    
    \b6_OKctIF[312]\ : SLE
      port map(D => \b4_nUAi[190]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[191]\);
    
    \b6_OKctIF[251]\ : SLE
      port map(D => \b4_nUAi[251]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[252]\);
    
    \b6_OKctIF[116]\ : SLE
      port map(D => \b4_nUAi[386]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[387]\);
    
    \b6_OKctIF[498]\ : SLE
      port map(D => \b4_nUAi[4]\, CLK => IICE_comm2iice_4, EN => 
        \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[5]\);
    
    \b6_OKctIF[409]\ : SLE
      port map(D => \b4_nUAi[93]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[94]\);
    
    \b6_OKctIF[489]\ : SLE
      port map(D => \b4_nUAi[13]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[14]\);
    
    b6_OKctIF4 : CFG2
      generic map(INIT => x"8")

      port map(A => b7_PSyi_9u, B => IICE_comm2iice_3, Y => 
        \b6_OKctIF4\);
    
    \b6_OKctIF[401]\ : SLE
      port map(D => \b4_nUAi[101]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[102]\);
    
    \b6_OKctIF[481]\ : SLE
      port map(D => \b4_nUAi[21]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[22]\);
    
    \b6_OKctIF[334]\ : SLE
      port map(D => \b4_nUAi[168]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[169]\);
    
    \b6_OKctIF[428]\ : SLE
      port map(D => \b4_nUAi[74]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[75]\);
    
    \b6_OKctIF[341]\ : SLE
      port map(D => \b4_nUAi[161]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[162]\);
    
    \b6_OKctIF[211]\ : SLE
      port map(D => \b4_nUAi[291]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[292]\);
    
    \b6_OKctIF[100]\ : SLE
      port map(D => \b4_nUAi[402]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[403]\);
    
    \b6_OKctIF[437]\ : SLE
      port map(D => \b4_nUAi[65]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[66]\);
    
    \b6_OKctIF[42]\ : SLE
      port map(D => \b4_nUAi[460]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[461]\);
    
    \b6_OKctIF[348]\ : SLE
      port map(D => \b4_nUAi[154]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[155]\);
    
    \b6_OKctIF[194]\ : SLE
      port map(D => \b4_nUAi[308]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[309]\);
    
    \b6_OKctIF[180]\ : SLE
      port map(D => \b4_nUAi[322]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[323]\);
    
    \b6_OKctIF[403]\ : SLE
      port map(D => \b4_nUAi[99]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[100]\);
    
    \b6_OKctIF[483]\ : SLE
      port map(D => \b4_nUAi[19]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[20]\);
    
    \b6_OKctIF[432]\ : SLE
      port map(D => \b4_nUAi[70]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[71]\);
    
    \b6_OKctIF[375]\ : SLE
      port map(D => \b4_nUAi[127]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[128]\);
    
    \b6_OKctIF[275]\ : SLE
      port map(D => \b4_nUAi[227]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[228]\);
    
    \b6_OKctIF[49]\ : SLE
      port map(D => \b4_nUAi[453]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[454]\);
    
    \b6_OKctIF[377]\ : SLE
      port map(D => \b4_nUAi[125]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[126]\);
    
    \b6_OKctIF[503]\ : SLE
      port map(D => IICE_comm2iice_0, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[0]\);
    
    \b6_OKctIF[390]\ : SLE
      port map(D => \b4_nUAi[112]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[113]\);
    
    \b6_OKctIF[103]\ : SLE
      port map(D => \b4_nUAi[399]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[400]\);
    
    \b6_OKctIF[183]\ : SLE
      port map(D => \b4_nUAi[319]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[320]\);
    
    \b6_OKctIF[440]\ : SLE
      port map(D => \b4_nUAi[62]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[63]\);
    
    \b6_OKctIF[124]\ : SLE
      port map(D => \b4_nUAi[378]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[379]\);
    
    \b6_OKctIF[264]\ : SLE
      port map(D => \b4_nUAi[238]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[239]\);
    
    \b6_OKctIF[197]\ : SLE
      port map(D => \b4_nUAi[305]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[306]\);
    
    \b6_OKctIF[102]\ : SLE
      port map(D => \b4_nUAi[400]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[401]\);
    
    \b6_OKctIF[320]\ : SLE
      port map(D => \b4_nUAi[182]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[183]\);
    
    \b6_OKctIF[182]\ : SLE
      port map(D => \b4_nUAi[320]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[321]\);
    
    \b6_OKctIF[40]\ : SLE
      port map(D => \b4_nUAi[462]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[463]\);
    
    \b6_OKctIF[268]\ : SLE
      port map(D => \b4_nUAi[234]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[235]\);
    
    \b6_OKctIF[465]\ : SLE
      port map(D => \b4_nUAi[37]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[38]\);
    
    \b6_OKctIF[127]\ : SLE
      port map(D => \b4_nUAi[375]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[376]\);
    
    \b6_OKctIF[458]\ : SLE
      port map(D => \b4_nUAi[44]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[45]\);
    
    \b6_OKctIF[3]\ : SLE
      port map(D => \b4_nUAi[499]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[500]\);
    
    \b6_OKctIF[296]\ : SLE
      port map(D => \b4_nUAi[206]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[207]\);
    
    \b6_OKctIF[335]\ : SLE
      port map(D => \b4_nUAi[167]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[168]\);
    
    \b6_OKctIF[235]\ : SLE
      port map(D => \b4_nUAi[267]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[268]\);
    
    \b6_OKctIF[337]\ : SLE
      port map(D => \b4_nUAi[165]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[166]\);
    
    \b6_OKctIF[469]\ : SLE
      port map(D => \b4_nUAi[33]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[34]\);
    
    \b6_OKctIF[154]\ : SLE
      port map(D => \b4_nUAi[348]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[349]\);
    
    \b6_OKctIF[226]\ : SLE
      port map(D => \b4_nUAi[276]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[277]\);
    
    \b6_OKctIF[461]\ : SLE
      port map(D => \b4_nUAi[41]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[42]\);
    
    \b6_OKctIF[418]\ : SLE
      port map(D => \b4_nUAi[84]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[85]\);
    
    \b6_OKctIF[344]\ : SLE
      port map(D => \b4_nUAi[158]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[159]\);
    
    \b6_OKctIF[350]\ : SLE
      port map(D => \b4_nUAi[152]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[153]\);
    
    \b6_OKctIF[447]\ : SLE
      port map(D => \b4_nUAi[55]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[56]\);
    
    \b6_OKctIF[160]\ : SLE
      port map(D => \b4_nUAi[342]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[343]\);
    
    \b6_OKctIF[404]\ : SLE
      port map(D => \b4_nUAi[98]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[99]\);
    
    \b6_OKctIF[24]\ : SLE
      port map(D => \b4_nUAi[478]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[479]\);
    
    \b6_OKctIF[484]\ : SLE
      port map(D => \b4_nUAi[18]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[19]\);
    
    \b6_OKctIF[463]\ : SLE
      port map(D => \b4_nUAi[39]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[40]\);
    
    \b6_OKctIF[442]\ : SLE
      port map(D => \b4_nUAi[60]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[61]\);
    
    \b6_OKctIF[178]\ : SLE
      port map(D => \b4_nUAi[324]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[325]\);
    
    \b6_OKctIF[391]\ : SLE
      port map(D => \b4_nUAi[111]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[112]\);
    
    \b6_OKctIF[157]\ : SLE
      port map(D => \b4_nUAi[345]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[346]\);
    
    \b6_OKctIF[398]\ : SLE
      port map(D => \b4_nUAi[104]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[105]\);
    
    \b6_OKctIF[163]\ : SLE
      port map(D => \b4_nUAi[339]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[340]\);
    
    \b6_OKctIF[114]\ : SLE
      port map(D => \b4_nUAi[388]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[389]\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \b6_OKctIF[21]\ : SLE
      port map(D => \b4_nUAi[481]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[482]\);
    
    \b6_OKctIF[321]\ : SLE
      port map(D => \b4_nUAi[181]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[182]\);
    
    \b6_OKctIF[310]\ : SLE
      port map(D => \b4_nUAi[192]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[193]\);
    
    \b6_OKctIF[490]\ : SLE
      port map(D => \b4_nUAi[12]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[13]\);
    
    \b6_OKctIF[328]\ : SLE
      port map(D => \b4_nUAi[174]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[175]\);
    
    \b6_OKctIF[162]\ : SLE
      port map(D => \b4_nUAi[340]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[341]\);
    
    \b6_OKctIF[5]\ : SLE
      port map(D => \b4_nUAi[497]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[498]\);
    
    \b6_OKctIF[27]\ : SLE
      port map(D => \b4_nUAi[475]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[476]\);
    
    \b6_OKctIF[207]\ : SLE
      port map(D => \b4_nUAi[295]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[296]\);
    
    \b6_OKctIF[287]\ : SLE
      port map(D => \b4_nUAi[215]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[216]\);
    
    \b6_OKctIF[256]\ : SLE
      port map(D => \b4_nUAi[246]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[247]\);
    
    \b6_OKctIF[54]\ : SLE
      port map(D => \b4_nUAi[448]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[449]\);
    
    \b6_OKctIF[273]\ : SLE
      port map(D => \b4_nUAi[229]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[230]\);
    
    \b6_OKctIF[117]\ : SLE
      port map(D => \b4_nUAi[385]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[386]\);
    
    \b6_OKctIF[26]\ : SLE
      port map(D => \b4_nUAi[476]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[477]\);
    
    \b6_OKctIF[23]\ : SLE
      port map(D => \b4_nUAi[479]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[480]\);
    
    \b6_OKctIF[373]\ : SLE
      port map(D => \b4_nUAi[129]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[130]\);
    
    \b6_OKctIF[420]\ : SLE
      port map(D => \b4_nUAi[82]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[83]\);
    
    \b6_OKctIF[376]\ : SLE
      port map(D => \b4_nUAi[126]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[127]\);
    
    \b6_OKctIF[171]\ : SLE
      port map(D => \b4_nUAi[331]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[332]\);
    
    \b6_OKctIF[51]\ : SLE
      port map(D => \b4_nUAi[451]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[452]\);
    
    \b6_OKctIF[345]\ : SLE
      port map(D => \b4_nUAi[157]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[158]\);
    
    \b6_OKctIF[245]\ : SLE
      port map(D => \b4_nUAi[257]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[258]\);
    
    \b6_OKctIF[138]\ : SLE
      port map(D => \b4_nUAi[364]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[365]\);
    
    \b6_OKctIF[347]\ : SLE
      port map(D => \b4_nUAi[155]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[156]\);
    
    \b6_OKctIF[216]\ : SLE
      port map(D => \b4_nUAi[286]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[287]\);
    
    \b6_OKctIF[57]\ : SLE
      port map(D => \b4_nUAi[445]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[446]\);
    
    \b6_OKctIF[351]\ : SLE
      port map(D => \b4_nUAi[151]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[152]\);
    
    \b6_OKctIF[56]\ : SLE
      port map(D => \b4_nUAi[446]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[447]\);
    
    \b6_OKctIF[53]\ : SLE
      port map(D => \b4_nUAi[449]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[450]\);
    
    \b6_OKctIF[358]\ : SLE
      port map(D => \b4_nUAi[144]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[145]\);
    
    \b6_OKctIF[202]\ : SLE
      port map(D => \b4_nUAi[300]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[301]\);
    
    \b6_OKctIF[38]\ : SLE
      port map(D => \b4_nUAi[464]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[465]\);
    
    \b6_OKctIF[35]\ : SLE
      port map(D => \b4_nUAi[467]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[468]\);
    
    \b6_OKctIF[282]\ : SLE
      port map(D => \b4_nUAi[220]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[221]\);
    
    \b6_OKctIF[501]\ : SLE
      port map(D => \b4_nUAi[1]\, CLK => IICE_comm2iice_4, EN => 
        \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[2]\);
    
    \b6_OKctIF[464]\ : SLE
      port map(D => \b4_nUAi[38]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[39]\);
    
    \b6_OKctIF[394]\ : SLE
      port map(D => \b4_nUAi[108]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[109]\);
    
    \b6_OKctIF[22]\ : SLE
      port map(D => \b4_nUAi[480]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[481]\);
    
    \b6_OKctIF[233]\ : SLE
      port map(D => \b4_nUAi[269]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[270]\);
    
    \b6_OKctIF[497]\ : SLE
      port map(D => \b4_nUAi[5]\, CLK => IICE_comm2iice_4, EN => 
        \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[6]\);
    
    \b6_OKctIF[333]\ : SLE
      port map(D => \b4_nUAi[169]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[170]\);
    
    \b6_OKctIF[29]\ : SLE
      port map(D => \b4_nUAi[473]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[474]\);
    
    \b6_OKctIF[492]\ : SLE
      port map(D => \b4_nUAi[10]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[11]\);
    
    \b6_OKctIF[450]\ : SLE
      port map(D => \b4_nUAi[52]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[53]\);
    
    \b6_OKctIF[302]\ : SLE
      port map(D => \b4_nUAi[200]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[201]\);
    
    \b6_OKctIF[382]\ : SLE
      port map(D => \b4_nUAi[120]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[121]\);
    
    \b6_OKctIF[336]\ : SLE
      port map(D => \b4_nUAi[166]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[167]\);
    
    \b6_OKctIF[324]\ : SLE
      port map(D => \b4_nUAi[178]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[179]\);
    
    \b6_OKctIF[311]\ : SLE
      port map(D => \b4_nUAi[191]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[192]\);
    
    \b6_OKctIF[131]\ : SLE
      port map(D => \b4_nUAi[371]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[372]\);
    
    \b6_OKctIF[106]\ : SLE
      port map(D => \b4_nUAi[396]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[397]\);
    
    \b6_OKctIF[9]\ : SLE
      port map(D => \b4_nUAi[493]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[494]\);
    
    \b6_OKctIF[318]\ : SLE
      port map(D => \b4_nUAi[184]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[185]\);
    
    \b6_OKctIF[186]\ : SLE
      port map(D => \b4_nUAi[316]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[317]\);
    
    \b6_OKctIF[427]\ : SLE
      port map(D => \b4_nUAi[75]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[76]\);
    
    \b6_OKctIF[422]\ : SLE
      port map(D => \b4_nUAi[80]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[81]\);
    
    \b6_OKctIF[379]\ : SLE
      port map(D => \b4_nUAi[123]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[124]\);
    
    \b6_OKctIF[267]\ : SLE
      port map(D => \b4_nUAi[235]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[236]\);
    
    \b6_OKctIF[476]\ : SLE
      port map(D => \b4_nUAi[26]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[27]\);
    
    \b6_OKctIF[20]\ : SLE
      port map(D => \b4_nUAi[482]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[483]\);
    
    \b6_OKctIF[52]\ : SLE
      port map(D => \b4_nUAi[450]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[451]\);
    
    \b6_OKctIF[410]\ : SLE
      port map(D => \b4_nUAi[92]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[93]\);
    
    \b6_OKctIF[201]\ : SLE
      port map(D => \b4_nUAi[301]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[302]\);
    
    \b6_OKctIF[179]\ : SLE
      port map(D => \b4_nUAi[323]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[324]\);
    
    \b6_OKctIF[59]\ : SLE
      port map(D => \b4_nUAi[443]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[444]\);
    
    \b6_OKctIF[281]\ : SLE
      port map(D => \b4_nUAi[221]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[222]\);
    
    \b6_OKctIF[279]\ : SLE
      port map(D => \b4_nUAi[223]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[224]\);
    
    \b6_OKctIF[148]\ : SLE
      port map(D => \b4_nUAi[354]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[355]\);
    
    \b6_OKctIF[18]\ : SLE
      port map(D => \b4_nUAi[484]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[485]\);
    
    \b6_OKctIF[15]\ : SLE
      port map(D => \b4_nUAi[487]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[488]\);
    
    \b6_OKctIF[270]\ : SLE
      port map(D => \b4_nUAi[232]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[233]\);
    
    \b6_OKctIF[395]\ : SLE
      port map(D => \b4_nUAi[107]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[108]\);
    
    \b6_OKctIF[295]\ : SLE
      port map(D => \b4_nUAi[207]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[208]\);
    
    \b6_OKctIF[175]\ : SLE
      port map(D => \b4_nUAi[327]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[328]\);
    
    \b6_OKctIF[397]\ : SLE
      port map(D => \b4_nUAi[105]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[106]\);
    
    \b6_OKctIF[354]\ : SLE
      port map(D => \b4_nUAi[148]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[149]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \b6_OKctIF[50]\ : SLE
      port map(D => \b4_nUAi[452]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[453]\);
    
    \b6_OKctIF[457]\ : SLE
      port map(D => \b4_nUAi[45]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[46]\);
    
    \b6_OKctIF[262]\ : SLE
      port map(D => \b4_nUAi[240]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[241]\);
    
    \b6_OKctIF[452]\ : SLE
      port map(D => \b4_nUAi[50]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[51]\);
    
    \b6_OKctIF[78]\ : SLE
      port map(D => \b4_nUAi[424]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[425]\);
    
    \b6_OKctIF[75]\ : SLE
      port map(D => \b4_nUAi[427]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[428]\);
    
    \b6_OKctIF[339]\ : SLE
      port map(D => \b4_nUAi[163]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[164]\);
    
    \b6_OKctIF[325]\ : SLE
      port map(D => \b4_nUAi[177]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[178]\);
    
    \b6_OKctIF[225]\ : SLE
      port map(D => \b4_nUAi[277]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[278]\);
    
    \b6_OKctIF[327]\ : SLE
      port map(D => \b4_nUAi[175]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[176]\);
    
    \b6_OKctIF[436]\ : SLE
      port map(D => \b4_nUAi[66]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[67]\);
    
    \b6_OKctIF[243]\ : SLE
      port map(D => \b4_nUAi[259]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[260]\);
    
    \b6_OKctIF[343]\ : SLE
      port map(D => \b4_nUAi[159]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[160]\);
    
    \b6_OKctIF[68]\ : SLE
      port map(D => \b4_nUAi[434]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[435]\);
    
    \b6_OKctIF[65]\ : SLE
      port map(D => \b4_nUAi[437]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[438]\);
    
    \b6_OKctIF[362]\ : SLE
      port map(D => \b4_nUAi[140]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[141]\);
    
    \b6_OKctIF[139]\ : SLE
      port map(D => \b4_nUAi[363]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[364]\);
    
    \b6_OKctIF[314]\ : SLE
      port map(D => \b4_nUAi[188]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[189]\);
    
    \b6_OKctIF[239]\ : SLE
      port map(D => \b4_nUAi[263]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[264]\);
    
    \b6_OKctIF[346]\ : SLE
      port map(D => \b4_nUAi[156]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[157]\);
    
    \b6_OKctIF[141]\ : SLE
      port map(D => \b4_nUAi[361]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[362]\);
    
    \b6_OKctIF[417]\ : SLE
      port map(D => \b4_nUAi[85]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[86]\);
    
    \b6_OKctIF[166]\ : SLE
      port map(D => \b4_nUAi[336]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[337]\);
    
    \b6_OKctIF[412]\ : SLE
      port map(D => \b4_nUAi[90]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[91]\);
    
    \b6_OKctIF[230]\ : SLE
      port map(D => \b4_nUAi[272]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[273]\);
    
    \b6_OKctIF[135]\ : SLE
      port map(D => \b4_nUAi[367]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[368]\);
    
    \b6_OKctIF[408]\ : SLE
      port map(D => \b4_nUAi[94]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[95]\);
    
    \b6_OKctIF[488]\ : SLE
      port map(D => \b4_nUAi[14]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[15]\);
    
    \b6_OKctIF[261]\ : SLE
      port map(D => \b4_nUAi[241]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[242]\);
    
    \b6_OKctIF[355]\ : SLE
      port map(D => \b4_nUAi[147]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[148]\);
    
    \b6_OKctIF[255]\ : SLE
      port map(D => \b4_nUAi[247]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[248]\);
    
    \b6_OKctIF[357]\ : SLE
      port map(D => \b4_nUAi[145]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[146]\);
    
    \b6_OKctIF[98]\ : SLE
      port map(D => \b4_nUAi[404]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[405]\);
    
    \b6_OKctIF[95]\ : SLE
      port map(D => \b4_nUAi[407]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[408]\);
    
    \b6_OKctIF[274]\ : SLE
      port map(D => \b4_nUAi[228]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[229]\);
    
    \b6_OKctIF[198]\ : SLE
      port map(D => \b4_nUAi[304]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[305]\);
    
    \b6_OKctIF[104]\ : SLE
      port map(D => \b4_nUAi[398]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[399]\);
    
    \b6_OKctIF[184]\ : SLE
      port map(D => \b4_nUAi[318]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[319]\);
    
    \b6_OKctIF[278]\ : SLE
      port map(D => \b4_nUAi[224]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[225]\);
    
    \b6_OKctIF[300]\ : SLE
      port map(D => \b4_nUAi[202]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[203]\);
    
    \b6_OKctIF[475]\ : SLE
      port map(D => \b4_nUAi[27]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[28]\);
    
    \b6_OKctIF[380]\ : SLE
      port map(D => \b4_nUAi[122]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[123]\);
    
    \b6_OKctIF[315]\ : SLE
      port map(D => \b4_nUAi[187]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[188]\);
    
    \b6_OKctIF[215]\ : SLE
      port map(D => \b4_nUAi[287]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[288]\);
    
    \b6_OKctIF[349]\ : SLE
      port map(D => \b4_nUAi[153]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[154]\);
    
    \b6_OKctIF[317]\ : SLE
      port map(D => \b4_nUAi[185]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[186]\);
    
    \b6_OKctIF[128]\ : SLE
      port map(D => \b4_nUAi[374]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[375]\);
    
    \b6_OKctIF[446]\ : SLE
      port map(D => \b4_nUAi[56]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[57]\);
    
    \b6_OKctIF[107]\ : SLE
      port map(D => \b4_nUAi[395]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[396]\);
    
    \b6_OKctIF[187]\ : SLE
      port map(D => \b4_nUAi[315]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[316]\);
    
    \b6_OKctIF[149]\ : SLE
      port map(D => \b4_nUAi[353]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[354]\);
    
    \b6_OKctIF[479]\ : SLE
      port map(D => \b4_nUAi[23]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[24]\);
    
    \b6_OKctIF[293]\ : SLE
      port map(D => \b4_nUAi[209]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[210]\);
    
    \b6_OKctIF[249]\ : SLE
      port map(D => \b4_nUAi[253]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[254]\);
    
    \b6_OKctIF[393]\ : SLE
      port map(D => \b4_nUAi[109]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[110]\);
    
    \b6_OKctIF[34]\ : SLE
      port map(D => \b4_nUAi[468]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[469]\);
    
    \b6_OKctIF[7]\ : SLE
      port map(D => \b4_nUAi[495]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[496]\);
    
    \b6_OKctIF[471]\ : SLE
      port map(D => \b4_nUAi[31]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[32]\);
    
    \b6_OKctIF[234]\ : SLE
      port map(D => \b4_nUAi[268]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[269]\);
    
    \b6_OKctIF[396]\ : SLE
      port map(D => \b4_nUAi[106]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[107]\);
    
    \b6_OKctIF[240]\ : SLE
      port map(D => \b4_nUAi[262]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[263]\);
    
    \b6_OKctIF[191]\ : SLE
      port map(D => \b4_nUAi[311]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[312]\);
    
    \b6_OKctIF[206]\ : SLE
      port map(D => \b4_nUAi[296]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[297]\);
    
    \b6_OKctIF[145]\ : SLE
      port map(D => \b4_nUAi[357]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[358]\);
    
    \b6_OKctIF[286]\ : SLE
      port map(D => \b4_nUAi[216]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[217]\);
    
    \b6_OKctIF[223]\ : SLE
      port map(D => \b4_nUAi[279]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[280]\);
    
    \b6_OKctIF[170]\ : SLE
      port map(D => \b4_nUAi[332]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[333]\);
    
    \b6_OKctIF[88]\ : SLE
      port map(D => \b4_nUAi[414]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[415]\);
    
    \b6_OKctIF[85]\ : SLE
      port map(D => \b4_nUAi[417]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[418]\);
    
    \b6_OKctIF[6]\ : SLE
      port map(D => \b4_nUAi[496]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[497]\);
    
    \b6_OKctIF[31]\ : SLE
      port map(D => \b4_nUAi[471]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[472]\);
    
    \b6_OKctIF[473]\ : SLE
      port map(D => \b4_nUAi[29]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[30]\);
    
    \b6_OKctIF[323]\ : SLE
      port map(D => \b4_nUAi[179]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[180]\);
    
    \b6_OKctIF[468]\ : SLE
      port map(D => \b4_nUAi[34]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[35]\);
    
    \b6_OKctIF[238]\ : SLE
      port map(D => \b4_nUAi[264]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[265]\);
    
    \b6_OKctIF[435]\ : SLE
      port map(D => \b4_nUAi[67]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[68]\);
    
    \b6_OKctIF[326]\ : SLE
      port map(D => \b4_nUAi[176]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[177]\);
    
    \b6_OKctIF[173]\ : SLE
      port map(D => \b4_nUAi[329]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[330]\);
    
    \b6_OKctIF[158]\ : SLE
      port map(D => \b4_nUAi[344]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[345]\);
    
    \b6_OKctIF[121]\ : SLE
      port map(D => \b4_nUAi[381]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[382]\);
    
    \b6_OKctIF[37]\ : SLE
      port map(D => \b4_nUAi[465]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[466]\);
    
    \b6_OKctIF[36]\ : SLE
      port map(D => \b4_nUAi[466]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[467]\);
    
    \b6_OKctIF[33]\ : SLE
      port map(D => \b4_nUAi[469]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[470]\);
    
    \b6_OKctIF[172]\ : SLE
      port map(D => \b4_nUAi[330]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[331]\);
    
    \b6_OKctIF[164]\ : SLE
      port map(D => \b4_nUAi[338]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[339]\);
    
    \b6_OKctIF[439]\ : SLE
      port map(D => \b4_nUAi[63]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[64]\);
    
    \b6_OKctIF[4]\ : SLE
      port map(D => \b4_nUAi[498]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[499]\);
    
    \b6_OKctIF[301]\ : SLE
      port map(D => \b4_nUAi[201]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[202]\);
    
    \b6_OKctIF[381]\ : SLE
      port map(D => \b4_nUAi[121]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[122]\);
    
    \b6_OKctIF[308]\ : SLE
      port map(D => \b4_nUAi[194]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[195]\);
    
    \b6_OKctIF[388]\ : SLE
      port map(D => \b4_nUAi[114]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[115]\);
    
    \b6_OKctIF[360]\ : SLE
      port map(D => \b4_nUAi[142]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[143]\);
    
    \b6_OKctIF[431]\ : SLE
      port map(D => \b4_nUAi[71]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[72]\);
    
    \b6_OKctIF[118]\ : SLE
      port map(D => \b4_nUAi[384]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[385]\);
    
    \b6_OKctIF[14]\ : SLE
      port map(D => \b4_nUAi[488]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[489]\);
    
    \b6_OKctIF[253]\ : SLE
      port map(D => \b4_nUAi[249]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[250]\);
    
    \b6_OKctIF[130]\ : SLE
      port map(D => \b4_nUAi[372]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[373]\);
    
    \b6_OKctIF[353]\ : SLE
      port map(D => \b4_nUAi[149]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[150]\);
    
    \b6_OKctIF[167]\ : SLE
      port map(D => \b4_nUAi[335]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[336]\);
    
    \b6_OKctIF[433]\ : SLE
      port map(D => \b4_nUAi[69]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[70]\);
    
    \b6_OKctIF[400]\ : SLE
      port map(D => \b4_nUAi[102]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[103]\);
    
    \b6_OKctIF[399]\ : SLE
      port map(D => \b4_nUAi[103]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[104]\);
    
    \b6_OKctIF[480]\ : SLE
      port map(D => \b4_nUAi[22]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[23]\);
    
    \b6_OKctIF[496]\ : SLE
      port map(D => \b4_nUAi[6]\, CLK => IICE_comm2iice_4, EN => 
        \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[7]\);
    
    \b6_OKctIF[356]\ : SLE
      port map(D => \b4_nUAi[146]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[147]\);
    
    \b6_OKctIF[151]\ : SLE
      port map(D => \b4_nUAi[351]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[352]\);
    
    \b6_OKctIF[11]\ : SLE
      port map(D => \b4_nUAi[491]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[492]\);
    
    \b6_OKctIF[133]\ : SLE
      port map(D => \b4_nUAi[369]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[370]\);
    
    \b6_OKctIF[74]\ : SLE
      port map(D => \b4_nUAi[428]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[429]\);
    
    \b6_OKctIF[32]\ : SLE
      port map(D => \b4_nUAi[470]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[471]\);
    
    \b6_OKctIF[199]\ : SLE
      port map(D => \b4_nUAi[303]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[304]\);
    
    \b6_OKctIF[299]\ : SLE
      port map(D => \b4_nUAi[203]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[204]\);
    
    \b6_OKctIF[244]\ : SLE
      port map(D => \b4_nUAi[258]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[259]\);
    
    \b6_OKctIF[329]\ : SLE
      port map(D => \b4_nUAi[173]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[174]\);
    
    \b6_OKctIF[39]\ : SLE
      port map(D => \b4_nUAi[463]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[464]\);
    
    \b6_OKctIF[213]\ : SLE
      port map(D => \b4_nUAi[289]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[290]\);
    
    \b6_OKctIF[17]\ : SLE
      port map(D => \b4_nUAi[485]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[486]\);
    
    \b6_OKctIF[426]\ : SLE
      port map(D => \b4_nUAi[76]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[77]\);
    
    \b6_OKctIF[266]\ : SLE
      port map(D => \b4_nUAi[236]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[237]\);
    
    \b6_OKctIF[132]\ : SLE
      port map(D => \b4_nUAi[370]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[371]\);
    
    \b6_OKctIF[64]\ : SLE
      port map(D => \b4_nUAi[438]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[439]\);
    
    \b6_OKctIF[313]\ : SLE
      port map(D => \b4_nUAi[189]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[190]\);
    
    \b6_OKctIF[474]\ : SLE
      port map(D => \b4_nUAi[28]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[29]\);
    
    \b6_OKctIF[16]\ : SLE
      port map(D => \b4_nUAi[486]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[487]\);
    
    \b6_OKctIF[13]\ : SLE
      port map(D => \b4_nUAi[489]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[490]\);
    
    \b6_OKctIF[71]\ : SLE
      port map(D => \b4_nUAi[431]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[432]\);
    
    \b6_OKctIF[290]\ : SLE
      port map(D => \b4_nUAi[212]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[213]\);
    
    \b6_OKctIF[248]\ : SLE
      port map(D => \b4_nUAi[254]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[255]\);
    
    \b6_OKctIF[195]\ : SLE
      port map(D => \b4_nUAi[307]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[308]\);
    
    \b6_OKctIF[129]\ : SLE
      port map(D => \b4_nUAi[373]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[374]\);
    
    \b6_OKctIF[445]\ : SLE
      port map(D => \b4_nUAi[57]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[58]\);
    
    \b6_OKctIF[316]\ : SLE
      port map(D => \b4_nUAi[186]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[187]\);
    
    \b6_OKctIF[229]\ : SLE
      port map(D => \b4_nUAi[273]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[274]\);
    
    \b6_OKctIF[111]\ : SLE
      port map(D => \b4_nUAi[391]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[392]\);
    
    \b6_OKctIF[61]\ : SLE
      port map(D => \b4_nUAi[441]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[442]\);
    
    \b6_OKctIF[77]\ : SLE
      port map(D => \b4_nUAi[425]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[426]\);
    
    \b6_OKctIF[30]\ : SLE
      port map(D => \b4_nUAi[472]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[473]\);
    
    \b6_OKctIF[220]\ : SLE
      port map(D => \b4_nUAi[282]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[283]\);
    
    \b6_OKctIF[125]\ : SLE
      port map(D => \b4_nUAi[377]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[378]\);
    
    \b6_OKctIF[76]\ : SLE
      port map(D => \b4_nUAi[426]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[427]\);
    
    \b6_OKctIF[73]\ : SLE
      port map(D => \b4_nUAi[429]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[430]\);
    
    \b6_OKctIF[449]\ : SLE
      port map(D => \b4_nUAi[53]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[54]\);
    
    \b6_OKctIF[304]\ : SLE
      port map(D => \b4_nUAi[198]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[199]\);
    
    \b6_OKctIF[67]\ : SLE
      port map(D => \b4_nUAi[435]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[436]\);
    
    \b6_OKctIF[384]\ : SLE
      port map(D => \b4_nUAi[118]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[119]\);
    
    \b6_OKctIF[361]\ : SLE
      port map(D => \b4_nUAi[141]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[142]\);
    
    \b6_OKctIF[277]\ : SLE
      port map(D => \b4_nUAi[225]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[226]\);
    
    \b6_OKctIF[407]\ : SLE
      port map(D => \b4_nUAi[95]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[96]\);
    
    \b6_OKctIF[66]\ : SLE
      port map(D => \b4_nUAi[436]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[437]\);
    
    \b6_OKctIF[63]\ : SLE
      port map(D => \b4_nUAi[439]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[440]\);
    
    \b6_OKctIF[487]\ : SLE
      port map(D => \b4_nUAi[15]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[16]\);
    
    \b6_OKctIF[368]\ : SLE
      port map(D => \b4_nUAi[134]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[135]\);
    
    \b6_OKctIF[441]\ : SLE
      port map(D => \b4_nUAi[61]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[62]\);
    
    \b6_OKctIF[402]\ : SLE
      port map(D => \b4_nUAi[100]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[101]\);
    
    \b6_OKctIF[359]\ : SLE
      port map(D => \b4_nUAi[143]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[144]\);
    
    \b6_OKctIF[482]\ : SLE
      port map(D => \b4_nUAi[20]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[21]\);
    
    \b6_OKctIF[94]\ : SLE
      port map(D => \b4_nUAi[408]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[409]\);
    
    \b6_OKctIF[456]\ : SLE
      port map(D => \b4_nUAi[46]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[47]\);
    
    \b6_OKctIF[140]\ : SLE
      port map(D => \b4_nUAi[362]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[363]\);
    
    \b6_OKctIF[12]\ : SLE
      port map(D => \b4_nUAi[490]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[491]\);
    
    \b6_OKctIF[443]\ : SLE
      port map(D => \b4_nUAi[59]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[60]\);
    
    \b6_OKctIF[434]\ : SLE
      port map(D => \b4_nUAi[68]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[69]\);
    
    \b6_OKctIF[19]\ : SLE
      port map(D => \b4_nUAi[483]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[484]\);
    
    \b6_OKctIF[159]\ : SLE
      port map(D => \b4_nUAi[343]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[344]\);
    
    \b6_OKctIF[460]\ : SLE
      port map(D => \b4_nUAi[42]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[43]\);
    
    \b6_OKctIF[259]\ : SLE
      port map(D => \b4_nUAi[243]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[244]\);
    
    \b6_OKctIF[91]\ : SLE
      port map(D => \b4_nUAi[411]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[412]\);
    
    \b6_OKctIF[143]\ : SLE
      port map(D => \b4_nUAi[359]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[360]\);
    
    \b6_OKctIF[500]\ : SLE
      port map(D => \b4_nUAi[2]\, CLK => IICE_comm2iice_4, EN => 
        \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[3]\);
    
    \b6_OKctIF[319]\ : SLE
      port map(D => \b4_nUAi[183]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[184]\);
    
    \b6_OKctIF[250]\ : SLE
      port map(D => \b4_nUAi[252]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[253]\);
    
    \b6_OKctIF[72]\ : SLE
      port map(D => \b4_nUAi[430]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[431]\);
    
    \b6_OKctIF[155]\ : SLE
      port map(D => \b4_nUAi[347]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[348]\);
    
    \b6_OKctIF[416]\ : SLE
      port map(D => \b4_nUAi[86]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[87]\);
    
    \b6_OKctIF[97]\ : SLE
      port map(D => \b4_nUAi[405]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[406]\);
    
    \b6_OKctIF[272]\ : SLE
      port map(D => \b4_nUAi[230]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[231]\);
    
    \b6_OKctIF[142]\ : SLE
      port map(D => \b4_nUAi[360]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[361]\);
    
    \b6_OKctIF[79]\ : SLE
      port map(D => \b4_nUAi[423]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[424]\);
    
    \b6_OKctIF[294]\ : SLE
      port map(D => \b4_nUAi[208]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[209]\);
    
    \b6_OKctIF[10]\ : SLE
      port map(D => \b4_nUAi[492]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[493]\);
    
    \b6_OKctIF[96]\ : SLE
      port map(D => \b4_nUAi[406]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[407]\);
    
    \b6_OKctIF[93]\ : SLE
      port map(D => \b4_nUAi[409]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[410]\);
    
    \b6_OKctIF[62]\ : SLE
      port map(D => \b4_nUAi[440]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[441]\);
    
    \b6_OKctIF[237]\ : SLE
      port map(D => \b4_nUAi[265]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[266]\);
    
    \b6_OKctIF[119]\ : SLE
      port map(D => \b4_nUAi[383]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[384]\);
    
    \b6_OKctIF[219]\ : SLE
      port map(D => \b4_nUAi[283]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[284]\);
    
    \b6_OKctIF[69]\ : SLE
      port map(D => \b4_nUAi[433]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[434]\);
    
    \b6_OKctIF[305]\ : SLE
      port map(D => \b4_nUAi[197]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[198]\);
    
    \b6_OKctIF[205]\ : SLE
      port map(D => \b4_nUAi[297]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[298]\);
    
    \b6_OKctIF[385]\ : SLE
      port map(D => \b4_nUAi[117]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[118]\);
    
    \b6_OKctIF[307]\ : SLE
      port map(D => \b4_nUAi[195]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[196]\);
    
    \b6_OKctIF[285]\ : SLE
      port map(D => \b4_nUAi[217]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[218]\);
    
    \b6_OKctIF[387]\ : SLE
      port map(D => \b4_nUAi[115]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[116]\);
    
    \b6_OKctIF[372]\ : SLE
      port map(D => \b4_nUAi[130]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[131]\);
    
    \b6_OKctIF[298]\ : SLE
      port map(D => \b4_nUAi[204]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[205]\);
    
    \b6_OKctIF[495]\ : SLE
      port map(D => \b4_nUAi[7]\, CLK => IICE_comm2iice_4, EN => 
        \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[8]\);
    
    \b6_OKctIF[224]\ : SLE
      port map(D => \b4_nUAi[278]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[279]\);
    
    \b6_OKctIF[210]\ : SLE
      port map(D => \b4_nUAi[292]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[293]\);
    
    \b6_OKctIF[115]\ : SLE
      port map(D => \b4_nUAi[387]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[388]\);
    
    \b6_OKctIF[0]\ : SLE
      port map(D => \b4_nUAi[502]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b12_PSyi_XlK_qHv);
    
    \b6_OKctIF[84]\ : SLE
      port map(D => \b4_nUAi[418]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[419]\);
    
    \b6_OKctIF[176]\ : SLE
      port map(D => \b4_nUAi[326]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[327]\);
    
    \b6_OKctIF[70]\ : SLE
      port map(D => \b4_nUAi[432]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[433]\);
    
    \b6_OKctIF[364]\ : SLE
      port map(D => \b4_nUAi[138]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[139]\);
    
    \b6_OKctIF[228]\ : SLE
      port map(D => \b4_nUAi[274]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[275]\);
    
    \b6_OKctIF[60]\ : SLE
      port map(D => \b4_nUAi[442]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[443]\);
    
    \b6_OKctIF[467]\ : SLE
      port map(D => \b4_nUAi[35]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[36]\);
    
    \b6_OKctIF[425]\ : SLE
      port map(D => \b4_nUAi[77]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[78]\);
    
    \b6_OKctIF[81]\ : SLE
      port map(D => \b4_nUAi[421]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[422]\);
    
    \b6_OKctIF[499]\ : SLE
      port map(D => \b4_nUAi[3]\, CLK => IICE_comm2iice_4, EN => 
        \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[4]\);
    
    \b6_OKctIF[462]\ : SLE
      port map(D => \b4_nUAi[40]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[41]\);
    
    \b6_OKctIF[271]\ : SLE
      port map(D => \b4_nUAi[231]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[232]\);
    
    \b6_OKctIF[232]\ : SLE
      port map(D => \b4_nUAi[270]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[271]\);
    
    \b6_OKctIF[92]\ : SLE
      port map(D => \b4_nUAi[410]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[411]\);
    
    \b6_OKctIF[491]\ : SLE
      port map(D => \b4_nUAi[11]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[12]\);
    
    \b6_OKctIF[444]\ : SLE
      port map(D => \b4_nUAi[58]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[59]\);
    
    \b6_OKctIF[99]\ : SLE
      port map(D => \b4_nUAi[403]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[404]\);
    
    \b6_OKctIF[87]\ : SLE
      port map(D => \b4_nUAi[415]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[416]\);
    
    \b6_OKctIF[429]\ : SLE
      port map(D => \b4_nUAi[73]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[74]\);
    
    \b6_OKctIF[190]\ : SLE
      port map(D => \b4_nUAi[312]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[313]\);
    
    \b6_OKctIF[86]\ : SLE
      port map(D => \b4_nUAi[416]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[417]\);
    
    \b6_OKctIF[83]\ : SLE
      port map(D => \b4_nUAi[419]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[420]\);
    
    \b6_OKctIF[493]\ : SLE
      port map(D => \b4_nUAi[9]\, CLK => IICE_comm2iice_4, EN => 
        \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[10]\);
    
    \b6_OKctIF[332]\ : SLE
      port map(D => \b4_nUAi[170]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[171]\);
    
    \b6_OKctIF[254]\ : SLE
      port map(D => \b4_nUAi[248]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[249]\);
    
    \b6_OKctIF[421]\ : SLE
      port map(D => \b4_nUAi[81]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[82]\);
    
    \b6_OKctIF[193]\ : SLE
      port map(D => \b4_nUAi[309]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[310]\);
    
    \b6_OKctIF[136]\ : SLE
      port map(D => \b4_nUAi[366]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[367]\);
    
    \b6_OKctIF[120]\ : SLE
      port map(D => \b4_nUAi[382]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[383]\);
    
    \b6_OKctIF[423]\ : SLE
      port map(D => \b4_nUAi[79]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[80]\);
    
    \b6_OKctIF[258]\ : SLE
      port map(D => \b4_nUAi[244]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[245]\);
    
    \b6_OKctIF[90]\ : SLE
      port map(D => \b4_nUAi[412]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[413]\);
    
    \b6_OKctIF[247]\ : SLE
      port map(D => \b4_nUAi[255]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[256]\);
    
    \b6_OKctIF[455]\ : SLE
      port map(D => \b4_nUAi[47]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[48]\);
    
    \b6_OKctIF[192]\ : SLE
      port map(D => \b4_nUAi[310]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[311]\);
    
    \b6_OKctIF[123]\ : SLE
      port map(D => \b4_nUAi[379]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[380]\);
    
    \b6_OKctIF[108]\ : SLE
      port map(D => \b4_nUAi[394]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[395]\);
    
    \b6_OKctIF[365]\ : SLE
      port map(D => \b4_nUAi[137]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[138]\);
    
    \b6_OKctIF[265]\ : SLE
      port map(D => \b4_nUAi[237]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[238]\);
    
    \b6_OKctIF[188]\ : SLE
      port map(D => \b4_nUAi[314]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[315]\);
    
    \b6_OKctIF[367]\ : SLE
      port map(D => \b4_nUAi[135]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[136]\);
    
    \b6_OKctIF[48]\ : SLE
      port map(D => \b4_nUAi[454]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[455]\);
    
    \b6_OKctIF[45]\ : SLE
      port map(D => \b4_nUAi[457]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[458]\);
    
    \b6_OKctIF[231]\ : SLE
      port map(D => \b4_nUAi[271]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[272]\);
    
    \b6_OKctIF[214]\ : SLE
      port map(D => \b4_nUAi[288]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[289]\);
    
    \b6_OKctIF[459]\ : SLE
      port map(D => \b4_nUAi[43]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[44]\);
    
    \b6_OKctIF[122]\ : SLE
      port map(D => \b4_nUAi[380]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[381]\);
    
    \b6_OKctIF[82]\ : SLE
      port map(D => \b4_nUAi[420]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[421]\);
    
    \b6_OKctIF[218]\ : SLE
      port map(D => \b4_nUAi[284]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[285]\);
    
    \b6_OKctIF[89]\ : SLE
      port map(D => \b4_nUAi[413]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[414]\);
    
    \b6_OKctIF[415]\ : SLE
      port map(D => \b4_nUAi[87]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[88]\);
    
    \b6_OKctIF[451]\ : SLE
      port map(D => \b4_nUAi[51]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[52]\);
    
    \b6_OKctIF[478]\ : SLE
      port map(D => \b4_nUAi[24]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[25]\);
    
    \b6_OKctIF[203]\ : SLE
      port map(D => \b4_nUAi[299]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[300]\);
    
    \b6_OKctIF[150]\ : SLE
      port map(D => \b4_nUAi[352]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[353]\);
    
    \b6_OKctIF[283]\ : SLE
      port map(D => \b4_nUAi[219]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[220]\);
    
    \b6_OKctIF[242]\ : SLE
      port map(D => \b4_nUAi[260]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[261]\);
    
    \b6_OKctIF[453]\ : SLE
      port map(D => \b4_nUAi[49]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[50]\);
    
    \b6_OKctIF[303]\ : SLE
      port map(D => \b4_nUAi[199]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[200]\);
    
    \b6_OKctIF[383]\ : SLE
      port map(D => \b4_nUAi[119]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[120]\);
    
    \b6_OKctIF[419]\ : SLE
      port map(D => \b4_nUAi[83]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[84]\);
    
    \b6_OKctIF[306]\ : SLE
      port map(D => \b4_nUAi[196]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[197]\);
    
    \b6_OKctIF[153]\ : SLE
      port map(D => \b4_nUAi[349]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[350]\);
    
    \b6_OKctIF[101]\ : SLE
      port map(D => \b4_nUAi[401]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[402]\);
    
    \b6_OKctIF[386]\ : SLE
      port map(D => \b4_nUAi[116]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[117]\);
    
    \b6_OKctIF[181]\ : SLE
      port map(D => \b4_nUAi[321]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[322]\);
    
    \b6_OKctIF[80]\ : SLE
      port map(D => \b4_nUAi[422]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[423]\);
    
    \b6_OKctIF[494]\ : SLE
      port map(D => \b4_nUAi[8]\, CLK => IICE_comm2iice_4, EN => 
        \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[9]\);
    
    \b6_OKctIF[1]\ : SLE
      port map(D => \b4_nUAi[501]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[502]\);
    
    \b6_OKctIF[342]\ : SLE
      port map(D => \b4_nUAi[160]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[161]\);
    
    \b6_OKctIF[174]\ : SLE
      port map(D => \b4_nUAi[328]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[329]\);
    
    \b6_OKctIF[411]\ : SLE
      port map(D => \b4_nUAi[91]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[92]\);
    
    \b6_OKctIF[152]\ : SLE
      port map(D => \b4_nUAi[350]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[351]\);
    
    \b6_OKctIF[146]\ : SLE
      port map(D => \b4_nUAi[356]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[357]\);
    
    \b6_OKctIF[110]\ : SLE
      port map(D => \b4_nUAi[392]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[393]\);
    
    \b6_OKctIF[370]\ : SLE
      port map(D => \b4_nUAi[132]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[133]\);
    
    \b6_OKctIF[413]\ : SLE
      port map(D => \b4_nUAi[89]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[90]\);
    
    \b6_OKctIF[424]\ : SLE
      port map(D => \b4_nUAi[78]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[79]\);
    
    \b6_OKctIF[177]\ : SLE
      port map(D => \b4_nUAi[325]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[326]\);
    
    \b6_OKctIF[113]\ : SLE
      port map(D => \b4_nUAi[389]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[390]\);
    
    \b6_OKctIF[438]\ : SLE
      port map(D => \b4_nUAi[64]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[65]\);
    
    \b6_OKctIF[168]\ : SLE
      port map(D => \b4_nUAi[334]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[335]\);
    
    \b6_OKctIF[297]\ : SLE
      port map(D => \b4_nUAi[205]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[206]\);
    
    \b6_OKctIF[241]\ : SLE
      port map(D => \b4_nUAi[261]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[262]\);
    
    \b6_OKctIF[112]\ : SLE
      port map(D => \b4_nUAi[390]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[391]\);
    
    \b6_OKctIF[227]\ : SLE
      port map(D => \b4_nUAi[275]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[276]\);
    
    \b6_OKctIF[276]\ : SLE
      port map(D => \b4_nUAi[226]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[227]\);
    
    \b6_OKctIF[134]\ : SLE
      port map(D => \b4_nUAi[368]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[369]\);
    
    \b6_OKctIF[309]\ : SLE
      port map(D => \b4_nUAi[193]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[194]\);
    
    \b6_OKctIF[389]\ : SLE
      port map(D => \b4_nUAi[113]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[114]\);
    
    \b6_OKctIF[406]\ : SLE
      port map(D => \b4_nUAi[96]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[97]\);
    
    \b6_OKctIF[486]\ : SLE
      port map(D => \b4_nUAi[16]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[17]\);
    
    \b6_OKctIF[330]\ : SLE
      port map(D => \b4_nUAi[172]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[173]\);
    
    \b6_OKctIF[263]\ : SLE
      port map(D => \b4_nUAi[239]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[240]\);
    
    \b6_OKctIF[454]\ : SLE
      port map(D => \b4_nUAi[48]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[49]\);
    
    \b6_OKctIF[363]\ : SLE
      port map(D => \b4_nUAi[139]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[140]\);
    
    \b6_OKctIF[109]\ : SLE
      port map(D => \b4_nUAi[393]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[394]\);
    
    \b6_OKctIF[209]\ : SLE
      port map(D => \b4_nUAi[293]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[294]\);
    
    \b6_OKctIF[189]\ : SLE
      port map(D => \b4_nUAi[313]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[314]\);
    
    \b6_OKctIF[292]\ : SLE
      port map(D => \b4_nUAi[210]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[211]\);
    
    \b6_OKctIF[289]\ : SLE
      port map(D => \b4_nUAi[213]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[214]\);
    
    \b6_OKctIF[137]\ : SLE
      port map(D => \b4_nUAi[365]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[366]\);
    
    \b6_OKctIF[502]\ : SLE
      port map(D => \b4_nUAi[0]\, CLK => IICE_comm2iice_4, EN => 
        \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[1]\);
    
    \b6_OKctIF[366]\ : SLE
      port map(D => \b4_nUAi[136]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[137]\);
    
    \b6_OKctIF[161]\ : SLE
      port map(D => \b4_nUAi[341]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[342]\);
    
    \b6_OKctIF[8]\ : SLE
      port map(D => \b4_nUAi[494]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[495]\);
    
    \b6_OKctIF[200]\ : SLE
      port map(D => \b4_nUAi[302]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[303]\);
    
    \b6_OKctIF[371]\ : SLE
      port map(D => \b4_nUAi[131]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[132]\);
    
    \b6_OKctIF[280]\ : SLE
      port map(D => \b4_nUAi[222]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[223]\);
    
    \b6_OKctIF[105]\ : SLE
      port map(D => \b4_nUAi[397]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[398]\);
    
    \b6_OKctIF[185]\ : SLE
      port map(D => \b4_nUAi[317]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[318]\);
    
    \b6_OKctIF[392]\ : SLE
      port map(D => \b4_nUAi[110]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[111]\);
    
    \b6_OKctIF[378]\ : SLE
      port map(D => \b4_nUAi[124]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[125]\);
    
    \b6_OKctIF[222]\ : SLE
      port map(D => \b4_nUAi[280]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[281]\);
    
    \b6_OKctIF[414]\ : SLE
      port map(D => \b4_nUAi[88]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[89]\);
    
    \b6_OKctIF[257]\ : SLE
      port map(D => \b4_nUAi[245]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[246]\);
    
    \b6_OKctIF[236]\ : SLE
      port map(D => \b4_nUAi[266]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[267]\);
    
    \b6_OKctIF[196]\ : SLE
      port map(D => \b4_nUAi[306]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[307]\);
    
    \b6_OKctIF[448]\ : SLE
      port map(D => \b4_nUAi[54]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[55]\);
    
    \b6_OKctIF[470]\ : SLE
      port map(D => \b4_nUAi[32]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[33]\);
    
    \b6_OKctIF[322]\ : SLE
      port map(D => \b4_nUAi[180]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[181]\);
    
    \b6_OKctIF[28]\ : SLE
      port map(D => \b4_nUAi[474]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[475]\);
    
    \b6_OKctIF[25]\ : SLE
      port map(D => \b4_nUAi[477]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[478]\);
    
    \b6_OKctIF[126]\ : SLE
      port map(D => \b4_nUAi[376]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[377]\);
    
    \b6_OKctIF[291]\ : SLE
      port map(D => \b4_nUAi[211]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[212]\);
    
    \b6_OKctIF[217]\ : SLE
      port map(D => \b4_nUAi[285]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[286]\);
    
    \b6_OKctIF[144]\ : SLE
      port map(D => \b4_nUAi[358]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[359]\);
    
    \b6_OKctIF[44]\ : SLE
      port map(D => \b4_nUAi[458]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[459]\);
    
    \b6_OKctIF[369]\ : SLE
      port map(D => \b4_nUAi[133]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[134]\);
    
    \b6_OKctIF[331]\ : SLE
      port map(D => \b4_nUAi[171]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[172]\);
    
    \b6_OKctIF[252]\ : SLE
      port map(D => \b4_nUAi[250]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[251]\);
    
    \b6_OKctIF[466]\ : SLE
      port map(D => \b4_nUAi[36]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[37]\);
    
    \b6_OKctIF[340]\ : SLE
      port map(D => \b4_nUAi[162]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[163]\);
    
    \b6_OKctIF[338]\ : SLE
      port map(D => \b4_nUAi[164]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[165]\);
    
    \b6_OKctIF[221]\ : SLE
      port map(D => \b4_nUAi[281]\, CLK => IICE_comm2iice_4, EN
         => \b6_OKctIF4\, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b4_nUAi[282]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_39_0 is

    port( b4_nUAi           : in    std_logic_vector(386 downto 384);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_39_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_39_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_24, b3_P_F_6_2_24, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(386), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(384), D => b4_nUAi(385), Y => b3_P_F_6_2_24);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(385), D => b4_nUAi(384), Y => b3_P_F_6_0_24);
    
    b3_P_F_6_0_RNILUCN2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_24, B => b4_nUAi(385), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_24, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(386), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(384), D => b4_nUAi(385), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_93_0 is

    port( b4_nUAi           : in    std_logic_vector(224 downto 222);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_93_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_93_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_69, b3_P_F_6_2_69, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNIQ05M1 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_69, B => b4_nUAi(223), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_69, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(224), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(222), D => b4_nUAi(223), Y => b3_P_F_6_2_69);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(223), D => b4_nUAi(222), Y => b3_P_F_6_0_69);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(224), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(222), D => b4_nUAi(223), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_16_0 is

    port( b4_nUAi           : in    std_logic_vector(455 downto 453);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_16_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_16_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_31, b3_P_F_6_2_31, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(455), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(453), D => b4_nUAi(454), Y => b3_P_F_6_2_31);
    
    b3_P_F_6_0_RNIIHKM3 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_31, B => b4_nUAi(454), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_31, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(454), D => b4_nUAi(453), Y => b3_P_F_6_0_31);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(455), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(453), D => b4_nUAi(454), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_40_0 is

    port( b4_nUAi           : in    std_logic_vector(383 downto 381);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_40_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_40_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_107, b3_P_F_6_2_107, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(383), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(381), D => b4_nUAi(382), Y => b3_P_F_6_2_107);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNI4QO92 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_107, B => b4_nUAi(382), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_107, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(382), D => b4_nUAi(381), Y => b3_P_F_6_0_107);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(383), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(381), D => b4_nUAi(382), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_153_0 is

    port( b4_nUAi           : in    std_logic_vector(44 downto 42);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_153_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_153_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_157, b3_P_F_6_2_157, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(44), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(42), D => b4_nUAi(43), Y => b3_P_F_6_2_157);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(43), D => b4_nUAi(42), Y => b3_P_F_6_0_157);
    
    b3_P_F_6_0_RNI88S03 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_157, B => b4_nUAi(43), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_157, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(44), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(42), D => b4_nUAi(43), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_96_0 is

    port( b4_nUAi           : in    std_logic_vector(215 downto 213);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_96_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_96_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_72, b3_P_F_6_2_72, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(215), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(213), D => b4_nUAi(214), Y => b3_P_F_6_2_72);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNI777O1 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_72, B => b4_nUAi(214), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_72, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(214), D => b4_nUAi(213), Y => b3_P_F_6_0_72);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(215), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(213), D => b4_nUAi(214), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_156_0 is

    port( b4_nUAi           : in    std_logic_vector(35 downto 33);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_156_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_156_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_51, b3_P_F_6_2_51, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNIUOOB3 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_51, B => b4_nUAi(34), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_51, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(35), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(33), D => b4_nUAi(34), Y => b3_P_F_6_2_51);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(34), D => b4_nUAi(33), Y => b3_P_F_6_0_51);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(35), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(33), D => b4_nUAi(34), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_47_0 is

    port( b4_nUAi           : in    std_logic_vector(362 downto 360);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_47_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_47_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_114, b3_P_F_6_2_114, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(362), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(360), D => b4_nUAi(361), Y => b3_P_F_6_2_114);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNIQRPL2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_114, B => b4_nUAi(361), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_114, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(361), D => b4_nUAi(360), Y => b3_P_F_6_0_114);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(362), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(360), D => b4_nUAi(361), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_97_0 is

    port( b4_nUAi           : in    std_logic_vector(212 downto 210);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_97_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_97_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_73, b3_P_F_6_2_73, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(212), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(210), D => b4_nUAi(211), Y => b3_P_F_6_2_73);
    
    b3_P_F_6_0_RNIGVRA2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_73, B => b4_nUAi(211), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_73, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(211), D => b4_nUAi(210), Y => b3_P_F_6_0_73);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(212), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(210), D => b4_nUAi(211), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_157_0 is

    port( b4_nUAi           : in    std_logic_vector(32 downto 30);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_157_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_157_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_52, b3_P_F_6_2_52, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(32), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(30), D => b4_nUAi(31), Y => b3_P_F_6_2_52);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(31), D => b4_nUAi(30), Y => b3_P_F_6_0_52);
    
    b3_P_F_6_0_RNI7HDU2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_52, B => b4_nUAi(31), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_52, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(32), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(30), D => b4_nUAi(31), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_116_0 is

    port( b4_nUAi           : in    std_logic_vector(155 downto 153);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_116_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_116_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_60, b3_P_F_6_2_60, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(155), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(153), D => b4_nUAi(154), Y => b3_P_F_6_2_60);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNIQLTU2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_60, B => b4_nUAi(154), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_60, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(154), D => b4_nUAi(153), Y => b3_P_F_6_0_60);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(155), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(153), D => b4_nUAi(154), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b9_O2yyf_fG2_x_9_0 is

    port( b6_2ZTGIf           : in    std_logic_vector(95 downto 80);
          b13_CZS0wfY_d_FH9_0 : out   std_logic
        );

end b9_O2yyf_fG2_x_9_0;

architecture DEF_ARCH of b9_O2yyf_fG2_x_9_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \o_11\, \o_10\, \o_9\, \o_8\, GND_net_1, VCC_net_1
         : std_logic;

begin 


    o_10 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(90), B => b6_2ZTGIf(89), C => 
        b6_2ZTGIf(88), D => b6_2ZTGIf(87), Y => \o_10\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    o_9 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(92), B => b6_2ZTGIf(91), C => 
        b6_2ZTGIf(81), D => b6_2ZTGIf(80), Y => \o_9\);
    
    o : CFG4
      generic map(INIT => x"8000")

      port map(A => \o_11\, B => \o_10\, C => \o_9\, D => \o_8\, 
        Y => b13_CZS0wfY_d_FH9_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    o_8 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(94), B => b6_2ZTGIf(93), C => 
        b6_2ZTGIf(83), D => b6_2ZTGIf(82), Y => \o_8\);
    
    o_11 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(95), B => b6_2ZTGIf(86), C => 
        b6_2ZTGIf(85), D => b6_2ZTGIf(84), Y => \o_11\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b9_O2yyf_fG2_x_6_0 is

    port( b6_2ZTGIf           : in    std_logic_vector(143 downto 128);
          b13_CZS0wfY_d_FH9_0 : out   std_logic
        );

end b9_O2yyf_fG2_x_6_0;

architecture DEF_ARCH of b9_O2yyf_fG2_x_6_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \o_11\, \o_10\, \o_9\, \o_8\, GND_net_1, VCC_net_1
         : std_logic;

begin 


    o_10 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(138), B => b6_2ZTGIf(137), C => 
        b6_2ZTGIf(136), D => b6_2ZTGIf(135), Y => \o_10\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    o_9 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(140), B => b6_2ZTGIf(139), C => 
        b6_2ZTGIf(129), D => b6_2ZTGIf(128), Y => \o_9\);
    
    o : CFG4
      generic map(INIT => x"8000")

      port map(A => \o_11\, B => \o_10\, C => \o_9\, D => \o_8\, 
        Y => b13_CZS0wfY_d_FH9_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    o_8 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(142), B => b6_2ZTGIf(141), C => 
        b6_2ZTGIf(131), D => b6_2ZTGIf(130), Y => \o_8\);
    
    o_11 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(143), B => b6_2ZTGIf(134), C => 
        b6_2ZTGIf(133), D => b6_2ZTGIf(132), Y => \o_11\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b9_O2yyf_fG2_x_5_0 is

    port( b6_2ZTGIf           : in    std_logic_vector(159 downto 144);
          b13_CZS0wfY_d_FH9_0 : out   std_logic
        );

end b9_O2yyf_fG2_x_5_0;

architecture DEF_ARCH of b9_O2yyf_fG2_x_5_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \o_11\, \o_10\, \o_9\, \o_8\, GND_net_1, VCC_net_1
         : std_logic;

begin 


    o_10 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(154), B => b6_2ZTGIf(153), C => 
        b6_2ZTGIf(152), D => b6_2ZTGIf(151), Y => \o_10\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    o_9 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(156), B => b6_2ZTGIf(155), C => 
        b6_2ZTGIf(145), D => b6_2ZTGIf(144), Y => \o_9\);
    
    o : CFG4
      generic map(INIT => x"8000")

      port map(A => \o_11\, B => \o_10\, C => \o_9\, D => \o_8\, 
        Y => b13_CZS0wfY_d_FH9_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    o_8 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(158), B => b6_2ZTGIf(157), C => 
        b6_2ZTGIf(147), D => b6_2ZTGIf(146), Y => \o_8\);
    
    o_11 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(159), B => b6_2ZTGIf(150), C => 
        b6_2ZTGIf(149), D => b6_2ZTGIf(148), Y => \o_11\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b9_O2yyf_fG2_x_14_0 is

    port( b6_2ZTGIf           : in    std_logic_vector(15 downto 0);
          b13_CZS0wfY_d_FH9_0 : out   std_logic
        );

end b9_O2yyf_fG2_x_14_0;

architecture DEF_ARCH of b9_O2yyf_fG2_x_14_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \o_11\, \o_10\, \o_9\, \o_8\, GND_net_1, VCC_net_1
         : std_logic;

begin 


    o_10 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(10), B => b6_2ZTGIf(9), C => 
        b6_2ZTGIf(8), D => b6_2ZTGIf(7), Y => \o_10\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    o_9 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(12), B => b6_2ZTGIf(11), C => 
        b6_2ZTGIf(1), D => b6_2ZTGIf(0), Y => \o_9\);
    
    o : CFG4
      generic map(INIT => x"8000")

      port map(A => \o_11\, B => \o_10\, C => \o_9\, D => \o_8\, 
        Y => b13_CZS0wfY_d_FH9_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    o_8 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(14), B => b6_2ZTGIf(13), C => 
        b6_2ZTGIf(3), D => b6_2ZTGIf(2), Y => \o_8\);
    
    o_11 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(15), B => b6_2ZTGIf(6), C => 
        b6_2ZTGIf(5), D => b6_2ZTGIf(4), Y => \o_11\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b9_O2yyf_fG2_x_10_0 is

    port( b6_2ZTGIf           : in    std_logic_vector(79 downto 64);
          b13_CZS0wfY_d_FH9_0 : out   std_logic
        );

end b9_O2yyf_fG2_x_10_0;

architecture DEF_ARCH of b9_O2yyf_fG2_x_10_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \o_11\, \o_10\, \o_9\, \o_8\, GND_net_1, VCC_net_1
         : std_logic;

begin 


    o_10 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(74), B => b6_2ZTGIf(73), C => 
        b6_2ZTGIf(72), D => b6_2ZTGIf(71), Y => \o_10\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    o_9 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(76), B => b6_2ZTGIf(75), C => 
        b6_2ZTGIf(65), D => b6_2ZTGIf(64), Y => \o_9\);
    
    o : CFG4
      generic map(INIT => x"8000")

      port map(A => \o_11\, B => \o_10\, C => \o_9\, D => \o_8\, 
        Y => b13_CZS0wfY_d_FH9_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    o_8 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(78), B => b6_2ZTGIf(77), C => 
        b6_2ZTGIf(67), D => b6_2ZTGIf(66), Y => \o_8\);
    
    o_11 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(79), B => b6_2ZTGIf(70), C => 
        b6_2ZTGIf(69), D => b6_2ZTGIf(68), Y => \o_11\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b9_O2yyf_fG2_x_11_0 is

    port( b6_2ZTGIf           : in    std_logic_vector(63 downto 48);
          b13_CZS0wfY_d_FH9_0 : out   std_logic
        );

end b9_O2yyf_fG2_x_11_0;

architecture DEF_ARCH of b9_O2yyf_fG2_x_11_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \o_11\, \o_10\, \o_9\, \o_8\, GND_net_1, VCC_net_1
         : std_logic;

begin 


    o_10 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(58), B => b6_2ZTGIf(57), C => 
        b6_2ZTGIf(56), D => b6_2ZTGIf(55), Y => \o_10\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    o_9 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(60), B => b6_2ZTGIf(59), C => 
        b6_2ZTGIf(49), D => b6_2ZTGIf(48), Y => \o_9\);
    
    o : CFG4
      generic map(INIT => x"8000")

      port map(A => \o_11\, B => \o_10\, C => \o_9\, D => \o_8\, 
        Y => b13_CZS0wfY_d_FH9_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    o_8 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(62), B => b6_2ZTGIf(61), C => 
        b6_2ZTGIf(51), D => b6_2ZTGIf(50), Y => \o_8\);
    
    o_11 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(63), B => b6_2ZTGIf(54), C => 
        b6_2ZTGIf(53), D => b6_2ZTGIf(52), Y => \o_11\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b9_O2yyf_fG2_x_12_0 is

    port( b6_2ZTGIf           : in    std_logic_vector(47 downto 32);
          b13_CZS0wfY_d_FH9_0 : out   std_logic
        );

end b9_O2yyf_fG2_x_12_0;

architecture DEF_ARCH of b9_O2yyf_fG2_x_12_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \o_11\, \o_10\, \o_9\, \o_8\, GND_net_1, VCC_net_1
         : std_logic;

begin 


    o_10 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(42), B => b6_2ZTGIf(41), C => 
        b6_2ZTGIf(40), D => b6_2ZTGIf(39), Y => \o_10\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    o_9 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(44), B => b6_2ZTGIf(43), C => 
        b6_2ZTGIf(33), D => b6_2ZTGIf(32), Y => \o_9\);
    
    o : CFG4
      generic map(INIT => x"8000")

      port map(A => \o_11\, B => \o_10\, C => \o_9\, D => \o_8\, 
        Y => b13_CZS0wfY_d_FH9_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    o_8 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(46), B => b6_2ZTGIf(45), C => 
        b6_2ZTGIf(35), D => b6_2ZTGIf(34), Y => \o_8\);
    
    o_11 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(47), B => b6_2ZTGIf(38), C => 
        b6_2ZTGIf(37), D => b6_2ZTGIf(36), Y => \o_11\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b9_O2yyf_fG2_x_7_0 is

    port( b6_2ZTGIf           : in    std_logic_vector(127 downto 112);
          b13_CZS0wfY_d_FH9_0 : out   std_logic
        );

end b9_O2yyf_fG2_x_7_0;

architecture DEF_ARCH of b9_O2yyf_fG2_x_7_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \o_11\, \o_10\, \o_9\, \o_8\, GND_net_1, VCC_net_1
         : std_logic;

begin 


    o_10 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(122), B => b6_2ZTGIf(121), C => 
        b6_2ZTGIf(120), D => b6_2ZTGIf(119), Y => \o_10\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    o_9 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(124), B => b6_2ZTGIf(123), C => 
        b6_2ZTGIf(113), D => b6_2ZTGIf(112), Y => \o_9\);
    
    o : CFG4
      generic map(INIT => x"8000")

      port map(A => \o_11\, B => \o_10\, C => \o_9\, D => \o_8\, 
        Y => b13_CZS0wfY_d_FH9_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    o_8 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(126), B => b6_2ZTGIf(125), C => 
        b6_2ZTGIf(115), D => b6_2ZTGIf(114), Y => \o_8\);
    
    o_11 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(127), B => b6_2ZTGIf(118), C => 
        b6_2ZTGIf(117), D => b6_2ZTGIf(116), Y => \o_11\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b9_O2yyf_fG2_x_4_0 is

    port( b6_2ZTGIf           : in    std_logic_vector(167 downto 160);
          b13_CZS0wfY_d_FH9_0 : out   std_logic
        );

end b9_O2yyf_fG2_x_4_0;

architecture DEF_ARCH of b9_O2yyf_fG2_x_4_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \o_3\, \o_4\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    o_4 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(163), B => b6_2ZTGIf(162), C => 
        b6_2ZTGIf(161), D => b6_2ZTGIf(160), Y => \o_4\);
    
    o_3 : CFG2
      generic map(INIT => x"8")

      port map(A => b6_2ZTGIf(164), B => b6_2ZTGIf(165), Y => 
        \o_3\);
    
    o : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(166), B => b6_2ZTGIf(167), C => 
        \o_4\, D => \o_3\, Y => b13_CZS0wfY_d_FH9_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b9_O2yyf_fG2_x_0_0 is

    port( b14_CZS0wfY_d_FH9m : in    std_logic_vector(10 downto 0);
          b10_nYBzIXrKbK_0   : out   std_logic
        );

end b9_O2yyf_fG2_x_0_0;

architecture DEF_ARCH of b9_O2yyf_fG2_x_0_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \o_4\, \o_6\, \o_8\, GND_net_1, VCC_net_1
         : std_logic;

begin 


    o_6 : CFG4
      generic map(INIT => x"8000")

      port map(A => b14_CZS0wfY_d_FH9m(4), B => 
        b14_CZS0wfY_d_FH9m(3), C => b14_CZS0wfY_d_FH9m(2), D => 
        b14_CZS0wfY_d_FH9m(1), Y => \o_6\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    o_4 : CFG2
      generic map(INIT => x"8")

      port map(A => b14_CZS0wfY_d_FH9m(8), B => 
        b14_CZS0wfY_d_FH9m(10), Y => \o_4\);
    
    o : CFG4
      generic map(INIT => x"8000")

      port map(A => b14_CZS0wfY_d_FH9m(0), B => 
        b14_CZS0wfY_d_FH9m(9), C => \o_8\, D => \o_4\, Y => 
        b10_nYBzIXrKbK_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    o_8 : CFG4
      generic map(INIT => x"8000")

      port map(A => b14_CZS0wfY_d_FH9m(5), B => \o_6\, C => 
        b14_CZS0wfY_d_FH9m(7), D => b14_CZS0wfY_d_FH9m(6), Y => 
        \o_8\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b9_O2yyf_fG2_x_13_0 is

    port( b6_2ZTGIf           : in    std_logic_vector(31 downto 16);
          b13_CZS0wfY_d_FH9_0 : out   std_logic
        );

end b9_O2yyf_fG2_x_13_0;

architecture DEF_ARCH of b9_O2yyf_fG2_x_13_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \o_11\, \o_10\, \o_9\, \o_8\, GND_net_1, VCC_net_1
         : std_logic;

begin 


    o_10 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(26), B => b6_2ZTGIf(25), C => 
        b6_2ZTGIf(24), D => b6_2ZTGIf(23), Y => \o_10\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    o_9 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(28), B => b6_2ZTGIf(27), C => 
        b6_2ZTGIf(17), D => b6_2ZTGIf(16), Y => \o_9\);
    
    o : CFG4
      generic map(INIT => x"8000")

      port map(A => \o_11\, B => \o_10\, C => \o_9\, D => \o_8\, 
        Y => b13_CZS0wfY_d_FH9_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    o_8 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(30), B => b6_2ZTGIf(29), C => 
        b6_2ZTGIf(19), D => b6_2ZTGIf(18), Y => \o_8\);
    
    o_11 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(31), B => b6_2ZTGIf(22), C => 
        b6_2ZTGIf(21), D => b6_2ZTGIf(20), Y => \o_11\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b9_O2yyf_fG2_x_8_0 is

    port( b6_2ZTGIf           : in    std_logic_vector(111 downto 96);
          b13_CZS0wfY_d_FH9_0 : out   std_logic
        );

end b9_O2yyf_fG2_x_8_0;

architecture DEF_ARCH of b9_O2yyf_fG2_x_8_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \o_11\, \o_10\, \o_9\, \o_8\, GND_net_1, VCC_net_1
         : std_logic;

begin 


    o_10 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(106), B => b6_2ZTGIf(105), C => 
        b6_2ZTGIf(104), D => b6_2ZTGIf(103), Y => \o_10\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    o_9 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(108), B => b6_2ZTGIf(107), C => 
        b6_2ZTGIf(97), D => b6_2ZTGIf(96), Y => \o_9\);
    
    o : CFG4
      generic map(INIT => x"8000")

      port map(A => \o_11\, B => \o_10\, C => \o_9\, D => \o_8\, 
        Y => b13_CZS0wfY_d_FH9_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    o_8 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(110), B => b6_2ZTGIf(109), C => 
        b6_2ZTGIf(99), D => b6_2ZTGIf(98), Y => \o_8\);
    
    o_11 : CFG4
      generic map(INIT => x"8000")

      port map(A => b6_2ZTGIf(111), B => b6_2ZTGIf(102), C => 
        b6_2ZTGIf(101), D => b6_2ZTGIf(100), Y => \o_11\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b16_CRGcTCua_eH4_uaL_x_0 is

    port( b6_2ZTGIf           : in    std_logic_vector(167 downto 0);
          b10_nYBzIXrKbK_0    : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic
        );

end b16_CRGcTCua_eH4_uaL_x_0;

architecture DEF_ARCH of b16_CRGcTCua_eH4_uaL_x_0 is 

  component b9_O2yyf_fG2_x_9_0
    port( b6_2ZTGIf           : in    std_logic_vector(95 downto 80) := (others => 'U');
          b13_CZS0wfY_d_FH9_0 : out   std_logic
        );
  end component;

  component b9_O2yyf_fG2_x_6_0
    port( b6_2ZTGIf           : in    std_logic_vector(143 downto 128) := (others => 'U');
          b13_CZS0wfY_d_FH9_0 : out   std_logic
        );
  end component;

  component b9_O2yyf_fG2_x_5_0
    port( b6_2ZTGIf           : in    std_logic_vector(159 downto 144) := (others => 'U');
          b13_CZS0wfY_d_FH9_0 : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component b9_O2yyf_fG2_x_14_0
    port( b6_2ZTGIf           : in    std_logic_vector(15 downto 0) := (others => 'U');
          b13_CZS0wfY_d_FH9_0 : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component b9_O2yyf_fG2_x_10_0
    port( b6_2ZTGIf           : in    std_logic_vector(79 downto 64) := (others => 'U');
          b13_CZS0wfY_d_FH9_0 : out   std_logic
        );
  end component;

  component b9_O2yyf_fG2_x_11_0
    port( b6_2ZTGIf           : in    std_logic_vector(63 downto 48) := (others => 'U');
          b13_CZS0wfY_d_FH9_0 : out   std_logic
        );
  end component;

  component b9_O2yyf_fG2_x_12_0
    port( b6_2ZTGIf           : in    std_logic_vector(47 downto 32) := (others => 'U');
          b13_CZS0wfY_d_FH9_0 : out   std_logic
        );
  end component;

  component b9_O2yyf_fG2_x_7_0
    port( b6_2ZTGIf           : in    std_logic_vector(127 downto 112) := (others => 'U');
          b13_CZS0wfY_d_FH9_0 : out   std_logic
        );
  end component;

  component b9_O2yyf_fG2_x_4_0
    port( b6_2ZTGIf           : in    std_logic_vector(167 downto 160) := (others => 'U');
          b13_CZS0wfY_d_FH9_0 : out   std_logic
        );
  end component;

  component b9_O2yyf_fG2_x_0_0
    port( b14_CZS0wfY_d_FH9m : in    std_logic_vector(10 downto 0) := (others => 'U');
          b10_nYBzIXrKbK_0   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component b9_O2yyf_fG2_x_13_0
    port( b6_2ZTGIf           : in    std_logic_vector(31 downto 16) := (others => 'U');
          b13_CZS0wfY_d_FH9_0 : out   std_logic
        );
  end component;

  component b9_O2yyf_fG2_x_8_0
    port( b6_2ZTGIf           : in    std_logic_vector(111 downto 96) := (others => 'U');
          b13_CZS0wfY_d_FH9_0 : out   std_logic
        );
  end component;

    signal \b14_CZS0wfY_d_FH9m[10]_net_1\, VCC_net_1, 
        \b13_CZS0wfY_d_FH9[10]\, GND_net_1, 
        \b14_CZS0wfY_d_FH9m[9]_net_1\, \b13_CZS0wfY_d_FH9[9]\, 
        \b14_CZS0wfY_d_FH9m[8]_net_1\, \b13_CZS0wfY_d_FH9[8]\, 
        \b14_CZS0wfY_d_FH9m[7]_net_1\, \b13_CZS0wfY_d_FH9[7]\, 
        \b14_CZS0wfY_d_FH9m[6]_net_1\, \b13_CZS0wfY_d_FH9[6]\, 
        \b14_CZS0wfY_d_FH9m[5]_net_1\, \b13_CZS0wfY_d_FH9[5]\, 
        \b14_CZS0wfY_d_FH9m[4]_net_1\, \b13_CZS0wfY_d_FH9[4]\, 
        \b14_CZS0wfY_d_FH9m[3]_net_1\, \b13_CZS0wfY_d_FH9[3]\, 
        \b14_CZS0wfY_d_FH9m[2]_net_1\, \b13_CZS0wfY_d_FH9[2]\, 
        \b14_CZS0wfY_d_FH9m[1]_net_1\, \b13_CZS0wfY_d_FH9[1]\, 
        \b14_CZS0wfY_d_FH9m[0]_net_1\, \b13_CZS0wfY_d_FH9[0]\
         : std_logic;

    for all : b9_O2yyf_fG2_x_9_0
	Use entity work.b9_O2yyf_fG2_x_9_0(DEF_ARCH);
    for all : b9_O2yyf_fG2_x_6_0
	Use entity work.b9_O2yyf_fG2_x_6_0(DEF_ARCH);
    for all : b9_O2yyf_fG2_x_5_0
	Use entity work.b9_O2yyf_fG2_x_5_0(DEF_ARCH);
    for all : b9_O2yyf_fG2_x_14_0
	Use entity work.b9_O2yyf_fG2_x_14_0(DEF_ARCH);
    for all : b9_O2yyf_fG2_x_10_0
	Use entity work.b9_O2yyf_fG2_x_10_0(DEF_ARCH);
    for all : b9_O2yyf_fG2_x_11_0
	Use entity work.b9_O2yyf_fG2_x_11_0(DEF_ARCH);
    for all : b9_O2yyf_fG2_x_12_0
	Use entity work.b9_O2yyf_fG2_x_12_0(DEF_ARCH);
    for all : b9_O2yyf_fG2_x_7_0
	Use entity work.b9_O2yyf_fG2_x_7_0(DEF_ARCH);
    for all : b9_O2yyf_fG2_x_4_0
	Use entity work.b9_O2yyf_fG2_x_4_0(DEF_ARCH);
    for all : b9_O2yyf_fG2_x_0_0
	Use entity work.b9_O2yyf_fG2_x_0_0(DEF_ARCH);
    for all : b9_O2yyf_fG2_x_13_0
	Use entity work.b9_O2yyf_fG2_x_13_0(DEF_ARCH);
    for all : b9_O2yyf_fG2_x_8_0
	Use entity work.b9_O2yyf_fG2_x_8_0(DEF_ARCH);
begin 


    b27_O2yyf_fG2_MiQA1E6_r_lnxob_c : b9_O2yyf_fG2_x_9_0
      port map(b6_2ZTGIf(95) => b6_2ZTGIf(95), b6_2ZTGIf(94) => 
        b6_2ZTGIf(94), b6_2ZTGIf(93) => b6_2ZTGIf(93), 
        b6_2ZTGIf(92) => b6_2ZTGIf(92), b6_2ZTGIf(91) => 
        b6_2ZTGIf(91), b6_2ZTGIf(90) => b6_2ZTGIf(90), 
        b6_2ZTGIf(89) => b6_2ZTGIf(89), b6_2ZTGIf(88) => 
        b6_2ZTGIf(88), b6_2ZTGIf(87) => b6_2ZTGIf(87), 
        b6_2ZTGIf(86) => b6_2ZTGIf(86), b6_2ZTGIf(85) => 
        b6_2ZTGIf(85), b6_2ZTGIf(84) => b6_2ZTGIf(84), 
        b6_2ZTGIf(83) => b6_2ZTGIf(83), b6_2ZTGIf(82) => 
        b6_2ZTGIf(82), b6_2ZTGIf(81) => b6_2ZTGIf(81), 
        b6_2ZTGIf(80) => b6_2ZTGIf(80), b13_CZS0wfY_d_FH9_0 => 
        \b13_CZS0wfY_d_FH9[5]\);
    
    b27_O2yyf_fG2_MiQA1E6_r_lnxob_F : b9_O2yyf_fG2_x_6_0
      port map(b6_2ZTGIf(143) => b6_2ZTGIf(143), b6_2ZTGIf(142)
         => b6_2ZTGIf(142), b6_2ZTGIf(141) => b6_2ZTGIf(141), 
        b6_2ZTGIf(140) => b6_2ZTGIf(140), b6_2ZTGIf(139) => 
        b6_2ZTGIf(139), b6_2ZTGIf(138) => b6_2ZTGIf(138), 
        b6_2ZTGIf(137) => b6_2ZTGIf(137), b6_2ZTGIf(136) => 
        b6_2ZTGIf(136), b6_2ZTGIf(135) => b6_2ZTGIf(135), 
        b6_2ZTGIf(134) => b6_2ZTGIf(134), b6_2ZTGIf(133) => 
        b6_2ZTGIf(133), b6_2ZTGIf(132) => b6_2ZTGIf(132), 
        b6_2ZTGIf(131) => b6_2ZTGIf(131), b6_2ZTGIf(130) => 
        b6_2ZTGIf(130), b6_2ZTGIf(129) => b6_2ZTGIf(129), 
        b6_2ZTGIf(128) => b6_2ZTGIf(128), b13_CZS0wfY_d_FH9_0 => 
        \b13_CZS0wfY_d_FH9[8]\);
    
    b27_O2yyf_fG2_MiQA1E6_r_lnxob_d : b9_O2yyf_fG2_x_5_0
      port map(b6_2ZTGIf(159) => b6_2ZTGIf(159), b6_2ZTGIf(158)
         => b6_2ZTGIf(158), b6_2ZTGIf(157) => b6_2ZTGIf(157), 
        b6_2ZTGIf(156) => b6_2ZTGIf(156), b6_2ZTGIf(155) => 
        b6_2ZTGIf(155), b6_2ZTGIf(154) => b6_2ZTGIf(154), 
        b6_2ZTGIf(153) => b6_2ZTGIf(153), b6_2ZTGIf(152) => 
        b6_2ZTGIf(152), b6_2ZTGIf(151) => b6_2ZTGIf(151), 
        b6_2ZTGIf(150) => b6_2ZTGIf(150), b6_2ZTGIf(149) => 
        b6_2ZTGIf(149), b6_2ZTGIf(148) => b6_2ZTGIf(148), 
        b6_2ZTGIf(147) => b6_2ZTGIf(147), b6_2ZTGIf(146) => 
        b6_2ZTGIf(146), b6_2ZTGIf(145) => b6_2ZTGIf(145), 
        b6_2ZTGIf(144) => b6_2ZTGIf(144), b13_CZS0wfY_d_FH9_0 => 
        \b13_CZS0wfY_d_FH9[9]\);
    
    \b14_CZS0wfY_d_FH9m[4]\ : SLE
      port map(D => \b13_CZS0wfY_d_FH9[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b14_CZS0wfY_d_FH9m[4]_net_1\);
    
    b27_O2yyf_fG2_MiQA1E6_r_lnxob_9 : b9_O2yyf_fG2_x_14_0
      port map(b6_2ZTGIf(15) => b6_2ZTGIf(15), b6_2ZTGIf(14) => 
        b6_2ZTGIf(14), b6_2ZTGIf(13) => b6_2ZTGIf(13), 
        b6_2ZTGIf(12) => b6_2ZTGIf(12), b6_2ZTGIf(11) => 
        b6_2ZTGIf(11), b6_2ZTGIf(10) => b6_2ZTGIf(10), 
        b6_2ZTGIf(9) => b6_2ZTGIf(9), b6_2ZTGIf(8) => 
        b6_2ZTGIf(8), b6_2ZTGIf(7) => b6_2ZTGIf(7), b6_2ZTGIf(6)
         => b6_2ZTGIf(6), b6_2ZTGIf(5) => b6_2ZTGIf(5), 
        b6_2ZTGIf(4) => b6_2ZTGIf(4), b6_2ZTGIf(3) => 
        b6_2ZTGIf(3), b6_2ZTGIf(2) => b6_2ZTGIf(2), b6_2ZTGIf(1)
         => b6_2ZTGIf(1), b6_2ZTGIf(0) => b6_2ZTGIf(0), 
        b13_CZS0wfY_d_FH9_0 => \b13_CZS0wfY_d_FH9[0]\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b27_O2yyf_fG2_MiQA1E6_r_lnxob_8 : b9_O2yyf_fG2_x_10_0
      port map(b6_2ZTGIf(79) => b6_2ZTGIf(79), b6_2ZTGIf(78) => 
        b6_2ZTGIf(78), b6_2ZTGIf(77) => b6_2ZTGIf(77), 
        b6_2ZTGIf(76) => b6_2ZTGIf(76), b6_2ZTGIf(75) => 
        b6_2ZTGIf(75), b6_2ZTGIf(74) => b6_2ZTGIf(74), 
        b6_2ZTGIf(73) => b6_2ZTGIf(73), b6_2ZTGIf(72) => 
        b6_2ZTGIf(72), b6_2ZTGIf(71) => b6_2ZTGIf(71), 
        b6_2ZTGIf(70) => b6_2ZTGIf(70), b6_2ZTGIf(69) => 
        b6_2ZTGIf(69), b6_2ZTGIf(68) => b6_2ZTGIf(68), 
        b6_2ZTGIf(67) => b6_2ZTGIf(67), b6_2ZTGIf(66) => 
        b6_2ZTGIf(66), b6_2ZTGIf(65) => b6_2ZTGIf(65), 
        b6_2ZTGIf(64) => b6_2ZTGIf(64), b13_CZS0wfY_d_FH9_0 => 
        \b13_CZS0wfY_d_FH9[4]\);
    
    b27_O2yyf_fG2_MiQA1E6_r_lnxob_I : b9_O2yyf_fG2_x_11_0
      port map(b6_2ZTGIf(63) => b6_2ZTGIf(63), b6_2ZTGIf(62) => 
        b6_2ZTGIf(62), b6_2ZTGIf(61) => b6_2ZTGIf(61), 
        b6_2ZTGIf(60) => b6_2ZTGIf(60), b6_2ZTGIf(59) => 
        b6_2ZTGIf(59), b6_2ZTGIf(58) => b6_2ZTGIf(58), 
        b6_2ZTGIf(57) => b6_2ZTGIf(57), b6_2ZTGIf(56) => 
        b6_2ZTGIf(56), b6_2ZTGIf(55) => b6_2ZTGIf(55), 
        b6_2ZTGIf(54) => b6_2ZTGIf(54), b6_2ZTGIf(53) => 
        b6_2ZTGIf(53), b6_2ZTGIf(52) => b6_2ZTGIf(52), 
        b6_2ZTGIf(51) => b6_2ZTGIf(51), b6_2ZTGIf(50) => 
        b6_2ZTGIf(50), b6_2ZTGIf(49) => b6_2ZTGIf(49), 
        b6_2ZTGIf(48) => b6_2ZTGIf(48), b13_CZS0wfY_d_FH9_0 => 
        \b13_CZS0wfY_d_FH9[3]\);
    
    \b14_CZS0wfY_d_FH9m[3]\ : SLE
      port map(D => \b13_CZS0wfY_d_FH9[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b14_CZS0wfY_d_FH9m[3]_net_1\);
    
    \b14_CZS0wfY_d_FH9m[1]\ : SLE
      port map(D => \b13_CZS0wfY_d_FH9[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b14_CZS0wfY_d_FH9m[1]_net_1\);
    
    \b14_CZS0wfY_d_FH9m[5]\ : SLE
      port map(D => \b13_CZS0wfY_d_FH9[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b14_CZS0wfY_d_FH9m[5]_net_1\);
    
    b27_O2yyf_fG2_MiQA1E6_r_lnxob_0 : b9_O2yyf_fG2_x_12_0
      port map(b6_2ZTGIf(47) => b6_2ZTGIf(47), b6_2ZTGIf(46) => 
        b6_2ZTGIf(46), b6_2ZTGIf(45) => b6_2ZTGIf(45), 
        b6_2ZTGIf(44) => b6_2ZTGIf(44), b6_2ZTGIf(43) => 
        b6_2ZTGIf(43), b6_2ZTGIf(42) => b6_2ZTGIf(42), 
        b6_2ZTGIf(41) => b6_2ZTGIf(41), b6_2ZTGIf(40) => 
        b6_2ZTGIf(40), b6_2ZTGIf(39) => b6_2ZTGIf(39), 
        b6_2ZTGIf(38) => b6_2ZTGIf(38), b6_2ZTGIf(37) => 
        b6_2ZTGIf(37), b6_2ZTGIf(36) => b6_2ZTGIf(36), 
        b6_2ZTGIf(35) => b6_2ZTGIf(35), b6_2ZTGIf(34) => 
        b6_2ZTGIf(34), b6_2ZTGIf(33) => b6_2ZTGIf(33), 
        b6_2ZTGIf(32) => b6_2ZTGIf(32), b13_CZS0wfY_d_FH9_0 => 
        \b13_CZS0wfY_d_FH9[2]\);
    
    \b14_CZS0wfY_d_FH9m[6]\ : SLE
      port map(D => \b13_CZS0wfY_d_FH9[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b14_CZS0wfY_d_FH9m[6]_net_1\);
    
    b27_O2yyf_fG2_MiQA1E6_r_lnxob_1 : b9_O2yyf_fG2_x_7_0
      port map(b6_2ZTGIf(127) => b6_2ZTGIf(127), b6_2ZTGIf(126)
         => b6_2ZTGIf(126), b6_2ZTGIf(125) => b6_2ZTGIf(125), 
        b6_2ZTGIf(124) => b6_2ZTGIf(124), b6_2ZTGIf(123) => 
        b6_2ZTGIf(123), b6_2ZTGIf(122) => b6_2ZTGIf(122), 
        b6_2ZTGIf(121) => b6_2ZTGIf(121), b6_2ZTGIf(120) => 
        b6_2ZTGIf(120), b6_2ZTGIf(119) => b6_2ZTGIf(119), 
        b6_2ZTGIf(118) => b6_2ZTGIf(118), b6_2ZTGIf(117) => 
        b6_2ZTGIf(117), b6_2ZTGIf(116) => b6_2ZTGIf(116), 
        b6_2ZTGIf(115) => b6_2ZTGIf(115), b6_2ZTGIf(114) => 
        b6_2ZTGIf(114), b6_2ZTGIf(113) => b6_2ZTGIf(113), 
        b6_2ZTGIf(112) => b6_2ZTGIf(112), b13_CZS0wfY_d_FH9_0 => 
        \b13_CZS0wfY_d_FH9[7]\);
    
    \b14_CZS0wfY_d_FH9m[9]\ : SLE
      port map(D => \b13_CZS0wfY_d_FH9[9]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b14_CZS0wfY_d_FH9m[9]_net_1\);
    
    \b14_CZS0wfY_d_FH9m[7]\ : SLE
      port map(D => \b13_CZS0wfY_d_FH9[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b14_CZS0wfY_d_FH9m[7]_net_1\);
    
    b28_O2yyf_fG2_MiQA1E6_r_lnxob_a6 : b9_O2yyf_fG2_x_4_0
      port map(b6_2ZTGIf(167) => b6_2ZTGIf(167), b6_2ZTGIf(166)
         => b6_2ZTGIf(166), b6_2ZTGIf(165) => b6_2ZTGIf(165), 
        b6_2ZTGIf(164) => b6_2ZTGIf(164), b6_2ZTGIf(163) => 
        b6_2ZTGIf(163), b6_2ZTGIf(162) => b6_2ZTGIf(162), 
        b6_2ZTGIf(161) => b6_2ZTGIf(161), b6_2ZTGIf(160) => 
        b6_2ZTGIf(160), b13_CZS0wfY_d_FH9_0 => 
        \b13_CZS0wfY_d_FH9[10]\);
    
    b25_O2yyf_fG2_MiQA1E6_Z_lnxob : b9_O2yyf_fG2_x_0_0
      port map(b14_CZS0wfY_d_FH9m(10) => 
        \b14_CZS0wfY_d_FH9m[10]_net_1\, b14_CZS0wfY_d_FH9m(9) => 
        \b14_CZS0wfY_d_FH9m[9]_net_1\, b14_CZS0wfY_d_FH9m(8) => 
        \b14_CZS0wfY_d_FH9m[8]_net_1\, b14_CZS0wfY_d_FH9m(7) => 
        \b14_CZS0wfY_d_FH9m[7]_net_1\, b14_CZS0wfY_d_FH9m(6) => 
        \b14_CZS0wfY_d_FH9m[6]_net_1\, b14_CZS0wfY_d_FH9m(5) => 
        \b14_CZS0wfY_d_FH9m[5]_net_1\, b14_CZS0wfY_d_FH9m(4) => 
        \b14_CZS0wfY_d_FH9m[4]_net_1\, b14_CZS0wfY_d_FH9m(3) => 
        \b14_CZS0wfY_d_FH9m[3]_net_1\, b14_CZS0wfY_d_FH9m(2) => 
        \b14_CZS0wfY_d_FH9m[2]_net_1\, b14_CZS0wfY_d_FH9m(1) => 
        \b14_CZS0wfY_d_FH9m[1]_net_1\, b14_CZS0wfY_d_FH9m(0) => 
        \b14_CZS0wfY_d_FH9m[0]_net_1\, b10_nYBzIXrKbK_0 => 
        b10_nYBzIXrKbK_0);
    
    \b14_CZS0wfY_d_FH9m[2]\ : SLE
      port map(D => \b13_CZS0wfY_d_FH9[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b14_CZS0wfY_d_FH9m[2]_net_1\);
    
    \b14_CZS0wfY_d_FH9m[0]\ : SLE
      port map(D => \b13_CZS0wfY_d_FH9[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b14_CZS0wfY_d_FH9m[0]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b27_O2yyf_fG2_MiQA1E6_r_lnxob_a : b9_O2yyf_fG2_x_13_0
      port map(b6_2ZTGIf(31) => b6_2ZTGIf(31), b6_2ZTGIf(30) => 
        b6_2ZTGIf(30), b6_2ZTGIf(29) => b6_2ZTGIf(29), 
        b6_2ZTGIf(28) => b6_2ZTGIf(28), b6_2ZTGIf(27) => 
        b6_2ZTGIf(27), b6_2ZTGIf(26) => b6_2ZTGIf(26), 
        b6_2ZTGIf(25) => b6_2ZTGIf(25), b6_2ZTGIf(24) => 
        b6_2ZTGIf(24), b6_2ZTGIf(23) => b6_2ZTGIf(23), 
        b6_2ZTGIf(22) => b6_2ZTGIf(22), b6_2ZTGIf(21) => 
        b6_2ZTGIf(21), b6_2ZTGIf(20) => b6_2ZTGIf(20), 
        b6_2ZTGIf(19) => b6_2ZTGIf(19), b6_2ZTGIf(18) => 
        b6_2ZTGIf(18), b6_2ZTGIf(17) => b6_2ZTGIf(17), 
        b6_2ZTGIf(16) => b6_2ZTGIf(16), b13_CZS0wfY_d_FH9_0 => 
        \b13_CZS0wfY_d_FH9[1]\);
    
    b27_O2yyf_fG2_MiQA1E6_r_lnxob_S : b9_O2yyf_fG2_x_8_0
      port map(b6_2ZTGIf(111) => b6_2ZTGIf(111), b6_2ZTGIf(110)
         => b6_2ZTGIf(110), b6_2ZTGIf(109) => b6_2ZTGIf(109), 
        b6_2ZTGIf(108) => b6_2ZTGIf(108), b6_2ZTGIf(107) => 
        b6_2ZTGIf(107), b6_2ZTGIf(106) => b6_2ZTGIf(106), 
        b6_2ZTGIf(105) => b6_2ZTGIf(105), b6_2ZTGIf(104) => 
        b6_2ZTGIf(104), b6_2ZTGIf(103) => b6_2ZTGIf(103), 
        b6_2ZTGIf(102) => b6_2ZTGIf(102), b6_2ZTGIf(101) => 
        b6_2ZTGIf(101), b6_2ZTGIf(100) => b6_2ZTGIf(100), 
        b6_2ZTGIf(99) => b6_2ZTGIf(99), b6_2ZTGIf(98) => 
        b6_2ZTGIf(98), b6_2ZTGIf(97) => b6_2ZTGIf(97), 
        b6_2ZTGIf(96) => b6_2ZTGIf(96), b13_CZS0wfY_d_FH9_0 => 
        \b13_CZS0wfY_d_FH9[6]\);
    
    \b14_CZS0wfY_d_FH9m[10]\ : SLE
      port map(D => \b13_CZS0wfY_d_FH9[10]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b14_CZS0wfY_d_FH9m[10]_net_1\);
    
    \b14_CZS0wfY_d_FH9m[8]\ : SLE
      port map(D => \b13_CZS0wfY_d_FH9[8]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b14_CZS0wfY_d_FH9m[8]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_117_0 is

    port( b4_nUAi           : in    std_logic_vector(152 downto 150);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_117_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_117_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_61, b3_P_F_6_2_61, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(152), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(150), D => b4_nUAi(151), Y => b3_P_F_6_2_61);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(151), D => b4_nUAi(150), Y => b3_P_F_6_0_61);
    
    b3_P_F_6_0_RNI56SG2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_61, B => b4_nUAi(151), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_61, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(152), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(150), D => b4_nUAi(151), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_85_0 is

    port( b4_nUAi           : in    std_logic_vector(248 downto 246);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_85_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_85_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_93, b3_P_F_6_2_93, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(248), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(246), D => b4_nUAi(247), Y => b3_P_F_6_2_93);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(247), D => b4_nUAi(246), Y => b3_P_F_6_0_93);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(248), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(246), D => b4_nUAi(247), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNIIJQ52 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_93, B => b4_nUAi(247), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_93, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_46_0 is

    port( b4_nUAi           : in    std_logic_vector(365 downto 363);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_46_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_46_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_113, b3_P_F_6_2_113, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(365), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(363), D => b4_nUAi(364), Y => b3_P_F_6_2_113);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNIH3532 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_113, B => b4_nUAi(364), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_113, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(364), D => b4_nUAi(363), Y => b3_P_F_6_0_113);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(365), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(363), D => b4_nUAi(364), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_142_0 is

    port( b4_nUAi           : in    std_logic_vector(77 downto 75);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_142_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_142_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_140, b3_P_F_6_2_140, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(77), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(75), D => b4_nUAi(76), Y => b3_P_F_6_2_140);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(76), D => b4_nUAi(75), Y => b3_P_F_6_0_140);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(77), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(75), D => b4_nUAi(76), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNI49IC2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_140, B => b4_nUAi(76), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_140, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_102_0 is

    port( b4_nUAi           : in    std_logic_vector(197 downto 195);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_102_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_102_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_78, b3_P_F_6_2_78, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(197), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(195), D => b4_nUAi(196), Y => b3_P_F_6_2_78);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNIEDH52 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_78, B => b4_nUAi(196), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_78, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(196), D => b4_nUAi(195), Y => b3_P_F_6_0_78);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(197), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(195), D => b4_nUAi(196), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_133_0 is

    port( b4_nUAi           : in    std_logic_vector(104 downto 102);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_133_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_133_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_45, b3_P_F_6_2_45, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(104), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(102), D => b4_nUAi(103), Y => b3_P_F_6_2_45);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNIVO5D2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_45, B => b4_nUAi(103), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_45, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(103), D => b4_nUAi(102), Y => b3_P_F_6_0_45);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(104), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(102), D => b4_nUAi(103), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_3_0 is

    port( b4_nUAi           : in    std_logic_vector(494 downto 492);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_3_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_3_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_151, b3_P_F_6_2_151, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(494), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(492), D => b4_nUAi(493), Y => b3_P_F_6_2_151);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(493), D => b4_nUAi(492), Y => b3_P_F_6_0_151);
    
    b3_P_F_6_0_RNI5JAV2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_151, B => b4_nUAi(493), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_151, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(494), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(492), D => b4_nUAi(493), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_1_0 is

    port( b4_nUAi           : in    std_logic_vector(500 downto 498);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_1_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_1_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_138, b3_P_F_6_2_138, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(500), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(498), D => b4_nUAi(499), Y => b3_P_F_6_2_138);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(499), D => b4_nUAi(498), Y => b3_P_F_6_0_138);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(500), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(498), D => b4_nUAi(499), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNIDJIE2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_138, B => b4_nUAi(499), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_138, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_103_0 is

    port( b4_nUAi           : in    std_logic_vector(194 downto 192);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_103_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_103_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_79, b3_P_F_6_2_79, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(194), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(192), D => b4_nUAi(193), Y => b3_P_F_6_2_79);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(193), D => b4_nUAi(192), Y => b3_P_F_6_0_79);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(194), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(192), D => b4_nUAi(193), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNIQC0U2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_79, B => b4_nUAi(193), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_79, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_23_0 is

    port( b4_nUAi           : in    std_logic_vector(434 downto 432);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_23_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_23_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_149, b3_P_F_6_2_149, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(434), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(432), D => b4_nUAi(433), Y => b3_P_F_6_2_149);
    
    b3_P_F_6_0_RNIAFVM3 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_149, B => b4_nUAi(433), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_149, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(433), D => b4_nUAi(432), Y => b3_P_F_6_0_149);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(434), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(432), D => b4_nUAi(433), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_21_0 is

    port( b4_nUAi           : in    std_logic_vector(440 downto 438);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_21_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_21_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_36, b3_P_F_6_2_36, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(440), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(438), D => b4_nUAi(439), Y => b3_P_F_6_2_36);
    
    b3_P_F_6_0_RNIPTMA3 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_36, B => b4_nUAi(439), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_36, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(439), D => b4_nUAi(438), Y => b3_P_F_6_0_36);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(440), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(438), D => b4_nUAi(439), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_14_0 is

    port( b4_nUAi           : in    std_logic_vector(461 downto 459);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_14_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_14_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_29, b3_P_F_6_2_29, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(461), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(459), D => b4_nUAi(460), Y => b3_P_F_6_2_29);
    
    b3_P_F_6_0_RNIKCQ63 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_29, B => b4_nUAi(460), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_29, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(460), D => b4_nUAi(459), Y => b3_P_F_6_0_29);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(461), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(459), D => b4_nUAi(460), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_143_0 is

    port( b4_nUAi           : in    std_logic_vector(74 downto 72);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_143_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_143_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_141, b3_P_F_6_2_141, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNIGO1B2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_141, B => b4_nUAi(73), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_141, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(74), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(72), D => b4_nUAi(73), Y => b3_P_F_6_2_141);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(73), D => b4_nUAi(72), Y => b3_P_F_6_0_141);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(74), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(72), D => b4_nUAi(73), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_145_0 is

    port( b4_nUAi           : in    std_logic_vector(68 downto 66);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_145_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_145_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_162, b3_P_F_6_2_162, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(68), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(66), D => b4_nUAi(67), Y => b3_P_F_6_2_162);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(67), D => b4_nUAi(66), Y => b3_P_F_6_0_162);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(68), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(66), D => b4_nUAi(67), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNIC57B2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_162, B => b4_nUAi(67), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_162, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_105_0 is

    port( b4_nUAi           : in    std_logic_vector(188 downto 186);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_105_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_105_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_49, b3_P_F_6_2_49, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNID1743 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_49, B => b4_nUAi(187), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_49, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(188), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(186), D => b4_nUAi(187), Y => b3_P_F_6_2_49);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(187), D => b4_nUAi(186), Y => b3_P_F_6_0_49);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(188), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(186), D => b4_nUAi(187), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_126_0 is

    port( b4_nUAi           : in    std_logic_vector(125 downto 123);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_126_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_126_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_38, b3_P_F_6_2_38, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(125), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(123), D => b4_nUAi(124), Y => b3_P_F_6_2_38);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNI15RI2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_38, B => b4_nUAi(124), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_38, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(124), D => b4_nUAi(123), Y => b3_P_F_6_0_38);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(125), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(123), D => b4_nUAi(124), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_89_0 is

    port( b4_nUAi           : in    std_logic_vector(236 downto 234);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_89_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_89_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_65, b3_P_F_6_2_65, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(236), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(234), D => b4_nUAi(235), Y => b3_P_F_6_2_65);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(235), D => b4_nUAi(234), Y => b3_P_F_6_0_65);
    
    b3_P_F_6_0_RNIN9832 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_65, B => b4_nUAi(235), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_65, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(236), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(234), D => b4_nUAi(235), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_149_0 is

    port( b4_nUAi           : in    std_logic_vector(56 downto 54);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_149_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_149_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_147, b3_P_F_6_2_147, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(56), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(54), D => b4_nUAi(55), Y => b3_P_F_6_2_147);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(55), D => b4_nUAi(54), Y => b3_P_F_6_0_147);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(56), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(54), D => b4_nUAi(55), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNIERPM2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_147, B => b4_nUAi(55), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_147, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_80_0 is

    port( b4_nUAi           : in    std_logic_vector(263 downto 261);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_80_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_80_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_88, b3_P_F_6_2_88, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(263), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(261), D => b4_nUAi(262), Y => b3_P_F_6_2_88);
    
    b3_P_F_6_0_RNIM53J2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_88, B => b4_nUAi(262), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_88, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(262), D => b4_nUAi(261), Y => b3_P_F_6_0_88);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(263), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(261), D => b4_nUAi(262), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_127_0 is

    port( b4_nUAi           : in    std_logic_vector(122 downto 120);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_127_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_127_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_39, b3_P_F_6_2_39, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(122), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(120), D => b4_nUAi(121), Y => b3_P_F_6_2_39);
    
    b3_P_F_6_0_RNIARPM2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_39, B => b4_nUAi(121), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_39, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(121), D => b4_nUAi(120), Y => b3_P_F_6_0_39);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(122), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(120), D => b4_nUAi(121), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_131_0 is

    port( b4_nUAi           : in    std_logic_vector(110 downto 108);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_131_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_131_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_43, b3_P_F_6_2_43, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(110), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(108), D => b4_nUAi(109), Y => b3_P_F_6_2_43);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(109), D => b4_nUAi(108), Y => b3_P_F_6_0_43);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(110), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(108), D => b4_nUAi(109), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNINBJ13 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_43, B => b4_nUAi(109), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_43, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_109_0 is

    port( b4_nUAi           : in    std_logic_vector(176 downto 174);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_109_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_109_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_3, b3_P_F_6_2_3, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(176), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(174), D => b4_nUAi(175), Y => b3_P_F_6_2_3);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(175), D => b4_nUAi(174), Y => b3_P_F_6_0_3);
    
    b3_P_F_6_0_RNI38992 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_3, B => b4_nUAi(175), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_3, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(176), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(174), D => b4_nUAi(175), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_44_0 is

    port( b4_nUAi           : in    std_logic_vector(371 downto 369);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_44_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_44_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_111, b3_P_F_6_2_111, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(371), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(369), D => b4_nUAi(370), Y => b3_P_F_6_2_111);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNICR202 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_111, B => b4_nUAi(370), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_111, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(370), D => b4_nUAi(369), Y => b3_P_F_6_0_111);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(371), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(369), D => b4_nUAi(370), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_88_0 is

    port( b4_nUAi           : in    std_logic_vector(239 downto 237);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_88_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_88_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_64, b3_P_F_6_2_64, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(239), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(237), D => b4_nUAi(238), Y => b3_P_F_6_2_64);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(238), D => b4_nUAi(237), Y => b3_P_F_6_0_64);
    
    b3_P_F_6_0_RNIO8702 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_64, B => b4_nUAi(238), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_64, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(239), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(237), D => b4_nUAi(238), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_148_0 is

    port( b4_nUAi           : in    std_logic_vector(59 downto 57);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_148_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_148_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_165, b3_P_F_6_2_165, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(59), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(57), D => b4_nUAi(58), Y => b3_P_F_6_2_165);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(58), D => b4_nUAi(57), Y => b3_P_F_6_0_165);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(59), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(57), D => b4_nUAi(58), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNIMAEK2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_165, B => b4_nUAi(58), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_165, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_33_0 is

    port( b4_nUAi           : in    std_logic_vector(404 downto 402);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_33_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_33_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_130, b3_P_F_6_2_130, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNIU6JR2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_130, B => b4_nUAi(403), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_130, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(404), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(402), D => b4_nUAi(403), Y => b3_P_F_6_2_130);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(403), D => b4_nUAi(402), Y => b3_P_F_6_0_130);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(404), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(402), D => b4_nUAi(403), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_108_0 is

    port( b4_nUAi           : in    std_logic_vector(179 downto 177);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_108_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_108_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_2, b3_P_F_6_2_2, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(179), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(177), D => b4_nUAi(178), Y => b3_P_F_6_2_2);
    
    b3_P_F_6_0_RNI47862 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_2, B => b4_nUAi(178), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_2, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(178), D => b4_nUAi(177), Y => b3_P_F_6_0_2);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(179), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(177), D => b4_nUAi(178), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_163_0 is

    port( b4_nUAi           : in    std_logic_vector(14 downto 12);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_163_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_163_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_58, b3_P_F_6_2_58, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(14), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(12), D => b4_nUAi(13), Y => b3_P_F_6_2_58);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(13), D => b4_nUAi(12), Y => b3_P_F_6_0_58);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(14), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(12), D => b4_nUAi(13), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNIM2MS2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_58, B => b4_nUAi(13), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_58, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_31_0 is

    port( b4_nUAi           : in    std_logic_vector(410 downto 408);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_31_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_31_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_128, b3_P_F_6_2_128, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNI81HC3 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_128, B => b4_nUAi(409), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_128, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(410), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(408), D => b4_nUAi(409), Y => b3_P_F_6_2_128);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(409), D => b4_nUAi(408), Y => b3_P_F_6_0_128);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(410), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(408), D => b4_nUAi(409), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_140_0 is

    port( b4_nUAi           : in    std_logic_vector(83 downto 81);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_140_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_140_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_103, b3_P_F_6_2_103, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(83), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(81), D => b4_nUAi(82), Y => b3_P_F_6_2_103);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(82), D => b4_nUAi(81), Y => b3_P_F_6_0_103);
    
    b3_P_F_6_0_RNI09RC2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_103, B => b4_nUAi(82), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_103, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(83), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(81), D => b4_nUAi(82), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_100_0 is

    port( b4_nUAi           : in    std_logic_vector(203 downto 201);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_100_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_100_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_76, b3_P_F_6_2_76, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(203), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(201), D => b4_nUAi(202), Y => b3_P_F_6_2_76);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNI15R52 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_76, B => b4_nUAi(202), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_76, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(202), D => b4_nUAi(201), Y => b3_P_F_6_0_76);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(203), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(201), D => b4_nUAi(202), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_53_0 is

    port( b4_nUAi           : in    std_logic_vector(344 downto 342);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_53_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_53_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_120, b3_P_F_6_2_120, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(344), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(342), D => b4_nUAi(343), Y => b3_P_F_6_2_120);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(343), D => b4_nUAi(342), Y => b3_P_F_6_0_120);
    
    b3_P_F_6_0_RNIUT7L1 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_120, B => b4_nUAi(343), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_120, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(344), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(342), D => b4_nUAi(343), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_71_0 is

    port( b4_nUAi           : in    std_logic_vector(290 downto 288);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_71_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_71_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_106, b3_P_F_6_2_106, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(290), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(288), D => b4_nUAi(289), Y => b3_P_F_6_2_106);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNI43M22 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_106, B => b4_nUAi(289), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_106, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(289), D => b4_nUAi(288), Y => b3_P_F_6_0_106);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(290), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(288), D => b4_nUAi(289), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_51_0 is

    port( b4_nUAi           : in    std_logic_vector(350 downto 348);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_51_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_51_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_118, b3_P_F_6_2_118, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(350), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(348), D => b4_nUAi(349), Y => b3_P_F_6_2_118);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNIM2SG1 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_118, B => b4_nUAi(349), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_118, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(349), D => b4_nUAi(348), Y => b3_P_F_6_0_118);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(350), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(348), D => b4_nUAi(349), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_63_0 is

    port( b4_nUAi           : in    std_logic_vector(314 downto 312);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_63_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_63_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_10, b3_P_F_6_2_10, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(314), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(312), D => b4_nUAi(313), Y => b3_P_F_6_2_10);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(313), D => b4_nUAi(312), Y => b3_P_F_6_0_10);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(314), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(312), D => b4_nUAi(313), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNIB4JP1 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_10, B => b4_nUAi(313), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_10, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_134_0 is

    port( b4_nUAi           : in    std_logic_vector(101 downto 99);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_134_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_134_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_46, b3_P_F_6_2_46, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNIAAOU1 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_46, B => b4_nUAi(100), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_46, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(101), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(99), D => b4_nUAi(100), Y => b3_P_F_6_2_46);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(100), D => b4_nUAi(99), Y => b3_P_F_6_0_46);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(101), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(99), D => b4_nUAi(100), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_61_0 is

    port( b4_nUAi           : in    std_logic_vector(320 downto 318);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_61_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_61_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_101, b3_P_F_6_2_101, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(320), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(318), D => b4_nUAi(319), Y => b3_P_F_6_2_101);
    
    b3_P_F_6_0_RNIQ08L1 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_101, B => b4_nUAi(319), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_101, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(319), D => b4_nUAi(318), Y => b3_P_F_6_0_101);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(320), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(318), D => b4_nUAi(319), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_119_0 is

    port( b4_nUAi           : in    std_logic_vector(146 downto 144);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_119_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_119_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_63, b3_P_F_6_2_63, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(146), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(144), D => b4_nUAi(145), Y => b3_P_F_6_2_63);
    
    b3_P_F_6_0_RNIADQ92 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_63, B => b4_nUAi(145), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_63, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(145), D => b4_nUAi(144), Y => b3_P_F_6_0_63);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(146), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(144), D => b4_nUAi(145), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_92_0 is

    port( b4_nUAi           : in    std_logic_vector(227 downto 225);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_92_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_92_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_68, b3_P_F_6_2_68, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(227), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(225), D => b4_nUAi(226), Y => b3_P_F_6_2_68);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(226), D => b4_nUAi(225), Y => b3_P_F_6_0_68);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(227), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(225), D => b4_nUAi(226), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNIEFTI2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_68, B => b4_nUAi(226), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_68, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_152_0 is

    port( b4_nUAi           : in    std_logic_vector(47 downto 45);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_152_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_152_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_156, b3_P_F_6_2_156, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(47), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(45), D => b4_nUAi(46), Y => b3_P_F_6_2_156);
    
    b3_P_F_6_0_RNI51F63 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_156, B => b4_nUAi(46), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_156, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(46), D => b4_nUAi(45), Y => b3_P_F_6_0_156);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(47), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(45), D => b4_nUAi(46), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_160_0 is

    port( b4_nUAi           : in    std_logic_vector(23 downto 21);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_160_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_160_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_55, b3_P_F_6_2_55, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(23), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(21), D => b4_nUAi(22), Y => b3_P_F_6_2_55);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(22), D => b4_nUAi(21), Y => b3_P_F_6_0_55);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(23), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(21), D => b4_nUAi(22), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNICKPT2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_55, B => b4_nUAi(22), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_55, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_112_0 is

    port( b4_nUAi           : in    std_logic_vector(167 downto 165);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_112_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_112_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_6, b3_P_F_6_2_6, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(167), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(165), D => b4_nUAi(166), Y => b3_P_F_6_2_6);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(166), D => b4_nUAi(165), Y => b3_P_F_6_0_6);
    
    b3_P_F_6_0_RNIH5VO2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_6, B => b4_nUAi(166), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_6, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(167), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(165), D => b4_nUAi(166), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_118_0 is

    port( b4_nUAi           : in    std_logic_vector(149 downto 147);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_118_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_118_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_62, b3_P_F_6_2_62, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNIK4762 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_62, B => b4_nUAi(148), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_62, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(149), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(147), D => b4_nUAi(148), Y => b3_P_F_6_2_62);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(148), D => b4_nUAi(147), Y => b3_P_F_6_0_62);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(149), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(147), D => b4_nUAi(148), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_136_0 is

    port( b4_nUAi           : in    std_logic_vector(95 downto 93);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_136_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_136_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_163, b3_P_F_6_2_163, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNICJ0B2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_163, B => b4_nUAi(94), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_163, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(95), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(93), D => b4_nUAi(94), Y => b3_P_F_6_2_163);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(94), D => b4_nUAi(93), Y => b3_P_F_6_0_163);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(95), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(93), D => b4_nUAi(94), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_95_0 is

    port( b4_nUAi           : in    std_logic_vector(218 downto 216);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_95_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_95_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_71, b3_P_F_6_2_71, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(218), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(216), D => b4_nUAi(217), Y => b3_P_F_6_2_71);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(217), D => b4_nUAi(216), Y => b3_P_F_6_0_71);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(218), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(216), D => b4_nUAi(217), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNID3JH2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_71, B => b4_nUAi(217), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_71, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_155_0 is

    port( b4_nUAi           : in    std_logic_vector(38 downto 36);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_155_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_155_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_159, b3_P_F_6_2_159, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(38), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(36), D => b4_nUAi(37), Y => b3_P_F_6_2_159);
    
    b3_P_F_6_0_RNI4L453 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_159, B => b4_nUAi(37), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_159, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(37), D => b4_nUAi(36), Y => b3_P_F_6_0_159);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(38), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(36), D => b4_nUAi(37), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_137_0 is

    port( b4_nUAi           : in    std_logic_vector(92 downto 90);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_137_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_137_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_160, b3_P_F_6_2_160, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNILBLT2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_160, B => b4_nUAi(91), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_160, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(92), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(90), D => b4_nUAi(91), Y => b3_P_F_6_2_160);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(91), D => b4_nUAi(90), Y => b3_P_F_6_0_160);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(92), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(90), D => b4_nUAi(91), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_5_0 is

    port( b4_nUAi           : in    std_logic_vector(488 downto 486);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_5_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_5_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_153, b3_P_F_6_2_153, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(488), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(486), D => b4_nUAi(487), Y => b3_P_F_6_2_153);
    
    b3_P_F_6_0_RNI84LS3 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_153, B => b4_nUAi(487), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_153, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(487), D => b4_nUAi(486), Y => b3_P_F_6_0_153);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(488), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(486), D => b4_nUAi(487), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_115_0 is

    port( b4_nUAi           : in    std_logic_vector(158 downto 156);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_115_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_115_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_9, b3_P_F_6_2_9, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(158), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(156), D => b4_nUAi(157), Y => b3_P_F_6_2_9);
    
    b3_P_F_6_0_RNI0I9O2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_9, B => b4_nUAi(157), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_9, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(157), D => b4_nUAi(156), Y => b3_P_F_6_0_9);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(158), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(156), D => b4_nUAi(157), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_25_0 is

    port( b4_nUAi           : in    std_logic_vector(428 downto 426);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_25_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_25_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_124, b3_P_F_6_2_124, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(428), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(426), D => b4_nUAi(427), Y => b3_P_F_6_2_124);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(427), D => b4_nUAi(426), Y => b3_P_F_6_0_124);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(428), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(426), D => b4_nUAi(427), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNI6TRL3 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_124, B => b4_nUAi(427), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_124, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_74_0 is

    port( b4_nUAi           : in    std_logic_vector(281 downto 279);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_74_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_74_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_82, b3_P_F_6_2_82, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(281), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(279), D => b4_nUAi(280), Y => b3_P_F_6_2_82);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(280), D => b4_nUAi(279), Y => b3_P_F_6_0_82);
    
    b3_P_F_6_0_RNIK9V82 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_82, B => b4_nUAi(280), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_82, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(281), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(279), D => b4_nUAi(280), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_161_0 is

    port( b4_nUAi           : in    std_logic_vector(20 downto 18);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_161_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_161_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_56, b3_P_F_6_2_56, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNI7IGO2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_56, B => b4_nUAi(19), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_56, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(20), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(18), D => b4_nUAi(19), Y => b3_P_F_6_2_56);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(19), D => b4_nUAi(18), Y => b3_P_F_6_0_56);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(20), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(18), D => b4_nUAi(19), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_2_0 is

    port( b4_nUAi           : in    std_logic_vector(497 downto 495);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_2_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_2_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_139, b3_P_F_6_2_139, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(497), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(495), D => b4_nUAi(496), Y => b3_P_F_6_2_139);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(496), D => b4_nUAi(495), Y => b3_P_F_6_0_139);
    
    b3_P_F_6_0_RNI9GM82 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_139, B => b4_nUAi(496), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_139, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(497), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(495), D => b4_nUAi(496), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_22_0 is

    port( b4_nUAi           : in    std_logic_vector(437 downto 435);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_22_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_22_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_37, b3_P_F_6_2_37, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(437), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(435), D => b4_nUAi(436), Y => b3_P_F_6_2_37);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNIUOF73 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_37, B => b4_nUAi(436), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_37, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(436), D => b4_nUAi(435), Y => b3_P_F_6_0_37);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(437), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(435), D => b4_nUAi(436), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_122_0 is

    port( b4_nUAi           : in    std_logic_vector(137 downto 135);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_122_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_122_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_34, b3_P_F_6_2_34, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(137), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(135), D => b4_nUAi(136), Y => b3_P_F_6_2_34);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNIOO8A2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_34, B => b4_nUAi(136), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_34, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(136), D => b4_nUAi(135), Y => b3_P_F_6_0_34);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(137), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(135), D => b4_nUAi(136), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_18_0 is

    port( b4_nUAi           : in    std_logic_vector(449 downto 447);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_18_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_18_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_144, b3_P_F_6_2_144, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(449), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(447), D => b4_nUAi(448), Y => b3_P_F_6_2_144);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(448), D => b4_nUAi(447), Y => b3_P_F_6_0_144);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(449), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(447), D => b4_nUAi(448), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNIHSE33 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_144, B => b4_nUAi(448), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_144, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_0_0 is

    port( b4_nUAi           : in    std_logic_vector(502 downto 501);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic;
          b12_PSyi_XlK_qHv  : in    std_logic
        );

end b8_1LbcQDr1_x_0_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_0_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_150, b3_P_F_6_2_150, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b12_PSyi_XlK_qHv, Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(501), D => b4_nUAi(502), Y => b3_P_F_6_2_150);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNISE9L2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_150, B => b4_nUAi(502), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_150, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(502), D => b4_nUAi(501), Y => b3_P_F_6_0_150);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b12_PSyi_XlK_qHv, B => \b3_P_F_6_4_1_1\, C
         => b4_nUAi(501), D => b4_nUAi(502), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_76_0 is

    port( b4_nUAi           : in    std_logic_vector(275 downto 273);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_76_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_76_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_84, b3_P_F_6_2_84, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(275), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(273), D => b4_nUAi(274), Y => b3_P_F_6_2_84);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(274), D => b4_nUAi(273), Y => b3_P_F_6_0_84);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(275), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(273), D => b4_nUAi(274), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNI6QIK2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_84, B => b4_nUAi(274), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_84, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_162_0 is

    port( b4_nUAi           : in    std_logic_vector(17 downto 15);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_162_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_162_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_57, b3_P_F_6_2_57, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(17), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(15), D => b4_nUAi(16), Y => b3_P_F_6_2_57);
    
    b3_P_F_6_0_RNIAR2P2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_57, B => b4_nUAi(16), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_57, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(16), D => b4_nUAi(15), Y => b3_P_F_6_0_57);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(17), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(15), D => b4_nUAi(16), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_19_0 is

    port( b4_nUAi           : in    std_logic_vector(446 downto 444);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_19_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_19_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_145, b3_P_F_6_2_145, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(446), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(444), D => b4_nUAi(445), Y => b3_P_F_6_2_145);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(445), D => b4_nUAi(444), Y => b3_P_F_6_0_145);
    
    b3_P_F_6_0_RNI4Q0N3 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_145, B => b4_nUAi(445), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_145, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(446), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(444), D => b4_nUAi(445), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_77_0 is

    port( b4_nUAi           : in    std_logic_vector(272 downto 270);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_77_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_77_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_85, b3_P_F_6_2_85, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(272), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(270), D => b4_nUAi(271), Y => b3_P_F_6_2_85);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(271), D => b4_nUAi(270), Y => b3_P_F_6_0_85);
    
    b3_P_F_6_0_RNIMF1R1 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_85, B => b4_nUAi(271), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_85, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(272), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(270), D => b4_nUAi(271), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_7_0 is

    port( b4_nUAi           : in    std_logic_vector(482 downto 480);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_7_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_7_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_155, b3_P_F_6_2_155, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(482), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(480), D => b4_nUAi(481), Y => b3_P_F_6_2_155);
    
    b3_P_F_6_0_RNIB0UL3 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_155, B => b4_nUAi(481), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_155, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(481), D => b4_nUAi(480), Y => b3_P_F_6_0_155);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(482), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(480), D => b4_nUAi(481), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_35_0 is

    port( b4_nUAi           : in    std_logic_vector(398 downto 396);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_35_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_35_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_20, b3_P_F_6_2_20, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(398), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(396), D => b4_nUAi(397), Y => b3_P_F_6_2_20);
    
    b3_P_F_6_0_RNIO3V12 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_20, B => b4_nUAi(397), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_20, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(397), D => b4_nUAi(396), Y => b3_P_F_6_0_20);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(398), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(396), D => b4_nUAi(397), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_20_0 is

    port( b4_nUAi           : in    std_logic_vector(443 downto 441);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_20_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_20_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_146, b3_P_F_6_2_146, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(443), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(441), D => b4_nUAi(442), Y => b3_P_F_6_2_146);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNIJPPH3 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_146, B => b4_nUAi(442), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_146, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(442), D => b4_nUAi(441), Y => b3_P_F_6_0_146);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(443), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(441), D => b4_nUAi(442), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_90_0 is

    port( b4_nUAi           : in    std_logic_vector(233 downto 231);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_90_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_90_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_66, b3_P_F_6_2_66, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(233), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(231), D => b4_nUAi(232), Y => b3_P_F_6_2_66);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNIHLRU1 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_66, B => b4_nUAi(232), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_66, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(232), D => b4_nUAi(231), Y => b3_P_F_6_0_66);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(233), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(231), D => b4_nUAi(232), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_150_0 is

    port( b4_nUAi           : in    std_logic_vector(53 downto 51);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_150_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_150_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_148, b3_P_F_6_2_148, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(53), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(51), D => b4_nUAi(52), Y => b3_P_F_6_2_148);
    
    b3_P_F_6_0_RNI87DI2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_148, B => b4_nUAi(52), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_148, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(52), D => b4_nUAi(51), Y => b3_P_F_6_0_148);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(53), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(51), D => b4_nUAi(52), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_113_0 is

    port( b4_nUAi           : in    std_logic_vector(164 downto 162);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_113_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_113_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_7, b3_P_F_6_2_7, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNI61RS2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_7, B => b4_nUAi(163), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_7, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(164), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(162), D => b4_nUAi(163), Y => b3_P_F_6_2_7);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(163), D => b4_nUAi(162), Y => b3_P_F_6_0_7);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(164), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(162), D => b4_nUAi(163), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_165_0 is

    port( b4_nUAi           : in    std_logic_vector(8 downto 6);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_165_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_165_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_131, b3_P_F_6_2_131, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(8), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(6), D => b4_nUAi(7), Y => b3_P_F_6_2_131);
    
    b3_P_F_6_0_RNI6NB42 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_131, B => b4_nUAi(7), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_131, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(7), D => b4_nUAi(6), Y => b3_P_F_6_0_131);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(8), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(6), D => b4_nUAi(7), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_110_0 is

    port( b4_nUAi           : in    std_logic_vector(173 downto 171);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_110_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_110_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_4, b3_P_F_6_2_4, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(173), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(171), D => b4_nUAi(172), Y => b3_P_F_6_2_4);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(172), D => b4_nUAi(171), Y => b3_P_F_6_0_4);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(173), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(171), D => b4_nUAi(172), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNITJS43 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_4, B => b4_nUAi(172), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_4, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_27_0 is

    port( b4_nUAi           : in    std_logic_vector(422 downto 420);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_27_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_27_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_126, b3_P_F_6_2_126, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(422), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(420), D => b4_nUAi(421), Y => b3_P_F_6_2_126);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(421), D => b4_nUAi(420), Y => b3_P_F_6_0_126);
    
    b3_P_F_6_0_RNI9BBJ3 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_126, B => b4_nUAi(421), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_126, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(422), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(420), D => b4_nUAi(421), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_129_0 is

    port( b4_nUAi           : in    std_logic_vector(116 downto 114);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_129_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_129_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_41, b3_P_F_6_2_41, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(116), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(114), D => b4_nUAi(115), Y => b3_P_F_6_2_41);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(115), D => b4_nUAi(114), Y => b3_P_F_6_0_41);
    
    b3_P_F_6_0_RNI0N3V2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_41, B => b4_nUAi(115), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_41, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(116), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(114), D => b4_nUAi(115), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_81_0 is

    port( b4_nUAi           : in    std_logic_vector(260 downto 258);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_81_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_81_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_89, b3_P_F_6_2_89, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(260), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(258), D => b4_nUAi(259), Y => b3_P_F_6_2_89);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNIJEVP1 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_89, B => b4_nUAi(259), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_89, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(259), D => b4_nUAi(258), Y => b3_P_F_6_0_89);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(260), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(258), D => b4_nUAi(259), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_125_0 is

    port( b4_nUAi           : in    std_logic_vector(128 downto 126);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_125_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_125_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_0, b3_P_F_6_2_0, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(128), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(126), D => b4_nUAi(127), Y => b3_P_F_6_2_0);
    
    b3_P_F_6_0_RNI7DAP2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_0, B => b4_nUAi(127), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_0, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(127), D => b4_nUAi(126), Y => b3_P_F_6_0_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(128), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(126), D => b4_nUAi(127), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_6_0 is

    port( b4_nUAi           : in    std_logic_vector(485 downto 483);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_6_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_6_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_154, b3_P_F_6_2_154, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNI28933 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_154, B => b4_nUAi(484), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_154, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(485), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(483), D => b4_nUAi(484), Y => b3_P_F_6_2_154);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(484), D => b4_nUAi(483), Y => b3_P_F_6_0_154);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(485), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(483), D => b4_nUAi(484), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_32_0 is

    port( b4_nUAi           : in    std_logic_vector(407 downto 405);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_32_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_32_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_129, b3_P_F_6_2_129, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(407), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(405), D => b4_nUAi(406), Y => b3_P_F_6_2_129);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(406), D => b4_nUAi(405), Y => b3_P_F_6_0_129);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(407), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(405), D => b4_nUAi(406), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNIDJOP2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_129, B => b4_nUAi(406), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_129, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_128_0 is

    port( b4_nUAi           : in    std_logic_vector(119 downto 117);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_128_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_128_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_40, b3_P_F_6_2_40, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(119), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(117), D => b4_nUAi(118), Y => b3_P_F_6_2_40);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(118), D => b4_nUAi(117), Y => b3_P_F_6_0_40);
    
    b3_P_F_6_0_RNI1M2S2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_40, B => b4_nUAi(118), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_40, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(119), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(117), D => b4_nUAi(118), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_26_0 is

    port( b4_nUAi           : in    std_logic_vector(425 downto 423);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_26_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_26_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_125, b3_P_F_6_2_125, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(425), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(423), D => b4_nUAi(424), Y => b3_P_F_6_2_125);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNI0LCF3 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_125, B => b4_nUAi(424), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_125, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(424), D => b4_nUAi(423), Y => b3_P_F_6_0_125);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(425), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(423), D => b4_nUAi(424), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_28_0 is

    port( b4_nUAi           : in    std_logic_vector(419 downto 417);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_28_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_28_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_17, b3_P_F_6_2_17, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNI9GSJ3 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_17, B => b4_nUAi(418), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_17, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(419), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(417), D => b4_nUAi(418), Y => b3_P_F_6_2_17);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(418), D => b4_nUAi(417), Y => b3_P_F_6_0_17);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(419), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(417), D => b4_nUAi(418), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_55_0 is

    port( b4_nUAi           : in    std_logic_vector(338 downto 336);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_55_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_55_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_122, b3_P_F_6_2_122, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNIQRK92 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_122, B => b4_nUAi(337), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_122, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(338), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(336), D => b4_nUAi(337), Y => b3_P_F_6_2_122);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(337), D => b4_nUAi(336), Y => b3_P_F_6_0_122);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(338), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(336), D => b4_nUAi(337), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_13_0 is

    port( b4_nUAi           : in    std_logic_vector(464 downto 462);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_13_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_13_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_28, b3_P_F_6_2_28, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(464), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(462), D => b4_nUAi(463), Y => b3_P_F_6_2_28);
    
    b3_P_F_6_0_RNI36NR3 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_28, B => b4_nUAi(463), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_28, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(463), D => b4_nUAi(462), Y => b3_P_F_6_0_28);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(464), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(462), D => b4_nUAi(463), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_65_0 is

    port( b4_nUAi           : in    std_logic_vector(308 downto 306);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_65_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_65_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_12, b3_P_F_6_2_12, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(308), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(306), D => b4_nUAi(307), Y => b3_P_F_6_2_12);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(307), D => b4_nUAi(306), Y => b3_P_F_6_0_12);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(308), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(306), D => b4_nUAi(307), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNI720E2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_12, B => b4_nUAi(307), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_12, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_29_0 is

    port( b4_nUAi           : in    std_logic_vector(416 downto 414);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_29_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_29_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_18, b3_P_F_6_2_18, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(416), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(414), D => b4_nUAi(415), Y => b3_P_F_6_2_18);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(415), D => b4_nUAi(414), Y => b3_P_F_6_0_18);
    
    b3_P_F_6_0_RNIS9403 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_18, B => b4_nUAi(415), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_18, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(416), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(414), D => b4_nUAi(415), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_11_0 is

    port( b4_nUAi           : in    std_logic_vector(470 downto 468);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_11_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_11_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_26, b3_P_F_6_2_26, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(470), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(468), D => b4_nUAi(469), Y => b3_P_F_6_2_26);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(469), D => b4_nUAi(468), Y => b3_P_F_6_0_26);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(470), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(468), D => b4_nUAi(469), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNIRABN3 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_26, B => b4_nUAi(469), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_26, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_30_0 is

    port( b4_nUAi           : in    std_logic_vector(413 downto 411);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_30_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_30_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_127, b3_P_F_6_2_127, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNIPKHI3 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_127, B => b4_nUAi(412), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_127, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(413), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(411), D => b4_nUAi(412), Y => b3_P_F_6_2_127);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(412), D => b4_nUAi(411), Y => b3_P_F_6_0_127);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(413), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(411), D => b4_nUAi(412), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_141_0 is

    port( b4_nUAi           : in    std_logic_vector(80 downto 78);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_141_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_141_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_104, b3_P_F_6_2_104, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(80), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(78), D => b4_nUAi(79), Y => b3_P_F_6_2_104);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(79), D => b4_nUAi(78), Y => b3_P_F_6_0_104);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(80), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(78), D => b4_nUAi(79), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNID0CV2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_104, B => b4_nUAi(79), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_104, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_167_0 is

    port( b4_nUAi           : in    std_logic_vector(2 downto 0);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_167_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_167_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_133, b3_P_F_6_2_133, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(2), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(0), D => b4_nUAi(1), Y => b3_P_F_6_2_133);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(1), D => b4_nUAi(0), Y => b3_P_F_6_0_133);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(2), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(0), D => b4_nUAi(1), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNI8TQK2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_133, B => b4_nUAi(1), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_133, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_37_0 is

    port( b4_nUAi           : in    std_logic_vector(392 downto 390);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_37_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_37_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_22, b3_P_F_6_2_22, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNIRV7R1 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_22, B => b4_nUAi(391), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_22, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(392), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(390), D => b4_nUAi(391), Y => b3_P_F_6_2_22);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(391), D => b4_nUAi(390), Y => b3_P_F_6_0_22);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(392), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(390), D => b4_nUAi(391), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_101_0 is

    port( b4_nUAi           : in    std_logic_vector(200 downto 198);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_101_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_101_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_77, b3_P_F_6_2_77, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNIUDNC2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_77, B => b4_nUAi(199), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_77, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(200), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(198), D => b4_nUAi(199), Y => b3_P_F_6_2_77);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(199), D => b4_nUAi(198), Y => b3_P_F_6_0_77);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(200), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(198), D => b4_nUAi(199), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_52_0 is

    port( b4_nUAi           : in    std_logic_vector(347 downto 345);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_52_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_52_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_119, b3_P_F_6_2_119, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(347), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(345), D => b4_nUAi(346), Y => b3_P_F_6_2_119);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(346), D => b4_nUAi(345), Y => b3_P_F_6_0_119);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(347), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(345), D => b4_nUAi(346), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNIR7VA2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_119, B => b4_nUAi(346), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_119, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_62_0 is

    port( b4_nUAi           : in    std_logic_vector(317 downto 315);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_62_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_62_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_102, b3_P_F_6_2_102, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(317), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(315), D => b4_nUAi(316), Y => b3_P_F_6_2_102);
    
    b3_P_F_6_0_RNIV5BF2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_102, B => b4_nUAi(316), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_102, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(316), D => b4_nUAi(315), Y => b3_P_F_6_0_102);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(317), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(315), D => b4_nUAi(316), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_69_0 is

    port( b4_nUAi           : in    std_logic_vector(296 downto 294);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_69_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_69_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_16, b3_P_F_6_2_16, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNIDE603 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_16, B => b4_nUAi(295), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_16, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(296), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(294), D => b4_nUAi(295), Y => b3_P_F_6_2_16);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(295), D => b4_nUAi(294), Y => b3_P_F_6_0_16);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(296), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(294), D => b4_nUAi(295), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_84_0 is

    port( b4_nUAi           : in    std_logic_vector(251 downto 249);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_84_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_84_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_92, b3_P_F_6_2_92, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNISU402 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_92, B => b4_nUAi(250), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_92, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(251), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(249), D => b4_nUAi(250), Y => b3_P_F_6_2_92);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(250), D => b4_nUAi(249), Y => b3_P_F_6_0_92);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(251), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(249), D => b4_nUAi(250), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_43_0 is

    port( b4_nUAi           : in    std_logic_vector(374 downto 372);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_43_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_43_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_110, b3_P_F_6_2_110, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(374), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(372), D => b4_nUAi(373), Y => b3_P_F_6_2_110);
    
    b3_P_F_6_0_RNI4A382 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_110, B => b4_nUAi(373), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_110, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(373), D => b4_nUAi(372), Y => b3_P_F_6_0_110);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(374), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(372), D => b4_nUAi(373), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_120_0 is

    port( b4_nUAi           : in    std_logic_vector(143 downto 141);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_120_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_120_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_32, b3_P_F_6_2_32, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNI4HJK2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_32, B => b4_nUAi(142), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_32, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(143), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(141), D => b4_nUAi(142), Y => b3_P_F_6_2_32);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(142), D => b4_nUAi(141), Y => b3_P_F_6_0_32);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(143), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(141), D => b4_nUAi(142), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_48_0 is

    port( b4_nUAi           : in    std_logic_vector(359 downto 357);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_48_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_48_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_115, b3_P_F_6_2_115, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(359), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(357), D => b4_nUAi(358), Y => b3_P_F_6_2_115);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(358), D => b4_nUAi(357), Y => b3_P_F_6_0_115);
    
    b3_P_F_6_0_RNI5K452 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_115, B => b4_nUAi(358), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_115, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(359), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(357), D => b4_nUAi(358), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_41_0 is

    port( b4_nUAi           : in    std_logic_vector(380 downto 378);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_41_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_41_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_108, b3_P_F_6_2_108, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(380), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(378), D => b4_nUAi(379), Y => b3_P_F_6_2_108);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(379), D => b4_nUAi(378), Y => b3_P_F_6_0_108);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(380), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(378), D => b4_nUAi(379), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNIJ6O32 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_108, B => b4_nUAi(379), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_108, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_36_0 is

    port( b4_nUAi           : in    std_logic_vector(395 downto 393);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_36_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_36_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_21, b3_P_F_6_2_21, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(395), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(393), D => b4_nUAi(394), Y => b3_P_F_6_2_21);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(394), D => b4_nUAi(393), Y => b3_P_F_6_0_21);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(395), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(393), D => b4_nUAi(394), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNII7J82 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_21, B => b4_nUAi(394), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_21, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_58_0 is

    port( b4_nUAi           : in    std_logic_vector(329 downto 327);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_58_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_58_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_98, b3_P_F_6_2_98, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(329), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(327), D => b4_nUAi(328), Y => b3_P_F_6_2_98);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(328), D => b4_nUAi(327), Y => b3_P_F_6_0_98);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(329), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(327), D => b4_nUAi(328), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNII7KS1 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_98, B => b4_nUAi(328), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_98, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_4_0 is

    port( b4_nUAi           : in    std_logic_vector(491 downto 489);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_4_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_4_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_152, b3_P_F_6_2_152, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(491), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(489), D => b4_nUAi(490), Y => b3_P_F_6_2_152);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNITV603 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_152, B => b4_nUAi(490), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_152, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(490), D => b4_nUAi(489), Y => b3_P_F_6_0_152);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(491), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(489), D => b4_nUAi(490), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_49_0 is

    port( b4_nUAi           : in    std_logic_vector(356 downto 354);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_49_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_49_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_116, b3_P_F_6_2_116, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(356), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(354), D => b4_nUAi(355), Y => b3_P_F_6_2_116);
    
    b3_P_F_6_0_RNIODCH2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_116, B => b4_nUAi(355), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_116, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(355), D => b4_nUAi(354), Y => b3_P_F_6_0_116);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(356), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(354), D => b4_nUAi(355), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_68_0 is

    port( b4_nUAi           : in    std_logic_vector(299 downto 297);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_68_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_68_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_15, b3_P_F_6_2_15, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNIED5T2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_15, B => b4_nUAi(298), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_15, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(299), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(297), D => b4_nUAi(298), Y => b3_P_F_6_2_15);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(298), D => b4_nUAi(297), Y => b3_P_F_6_0_15);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(299), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(297), D => b4_nUAi(298), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_132_0 is

    port( b4_nUAi           : in    std_logic_vector(107 downto 105);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_132_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_132_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_44, b3_P_F_6_2_44, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(107), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(105), D => b4_nUAi(106), Y => b3_P_F_6_2_44);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(106), D => b4_nUAi(105), Y => b3_P_F_6_0_44);
    
    b3_P_F_6_0_RNIEKPE2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_44, B => b4_nUAi(106), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_44, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(107), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(105), D => b4_nUAi(106), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_59_0 is

    port( b4_nUAi           : in    std_logic_vector(326 downto 324);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_59_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_59_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_99, b3_P_F_6_2_99, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(326), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(324), D => b4_nUAi(325), Y => b3_P_F_6_2_99);
    
    b3_P_F_6_0_RNIE9R82 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_99, B => b4_nUAi(325), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_99, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(325), D => b4_nUAi(324), Y => b3_P_F_6_0_99);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(326), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(324), D => b4_nUAi(325), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_164_0 is

    port( b4_nUAi           : in    std_logic_vector(11 downto 9);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_164_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_164_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_59, b3_P_F_6_2_59, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(11), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(9), D => b4_nUAi(10), Y => b3_P_F_6_2_59);
    
    b3_P_F_6_0_RNIJQ2I2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_59, B => b4_nUAi(10), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_59, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(10), D => b4_nUAi(9), Y => b3_P_F_6_0_59);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(11), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(9), D => b4_nUAi(10), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_50_0 is

    port( b4_nUAi           : in    std_logic_vector(353 downto 351);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_50_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_50_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_117, b3_P_F_6_2_117, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(353), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(351), D => b4_nUAi(352), Y => b3_P_F_6_2_117);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNIU0P32 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_117, B => b4_nUAi(352), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_117, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(352), D => b4_nUAi(351), Y => b3_P_F_6_0_117);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(353), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(351), D => b4_nUAi(352), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_24_0 is

    port( b4_nUAi           : in    std_logic_vector(431 downto 429);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_24_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_24_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_123, b3_P_F_6_2_123, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNIRSOB3 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_123, B => b4_nUAi(430), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_123, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(431), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(429), D => b4_nUAi(430), Y => b3_P_F_6_2_123);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(430), D => b4_nUAi(429), Y => b3_P_F_6_0_123);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(431), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(429), D => b4_nUAi(430), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_60_0 is

    port( b4_nUAi           : in    std_logic_vector(323 downto 321);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_60_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_60_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_100, b3_P_F_6_2_100, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(323), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(321), D => b4_nUAi(322), Y => b3_P_F_6_2_100);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(322), D => b4_nUAi(321), Y => b3_P_F_6_0_100);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(323), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(321), D => b4_nUAi(322), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNIBK8R1 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_100, B => b4_nUAi(322), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_100, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_57_0 is

    port( b4_nUAi           : in    std_logic_vector(332 downto 330);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_57_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_57_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_97, b3_P_F_6_2_97, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(332), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(330), D => b4_nUAi(331), Y => b3_P_F_6_2_97);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(331), D => b4_nUAi(330), Y => b3_P_F_6_0_97);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(332), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(330), D => b4_nUAi(331), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNITNT22 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_97, B => b4_nUAi(331), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_97, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_67_0 is

    port( b4_nUAi           : in    std_logic_vector(302 downto 300);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_67_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_67_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_14, b3_P_F_6_2_14, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(302), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(300), D => b4_nUAi(301), Y => b3_P_F_6_2_14);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(301), D => b4_nUAi(300), Y => b3_P_F_6_0_14);
    
    b3_P_F_6_0_RNIDSRN2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_14, B => b4_nUAi(301), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_14, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(302), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(300), D => b4_nUAi(301), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_86_0 is

    port( b4_nUAi           : in    std_logic_vector(245 downto 243);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_86_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_86_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_94, b3_P_F_6_2_94, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(245), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(243), D => b4_nUAi(244), Y => b3_P_F_6_2_94);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNICNEC2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_94, B => b4_nUAi(244), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_94, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(244), D => b4_nUAi(243), Y => b3_P_F_6_0_94);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(245), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(243), D => b4_nUAi(244), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_87_0 is

    port( b4_nUAi           : in    std_logic_vector(242 downto 240);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_87_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_87_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_95, b3_P_F_6_2_95, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(242), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(240), D => b4_nUAi(241), Y => b3_P_F_6_2_95);
    
    b3_P_F_6_0_RNILF3V1 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_95, B => b4_nUAi(241), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_95, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(241), D => b4_nUAi(240), Y => b3_P_F_6_0_95);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(242), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(240), D => b4_nUAi(241), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_135_0 is

    port( b4_nUAi           : in    std_logic_vector(98 downto 96);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_135_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_135_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_47, b3_P_F_6_2_47, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(98), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(96), D => b4_nUAi(97), Y => b3_P_F_6_2_47);
    
    b3_P_F_6_0_RNI97D42 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_47, B => b4_nUAi(97), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_47, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(97), D => b4_nUAi(96), Y => b3_P_F_6_0_47);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(98), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(96), D => b4_nUAi(97), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_56_0 is

    port( b4_nUAi           : in    std_logic_vector(335 downto 333);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_56_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_56_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_96, b3_P_F_6_2_96, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(335), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(333), D => b4_nUAi(334), Y => b3_P_F_6_2_96);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(334), D => b4_nUAi(333), Y => b3_P_F_6_0_96);
    
    b3_P_F_6_0_RNIKV8G1 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_96, B => b4_nUAi(334), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_96, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(335), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(333), D => b4_nUAi(334), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_144_0 is

    port( b4_nUAi           : in    std_logic_vector(71 downto 69);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_144_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_144_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_142, b3_P_F_6_2_142, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(71), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(69), D => b4_nUAi(70), Y => b3_P_F_6_2_142);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNID8I53 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_142, B => b4_nUAi(70), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_142, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(70), D => b4_nUAi(69), Y => b3_P_F_6_0_142);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(71), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(69), D => b4_nUAi(70), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_104_0 is

    port( b4_nUAi           : in    std_logic_vector(191 downto 189);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_104_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_104_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_48, b3_P_F_6_2_48, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(191), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(189), D => b4_nUAi(190), Y => b3_P_F_6_2_48);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(190), D => b4_nUAi(189), Y => b3_P_F_6_0_48);
    
    b3_P_F_6_0_RNIE4IU2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_48, B => b4_nUAi(190), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_48, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(191), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(189), D => b4_nUAi(190), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_66_0 is

    port( b4_nUAi           : in    std_logic_vector(305 downto 303);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_66_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_66_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_13, b3_P_F_6_2_13, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(305), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(303), D => b4_nUAi(304), Y => b3_P_F_6_2_13);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(304), D => b4_nUAi(303), Y => b3_P_F_6_0_13);
    
    b3_P_F_6_0_RNIOKCL1 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_13, B => b4_nUAi(304), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_13, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(305), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(303), D => b4_nUAi(304), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_34_0 is

    port( b4_nUAi           : in    std_logic_vector(401 downto 399);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_34_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_34_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_19, b3_P_F_6_2_19, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(401), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(399), D => b4_nUAi(400), Y => b3_P_F_6_2_19);
    
    b3_P_F_6_0_RNIDVG52 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_19, B => b4_nUAi(400), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_19, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(400), D => b4_nUAi(399), Y => b3_P_F_6_0_19);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(401), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(399), D => b4_nUAi(400), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_72_0 is

    port( b4_nUAi           : in    std_logic_vector(287 downto 285);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_72_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_72_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_80, b3_P_F_6_2_80, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNIRBSF2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_80, B => b4_nUAi(286), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_80, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(287), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(285), D => b4_nUAi(286), Y => b3_P_F_6_2_80);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(286), D => b4_nUAi(285), Y => b3_P_F_6_0_80);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(287), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(285), D => b4_nUAi(286), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_159_0 is

    port( b4_nUAi           : in    std_logic_vector(26 downto 24);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_159_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_159_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_54, b3_P_F_6_2_54, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(26), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(24), D => b4_nUAi(25), Y => b3_P_F_6_2_54);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNIU8IL2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_54, B => b4_nUAi(25), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_54, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(25), D => b4_nUAi(24), Y => b3_P_F_6_0_54);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(26), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(24), D => b4_nUAi(25), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_146_0 is

    port( b4_nUAi           : in    std_logic_vector(65 downto 63);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_146_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_146_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_166, b3_P_F_6_2_166, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNI69RH2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_166, B => b4_nUAi(64), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_166, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(65), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(63), D => b4_nUAi(64), Y => b3_P_F_6_2_166);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(64), D => b4_nUAi(63), Y => b3_P_F_6_0_166);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(65), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(63), D => b4_nUAi(64), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_106_0 is

    port( b4_nUAi           : in    std_logic_vector(185 downto 183);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_106_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_106_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_50, b3_P_F_6_2_50, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(185), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(183), D => b4_nUAi(184), Y => b3_P_F_6_2_50);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNIGPCB2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_50, B => b4_nUAi(184), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_50, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(184), D => b4_nUAi(183), Y => b3_P_F_6_0_50);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(185), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(183), D => b4_nUAi(184), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_147_0 is

    port( b4_nUAi           : in    std_logic_vector(62 downto 60);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_147_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_147_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_164, b3_P_F_6_2_164, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(62), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(60), D => b4_nUAi(61), Y => b3_P_F_6_2_164);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNIV5N53 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_164, B => b4_nUAi(61), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_164, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(61), D => b4_nUAi(60), Y => b3_P_F_6_0_164);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(62), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(60), D => b4_nUAi(61), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_107_0 is

    port( b4_nUAi           : in    std_logic_vector(182 downto 180);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_107_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_107_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_1, b3_P_F_6_2_1, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(182), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(180), D => b4_nUAi(181), Y => b3_P_F_6_2_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(181), D => b4_nUAi(180), Y => b3_P_F_6_0_1);
    
    b3_P_F_6_0_RNIPH1U2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_1, B => b4_nUAi(181), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_1, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(182), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(180), D => b4_nUAi(181), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_75_0 is

    port( b4_nUAi           : in    std_logic_vector(278 downto 276);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_75_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_75_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_83, b3_P_F_6_2_83, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(278), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(276), D => b4_nUAi(277), Y => b3_P_F_6_2_83);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(277), D => b4_nUAi(276), Y => b3_P_F_6_0_83);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(278), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(276), D => b4_nUAi(277), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNIJ6KE2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_83, B => b4_nUAi(277), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_83, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_91_0 is

    port( b4_nUAi           : in    std_logic_vector(230 downto 228);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_91_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_91_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_67, b3_P_F_6_2_67, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(230), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(228), D => b4_nUAi(229), Y => b3_P_F_6_2_67);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(229), D => b4_nUAi(228), Y => b3_P_F_6_0_67);
    
    b3_P_F_6_0_RNIEUN52 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_67, B => b4_nUAi(229), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_67, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(230), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(228), D => b4_nUAi(229), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_151_0 is

    port( b4_nUAi           : in    std_logic_vector(50 downto 48);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_151_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_151_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_161, b3_P_F_6_2_161, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(50), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(48), D => b4_nUAi(49), Y => b3_P_F_6_2_161);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(49), D => b4_nUAi(48), Y => b3_P_F_6_0_161);
    
    b3_P_F_6_0_RNIEO8P2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_161, B => b4_nUAi(49), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_161, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(50), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(48), D => b4_nUAi(49), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_123_0 is

    port( b4_nUAi           : in    std_logic_vector(134 downto 132);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_123_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_123_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_35, b3_P_F_6_2_35, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(134), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(132), D => b4_nUAi(133), Y => b3_P_F_6_2_35);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNI4FOP2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_35, B => b4_nUAi(133), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_35, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(133), D => b4_nUAi(132), Y => b3_P_F_6_0_35);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(134), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(132), D => b4_nUAi(133), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_130_0 is

    port( b4_nUAi           : in    std_logic_vector(113 downto 111);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_130_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_130_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_42, b3_P_F_6_2_42, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNIQ2NQ2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_42, B => b4_nUAi(112), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_42, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(113), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(111), D => b4_nUAi(112), Y => b3_P_F_6_2_42);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(112), D => b4_nUAi(111), Y => b3_P_F_6_0_42);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(113), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(111), D => b4_nUAi(112), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_54_0 is

    port( b4_nUAi           : in    std_logic_vector(341 downto 339);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_54_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_54_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_121, b3_P_F_6_2_121, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNIFN6D2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_121, B => b4_nUAi(340), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_121, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(341), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(339), D => b4_nUAi(340), Y => b3_P_F_6_2_121);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(340), D => b4_nUAi(339), Y => b3_P_F_6_0_121);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(341), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(339), D => b4_nUAi(340), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_79_0 is

    port( b4_nUAi           : in    std_logic_vector(266 downto 264);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_79_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_79_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_87, b3_P_F_6_2_87, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(266), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(264), D => b4_nUAi(265), Y => b3_P_F_6_2_87);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(265), D => b4_nUAi(264), Y => b3_P_F_6_0_87);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(266), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(264), D => b4_nUAi(265), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNISPFN1 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_87, B => b4_nUAi(265), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_87, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_64_0 is

    port( b4_nUAi           : in    std_logic_vector(311 downto 309);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_64_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_64_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_11, b3_P_F_6_2_11, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(311), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(309), D => b4_nUAi(310), Y => b3_P_F_6_2_11);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(310), D => b4_nUAi(309), Y => b3_P_F_6_0_11);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(311), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(309), D => b4_nUAi(310), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNISTHH1 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_11, B => b4_nUAi(310), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_11, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_111_0 is

    port( b4_nUAi           : in    std_logic_vector(170 downto 168);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_111_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_111_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_5, b3_P_F_6_2_5, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(170), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(168), D => b4_nUAi(169), Y => b3_P_F_6_2_5);
    
    b3_P_F_6_0_RNIQSOB2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_5, B => b4_nUAi(169), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_5, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(169), D => b4_nUAi(168), Y => b3_P_F_6_0_5);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(170), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(168), D => b4_nUAi(169), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_83_0 is

    port( b4_nUAi           : in    std_logic_vector(254 downto 252);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_83_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_83_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_91, b3_P_F_6_2_91, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(254), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(252), D => b4_nUAi(253), Y => b3_P_F_6_2_91);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(253), D => b4_nUAi(252), Y => b3_P_F_6_0_91);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(254), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(252), D => b4_nUAi(253), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNIV4R12 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_91, B => b4_nUAi(253), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_91, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_15_0 is

    port( b4_nUAi           : in    std_logic_vector(458 downto 456);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_15_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_15_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_30, b3_P_F_6_2_30, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(458), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(456), D => b4_nUAi(457), Y => b3_P_F_6_2_30);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(457), D => b4_nUAi(456), Y => b3_P_F_6_0_30);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(458), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(456), D => b4_nUAi(457), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNIF51G3 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_30, B => b4_nUAi(457), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_30, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_78_0 is

    port( b4_nUAi           : in    std_logic_vector(269 downto 267);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_78_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_78_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_86, b3_P_F_6_2_86, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(269), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(267), D => b4_nUAi(268), Y => b3_P_F_6_2_86);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(268), D => b4_nUAi(267), Y => b3_P_F_6_0_86);
    
    b3_P_F_6_0_RNITOEK1 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_86, B => b4_nUAi(268), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_86, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(269), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(267), D => b4_nUAi(268), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_166_0 is

    port( b4_nUAi           : in    std_logic_vector(5 downto 3);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_166_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_166_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_132, b3_P_F_6_2_132, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNI3A4V2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_132, B => b4_nUAi(4), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_132, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(5), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(3), D => b4_nUAi(4), Y => b3_P_F_6_2_132);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(4), D => b4_nUAi(3), Y => b3_P_F_6_0_132);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(5), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(3), D => b4_nUAi(4), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_12_0 is

    port( b4_nUAi           : in    std_logic_vector(467 downto 465);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_12_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_12_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_27, b3_P_F_6_2_27, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(467), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(465), D => b4_nUAi(466), Y => b3_P_F_6_2_27);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(466), D => b4_nUAi(465), Y => b3_P_F_6_0_27);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(467), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(465), D => b4_nUAi(466), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNIN7FH3 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_27, B => b4_nUAi(466), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_27, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_73_0 is

    port( b4_nUAi           : in    std_logic_vector(284 downto 282);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_73_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_73_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_81, b3_P_F_6_2_81, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNI08JO2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_81, B => b4_nUAi(283), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_81, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(284), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(282), D => b4_nUAi(283), Y => b3_P_F_6_2_81);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(283), D => b4_nUAi(282), Y => b3_P_F_6_0_81);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(284), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(282), D => b4_nUAi(283), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_45_0 is

    port( b4_nUAi           : in    std_logic_vector(368 downto 366);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_45_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_45_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_112, b3_P_F_6_2_112, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(368), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(366), D => b4_nUAi(367), Y => b3_P_F_6_2_112);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNINVGS1 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_112, B => b4_nUAi(367), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_112, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(367), D => b4_nUAi(366), Y => b3_P_F_6_0_112);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(368), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(366), D => b4_nUAi(367), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_158_0 is

    port( b4_nUAi           : in    std_logic_vector(29 downto 27);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_158_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_158_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_53, b3_P_F_6_2_53, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(29), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(27), D => b4_nUAi(28), Y => b3_P_F_6_2_53);
    
    b3_P_F_6_0_RNIMVHI2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_53, B => b4_nUAi(28), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_53, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(28), D => b4_nUAi(27), Y => b3_P_F_6_0_53);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(29), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(27), D => b4_nUAi(28), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_8_0 is

    port( b4_nUAi           : in    std_logic_vector(479 downto 477);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_8_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_8_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_134, b3_P_F_6_2_134, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(479), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(477), D => b4_nUAi(478), Y => b3_P_F_6_2_134);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(478), D => b4_nUAi(477), Y => b3_P_F_6_0_134);
    
    b3_P_F_6_0_RNIA9OU2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_134, B => b4_nUAi(478), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_134, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(479), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(477), D => b4_nUAi(478), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_139_0 is

    port( b4_nUAi           : in    std_logic_vector(86 downto 84);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_139_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_139_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_137, b3_P_F_6_2_137, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(86), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(84), D => b4_nUAi(85), Y => b3_P_F_6_2_137);
    
    b3_P_F_6_0_RNI6T7H2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_137, B => b4_nUAi(85), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_137, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(85), D => b4_nUAi(84), Y => b3_P_F_6_0_137);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(86), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(84), D => b4_nUAi(85), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_9_0 is

    port( b4_nUAi           : in    std_logic_vector(476 downto 474);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_9_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_9_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_135, b3_P_F_6_2_135, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(476), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(474), D => b4_nUAi(475), Y => b3_P_F_6_2_135);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(475), D => b4_nUAi(474), Y => b3_P_F_6_0_135);
    
    b3_P_F_6_0_RNIT20B3 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_135, B => b4_nUAi(475), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_135, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(476), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(474), D => b4_nUAi(475), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_99_0 is

    port( b4_nUAi           : in    std_logic_vector(206 downto 204);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_99_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_99_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_75, b3_P_F_6_2_75, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(206), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(204), D => b4_nUAi(205), Y => b3_P_F_6_2_75);
    
    b3_P_F_6_0_RNIKFD62 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_75, B => b4_nUAi(205), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_75, Y => b6_2ZTGIf_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(205), D => b4_nUAi(204), Y => b3_P_F_6_0_75);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(206), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(204), D => b4_nUAi(205), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_70_0 is

    port( b4_nUAi           : in    std_logic_vector(293 downto 291);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_70_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_70_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_105, b3_P_F_6_2_105, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNI7QPR2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_105, B => b4_nUAi(292), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_105, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(293), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(291), D => b4_nUAi(292), Y => b3_P_F_6_2_105);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(292), D => b4_nUAi(291), Y => b3_P_F_6_0_105);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(293), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(291), D => b4_nUAi(292), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_94_0 is

    port( b4_nUAi           : in    std_logic_vector(221 downto 219);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_94_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_94_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_70, b3_P_F_6_2_70, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(221), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(219), D => b4_nUAi(220), Y => b3_P_F_6_2_70);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(220), D => b4_nUAi(219), Y => b3_P_F_6_0_70);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(221), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(219), D => b4_nUAi(220), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNIE6UB2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_70, B => b4_nUAi(220), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_70, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_154_0 is

    port( b4_nUAi           : in    std_logic_vector(41 downto 39);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_154_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_154_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_158, b3_P_F_6_2_158, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(41), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(39), D => b4_nUAi(40), Y => b3_P_F_6_2_158);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(40), D => b4_nUAi(39), Y => b3_P_F_6_0_158);
    
    b3_P_F_6_0_RNI5OFV2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_158, B => b4_nUAi(40), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_158, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(41), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(39), D => b4_nUAi(40), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_124_0 is

    port( b4_nUAi           : in    std_logic_vector(131 downto 129);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_124_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_124_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \b3_P_F_6_0\, \b3_P_F_6_2\, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(131), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(129), D => b4_nUAi(130), Y => \b3_P_F_6_2\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(130), D => b4_nUAi(129), Y => \b3_P_F_6_0\);
    
    b3_P_F_6_0_RNI1GIU2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => \b3_P_F_6_0\, B => b4_nUAi(130), C => 
        \b3_P_F_6_4_1\, D => \b3_P_F_6_2\, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(131), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(129), D => b4_nUAi(130), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_10_0 is

    port( b4_nUAi           : in    std_logic_vector(473 downto 471);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_10_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_10_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_25, b3_P_F_6_2_25, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(473), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(471), D => b4_nUAi(472), Y => b3_P_F_6_2_25);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNICUBT2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_25, B => b4_nUAi(472), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_25, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(472), D => b4_nUAi(471), Y => b3_P_F_6_0_25);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(473), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(471), D => b4_nUAi(472), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_42_0 is

    port( b4_nUAi           : in    std_logic_vector(377 downto 375);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_42_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_42_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_109, b3_P_F_6_2_109, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(377), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(375), D => b4_nUAi(376), Y => b3_P_F_6_2_109);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNIOBRT1 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_109, B => b4_nUAi(376), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_109, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(376), D => b4_nUAi(375), Y => b3_P_F_6_0_109);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(377), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(375), D => b4_nUAi(376), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_114_0 is

    port( b4_nUAi           : in    std_logic_vector(161 downto 159);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_114_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_114_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_8, b3_P_F_6_2_8, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNI1LKI2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_8, B => b4_nUAi(160), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_8, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(161), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(159), D => b4_nUAi(160), Y => b3_P_F_6_2_8);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(160), D => b4_nUAi(159), Y => b3_P_F_6_0_8);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(161), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(159), D => b4_nUAi(160), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_138_0 is

    port( b4_nUAi           : in    std_logic_vector(89 downto 87);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_138_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_138_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_136, b3_P_F_6_2_136, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    b3_P_F_6_0_RNIG46E2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_136, B => b4_nUAi(88), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_136, Y => b6_2ZTGIf_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(89), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(87), D => b4_nUAi(88), Y => b3_P_F_6_2_136);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(88), D => b4_nUAi(87), Y => b3_P_F_6_0_136);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(89), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(87), D => b4_nUAi(88), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_17_0 is

    port( b4_nUAi           : in    std_logic_vector(452 downto 450);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_17_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_17_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_143, b3_P_F_6_2_143, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(452), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(450), D => b4_nUAi(451), Y => b3_P_F_6_2_143);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(451), D => b4_nUAi(450), Y => b3_P_F_6_0_143);
    
    b3_P_F_6_0_RNIR9993 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_143, B => b4_nUAi(451), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_143, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(452), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(450), D => b4_nUAi(451), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_98_0 is

    port( b4_nUAi           : in    std_logic_vector(209 downto 207);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_98_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_98_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_74, b3_P_F_6_2_74, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(209), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(207), D => b4_nUAi(208), Y => b3_P_F_6_2_74);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNILEC32 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_74, B => b4_nUAi(208), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_74, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(208), D => b4_nUAi(207), Y => b3_P_F_6_0_74);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(209), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(207), D => b4_nUAi(208), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_121_0 is

    port( b4_nUAi           : in    std_logic_vector(140 downto 138);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_121_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_121_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_33, b3_P_F_6_2_33, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(140), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(138), D => b4_nUAi(139), Y => b3_P_F_6_2_33);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNI189N2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_33, B => b4_nUAi(139), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_33, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(139), D => b4_nUAi(138), Y => b3_P_F_6_0_33);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(140), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(138), D => b4_nUAi(139), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_38_0 is

    port( b4_nUAi           : in    std_logic_vector(389 downto 387);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_38_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_38_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_23, b3_P_F_6_2_23, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(389), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(387), D => b4_nUAi(388), Y => b3_P_F_6_2_23);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0_RNI255B2 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_23, B => b4_nUAi(388), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_23, Y => b6_2ZTGIf_0);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(388), D => b4_nUAi(387), Y => b3_P_F_6_0_23);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(389), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(387), D => b4_nUAi(388), Y => \b3_P_F_6_4_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_1LbcQDr1_x_82_0 is

    port( b4_nUAi           : in    std_logic_vector(257 downto 255);
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic;
          mdiclink_reg_0    : in    std_logic
        );

end b8_1LbcQDr1_x_82_0;

architecture DEF_ARCH of b8_1LbcQDr1_x_82_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal b3_P_F_6_0_90, b3_P_F_6_2_90, \b3_P_F_6_4_1_1\, 
        \b3_P_F_6_4_1\, GND_net_1, VCC_net_1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b3_P_F_6_4_1_1 : CFG3
      generic map(INIT => x"71")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(257), Y => \b3_P_F_6_4_1_1\);
    
    b3_P_F_6_2 : CFG4
      generic map(INIT => x"F045")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(255), D => b4_nUAi(256), Y => b3_P_F_6_2_90);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_P_F_6_0 : CFG4
      generic map(INIT => x"F20A")

      port map(A => mdiclink_reg_0, B => b11_OFWNT9L_8tZ_0, C => 
        b4_nUAi(256), D => b4_nUAi(255), Y => b3_P_F_6_0_90);
    
    b3_P_F_6_4_1 : CFG4
      generic map(INIT => x"9855")

      port map(A => b4_nUAi(257), B => \b3_P_F_6_4_1_1\, C => 
        b4_nUAi(255), D => b4_nUAi(256), Y => \b3_P_F_6_4_1\);
    
    b3_P_F_6_0_RNIAN572 : CFG4
      generic map(INIT => x"2F2C")

      port map(A => b3_P_F_6_0_90, B => b4_nUAi(256), C => 
        \b3_P_F_6_4_1\, D => b3_P_F_6_2_90, Y => b6_2ZTGIf_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b13_PSyil9s1fkJ_L_x is

    port( mdiclink_reg        : in    std_logic_vector(167 downto 0);
          b11_OFWNT9L_8tZ     : in    std_logic_vector(167 downto 0);
          b4_nUAi             : in    std_logic_vector(502 downto 0);
          b10_nYBzIXrKbK_0    : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          b12_PSyi_XlK_qHv    : in    std_logic
        );

end b13_PSyil9s1fkJ_L_x;

architecture DEF_ARCH of b13_PSyil9s1fkJ_L_x is 

  component b8_1LbcQDr1_x_39_0
    port( b4_nUAi           : in    std_logic_vector(386 downto 384) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_93_0
    port( b4_nUAi           : in    std_logic_vector(224 downto 222) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_16_0
    port( b4_nUAi           : in    std_logic_vector(455 downto 453) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_40_0
    port( b4_nUAi           : in    std_logic_vector(383 downto 381) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_153_0
    port( b4_nUAi           : in    std_logic_vector(44 downto 42) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_96_0
    port( b4_nUAi           : in    std_logic_vector(215 downto 213) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_156_0
    port( b4_nUAi           : in    std_logic_vector(35 downto 33) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_47_0
    port( b4_nUAi           : in    std_logic_vector(362 downto 360) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_97_0
    port( b4_nUAi           : in    std_logic_vector(212 downto 210) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_157_0
    port( b4_nUAi           : in    std_logic_vector(32 downto 30) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_116_0
    port( b4_nUAi           : in    std_logic_vector(155 downto 153) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b16_CRGcTCua_eH4_uaL_x_0
    port( b6_2ZTGIf           : in    std_logic_vector(167 downto 0) := (others => 'U');
          b10_nYBzIXrKbK_0    : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_117_0
    port( b4_nUAi           : in    std_logic_vector(152 downto 150) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_85_0
    port( b4_nUAi           : in    std_logic_vector(248 downto 246) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_46_0
    port( b4_nUAi           : in    std_logic_vector(365 downto 363) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_142_0
    port( b4_nUAi           : in    std_logic_vector(77 downto 75) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_102_0
    port( b4_nUAi           : in    std_logic_vector(197 downto 195) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_133_0
    port( b4_nUAi           : in    std_logic_vector(104 downto 102) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_3_0
    port( b4_nUAi           : in    std_logic_vector(494 downto 492) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_1_0
    port( b4_nUAi           : in    std_logic_vector(500 downto 498) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_103_0
    port( b4_nUAi           : in    std_logic_vector(194 downto 192) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_23_0
    port( b4_nUAi           : in    std_logic_vector(434 downto 432) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_21_0
    port( b4_nUAi           : in    std_logic_vector(440 downto 438) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_14_0
    port( b4_nUAi           : in    std_logic_vector(461 downto 459) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_143_0
    port( b4_nUAi           : in    std_logic_vector(74 downto 72) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_145_0
    port( b4_nUAi           : in    std_logic_vector(68 downto 66) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_105_0
    port( b4_nUAi           : in    std_logic_vector(188 downto 186) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_126_0
    port( b4_nUAi           : in    std_logic_vector(125 downto 123) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_89_0
    port( b4_nUAi           : in    std_logic_vector(236 downto 234) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_149_0
    port( b4_nUAi           : in    std_logic_vector(56 downto 54) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_80_0
    port( b4_nUAi           : in    std_logic_vector(263 downto 261) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_127_0
    port( b4_nUAi           : in    std_logic_vector(122 downto 120) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_131_0
    port( b4_nUAi           : in    std_logic_vector(110 downto 108) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_109_0
    port( b4_nUAi           : in    std_logic_vector(176 downto 174) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_44_0
    port( b4_nUAi           : in    std_logic_vector(371 downto 369) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component b8_1LbcQDr1_x_88_0
    port( b4_nUAi           : in    std_logic_vector(239 downto 237) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_148_0
    port( b4_nUAi           : in    std_logic_vector(59 downto 57) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_33_0
    port( b4_nUAi           : in    std_logic_vector(404 downto 402) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_108_0
    port( b4_nUAi           : in    std_logic_vector(179 downto 177) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_163_0
    port( b4_nUAi           : in    std_logic_vector(14 downto 12) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_31_0
    port( b4_nUAi           : in    std_logic_vector(410 downto 408) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_140_0
    port( b4_nUAi           : in    std_logic_vector(83 downto 81) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_100_0
    port( b4_nUAi           : in    std_logic_vector(203 downto 201) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_53_0
    port( b4_nUAi           : in    std_logic_vector(344 downto 342) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_71_0
    port( b4_nUAi           : in    std_logic_vector(290 downto 288) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_51_0
    port( b4_nUAi           : in    std_logic_vector(350 downto 348) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_63_0
    port( b4_nUAi           : in    std_logic_vector(314 downto 312) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_134_0
    port( b4_nUAi           : in    std_logic_vector(101 downto 99) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_61_0
    port( b4_nUAi           : in    std_logic_vector(320 downto 318) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_119_0
    port( b4_nUAi           : in    std_logic_vector(146 downto 144) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_92_0
    port( b4_nUAi           : in    std_logic_vector(227 downto 225) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_152_0
    port( b4_nUAi           : in    std_logic_vector(47 downto 45) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_160_0
    port( b4_nUAi           : in    std_logic_vector(23 downto 21) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_112_0
    port( b4_nUAi           : in    std_logic_vector(167 downto 165) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_118_0
    port( b4_nUAi           : in    std_logic_vector(149 downto 147) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component b8_1LbcQDr1_x_136_0
    port( b4_nUAi           : in    std_logic_vector(95 downto 93) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_95_0
    port( b4_nUAi           : in    std_logic_vector(218 downto 216) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_155_0
    port( b4_nUAi           : in    std_logic_vector(38 downto 36) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_137_0
    port( b4_nUAi           : in    std_logic_vector(92 downto 90) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_5_0
    port( b4_nUAi           : in    std_logic_vector(488 downto 486) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_115_0
    port( b4_nUAi           : in    std_logic_vector(158 downto 156) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_25_0
    port( b4_nUAi           : in    std_logic_vector(428 downto 426) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_74_0
    port( b4_nUAi           : in    std_logic_vector(281 downto 279) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_161_0
    port( b4_nUAi           : in    std_logic_vector(20 downto 18) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_2_0
    port( b4_nUAi           : in    std_logic_vector(497 downto 495) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_22_0
    port( b4_nUAi           : in    std_logic_vector(437 downto 435) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_122_0
    port( b4_nUAi           : in    std_logic_vector(137 downto 135) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_18_0
    port( b4_nUAi           : in    std_logic_vector(449 downto 447) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_0_0
    port( b4_nUAi           : in    std_logic_vector(502 downto 501) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U';
          b12_PSyi_XlK_qHv  : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_76_0
    port( b4_nUAi           : in    std_logic_vector(275 downto 273) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_162_0
    port( b4_nUAi           : in    std_logic_vector(17 downto 15) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_19_0
    port( b4_nUAi           : in    std_logic_vector(446 downto 444) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_77_0
    port( b4_nUAi           : in    std_logic_vector(272 downto 270) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_7_0
    port( b4_nUAi           : in    std_logic_vector(482 downto 480) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_35_0
    port( b4_nUAi           : in    std_logic_vector(398 downto 396) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_20_0
    port( b4_nUAi           : in    std_logic_vector(443 downto 441) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_90_0
    port( b4_nUAi           : in    std_logic_vector(233 downto 231) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_150_0
    port( b4_nUAi           : in    std_logic_vector(53 downto 51) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_113_0
    port( b4_nUAi           : in    std_logic_vector(164 downto 162) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_165_0
    port( b4_nUAi           : in    std_logic_vector(8 downto 6) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_110_0
    port( b4_nUAi           : in    std_logic_vector(173 downto 171) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_27_0
    port( b4_nUAi           : in    std_logic_vector(422 downto 420) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_129_0
    port( b4_nUAi           : in    std_logic_vector(116 downto 114) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_81_0
    port( b4_nUAi           : in    std_logic_vector(260 downto 258) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_125_0
    port( b4_nUAi           : in    std_logic_vector(128 downto 126) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_6_0
    port( b4_nUAi           : in    std_logic_vector(485 downto 483) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_32_0
    port( b4_nUAi           : in    std_logic_vector(407 downto 405) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_128_0
    port( b4_nUAi           : in    std_logic_vector(119 downto 117) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_26_0
    port( b4_nUAi           : in    std_logic_vector(425 downto 423) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_28_0
    port( b4_nUAi           : in    std_logic_vector(419 downto 417) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_55_0
    port( b4_nUAi           : in    std_logic_vector(338 downto 336) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_13_0
    port( b4_nUAi           : in    std_logic_vector(464 downto 462) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_65_0
    port( b4_nUAi           : in    std_logic_vector(308 downto 306) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_29_0
    port( b4_nUAi           : in    std_logic_vector(416 downto 414) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_11_0
    port( b4_nUAi           : in    std_logic_vector(470 downto 468) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_30_0
    port( b4_nUAi           : in    std_logic_vector(413 downto 411) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_141_0
    port( b4_nUAi           : in    std_logic_vector(80 downto 78) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_167_0
    port( b4_nUAi           : in    std_logic_vector(2 downto 0) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_37_0
    port( b4_nUAi           : in    std_logic_vector(392 downto 390) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_101_0
    port( b4_nUAi           : in    std_logic_vector(200 downto 198) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_52_0
    port( b4_nUAi           : in    std_logic_vector(347 downto 345) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_62_0
    port( b4_nUAi           : in    std_logic_vector(317 downto 315) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_69_0
    port( b4_nUAi           : in    std_logic_vector(296 downto 294) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_84_0
    port( b4_nUAi           : in    std_logic_vector(251 downto 249) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_43_0
    port( b4_nUAi           : in    std_logic_vector(374 downto 372) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_120_0
    port( b4_nUAi           : in    std_logic_vector(143 downto 141) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_48_0
    port( b4_nUAi           : in    std_logic_vector(359 downto 357) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_41_0
    port( b4_nUAi           : in    std_logic_vector(380 downto 378) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_36_0
    port( b4_nUAi           : in    std_logic_vector(395 downto 393) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_58_0
    port( b4_nUAi           : in    std_logic_vector(329 downto 327) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_4_0
    port( b4_nUAi           : in    std_logic_vector(491 downto 489) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_49_0
    port( b4_nUAi           : in    std_logic_vector(356 downto 354) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_68_0
    port( b4_nUAi           : in    std_logic_vector(299 downto 297) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_132_0
    port( b4_nUAi           : in    std_logic_vector(107 downto 105) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_59_0
    port( b4_nUAi           : in    std_logic_vector(326 downto 324) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_164_0
    port( b4_nUAi           : in    std_logic_vector(11 downto 9) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_50_0
    port( b4_nUAi           : in    std_logic_vector(353 downto 351) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_24_0
    port( b4_nUAi           : in    std_logic_vector(431 downto 429) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_60_0
    port( b4_nUAi           : in    std_logic_vector(323 downto 321) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_57_0
    port( b4_nUAi           : in    std_logic_vector(332 downto 330) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_67_0
    port( b4_nUAi           : in    std_logic_vector(302 downto 300) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_86_0
    port( b4_nUAi           : in    std_logic_vector(245 downto 243) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_87_0
    port( b4_nUAi           : in    std_logic_vector(242 downto 240) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_135_0
    port( b4_nUAi           : in    std_logic_vector(98 downto 96) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_56_0
    port( b4_nUAi           : in    std_logic_vector(335 downto 333) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_144_0
    port( b4_nUAi           : in    std_logic_vector(71 downto 69) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_104_0
    port( b4_nUAi           : in    std_logic_vector(191 downto 189) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_66_0
    port( b4_nUAi           : in    std_logic_vector(305 downto 303) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_34_0
    port( b4_nUAi           : in    std_logic_vector(401 downto 399) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_72_0
    port( b4_nUAi           : in    std_logic_vector(287 downto 285) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_159_0
    port( b4_nUAi           : in    std_logic_vector(26 downto 24) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_146_0
    port( b4_nUAi           : in    std_logic_vector(65 downto 63) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_106_0
    port( b4_nUAi           : in    std_logic_vector(185 downto 183) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_147_0
    port( b4_nUAi           : in    std_logic_vector(62 downto 60) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_107_0
    port( b4_nUAi           : in    std_logic_vector(182 downto 180) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_75_0
    port( b4_nUAi           : in    std_logic_vector(278 downto 276) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_91_0
    port( b4_nUAi           : in    std_logic_vector(230 downto 228) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_151_0
    port( b4_nUAi           : in    std_logic_vector(50 downto 48) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_123_0
    port( b4_nUAi           : in    std_logic_vector(134 downto 132) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_130_0
    port( b4_nUAi           : in    std_logic_vector(113 downto 111) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_54_0
    port( b4_nUAi           : in    std_logic_vector(341 downto 339) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_79_0
    port( b4_nUAi           : in    std_logic_vector(266 downto 264) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_64_0
    port( b4_nUAi           : in    std_logic_vector(311 downto 309) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_111_0
    port( b4_nUAi           : in    std_logic_vector(170 downto 168) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_83_0
    port( b4_nUAi           : in    std_logic_vector(254 downto 252) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_15_0
    port( b4_nUAi           : in    std_logic_vector(458 downto 456) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_78_0
    port( b4_nUAi           : in    std_logic_vector(269 downto 267) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_166_0
    port( b4_nUAi           : in    std_logic_vector(5 downto 3) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_12_0
    port( b4_nUAi           : in    std_logic_vector(467 downto 465) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_73_0
    port( b4_nUAi           : in    std_logic_vector(284 downto 282) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_45_0
    port( b4_nUAi           : in    std_logic_vector(368 downto 366) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_158_0
    port( b4_nUAi           : in    std_logic_vector(29 downto 27) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_8_0
    port( b4_nUAi           : in    std_logic_vector(479 downto 477) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_139_0
    port( b4_nUAi           : in    std_logic_vector(86 downto 84) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_9_0
    port( b4_nUAi           : in    std_logic_vector(476 downto 474) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_99_0
    port( b4_nUAi           : in    std_logic_vector(206 downto 204) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_70_0
    port( b4_nUAi           : in    std_logic_vector(293 downto 291) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_94_0
    port( b4_nUAi           : in    std_logic_vector(221 downto 219) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_154_0
    port( b4_nUAi           : in    std_logic_vector(41 downto 39) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_124_0
    port( b4_nUAi           : in    std_logic_vector(131 downto 129) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_10_0
    port( b4_nUAi           : in    std_logic_vector(473 downto 471) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_42_0
    port( b4_nUAi           : in    std_logic_vector(377 downto 375) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_114_0
    port( b4_nUAi           : in    std_logic_vector(161 downto 159) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_138_0
    port( b4_nUAi           : in    std_logic_vector(89 downto 87) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_17_0
    port( b4_nUAi           : in    std_logic_vector(452 downto 450) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_98_0
    port( b4_nUAi           : in    std_logic_vector(209 downto 207) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_121_0
    port( b4_nUAi           : in    std_logic_vector(140 downto 138) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_38_0
    port( b4_nUAi           : in    std_logic_vector(389 downto 387) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

  component b8_1LbcQDr1_x_82_0
    port( b4_nUAi           : in    std_logic_vector(257 downto 255) := (others => 'U');
          b6_2ZTGIf_0       : out   std_logic;
          b11_OFWNT9L_8tZ_0 : in    std_logic := 'U';
          mdiclink_reg_0    : in    std_logic := 'U'
        );
  end component;

    signal \b6_2ZTGIf[0]\, \b6_2ZTGIf[1]\, \b6_2ZTGIf[2]\, 
        \b6_2ZTGIf[3]\, \b6_2ZTGIf[4]\, \b6_2ZTGIf[5]\, 
        \b6_2ZTGIf[6]\, \b6_2ZTGIf[7]\, \b6_2ZTGIf[8]\, 
        \b6_2ZTGIf[9]\, \b6_2ZTGIf[10]\, \b6_2ZTGIf[11]\, 
        \b6_2ZTGIf[12]\, \b6_2ZTGIf[13]\, \b6_2ZTGIf[14]\, 
        \b6_2ZTGIf[15]\, \b6_2ZTGIf[16]\, \b6_2ZTGIf[17]\, 
        \b6_2ZTGIf[18]\, \b6_2ZTGIf[19]\, \b6_2ZTGIf[20]\, 
        \b6_2ZTGIf[21]\, \b6_2ZTGIf[22]\, \b6_2ZTGIf[23]\, 
        \b6_2ZTGIf[24]\, \b6_2ZTGIf[25]\, \b6_2ZTGIf[26]\, 
        \b6_2ZTGIf[27]\, \b6_2ZTGIf[28]\, \b6_2ZTGIf[29]\, 
        \b6_2ZTGIf[30]\, \b6_2ZTGIf[31]\, \b6_2ZTGIf[32]\, 
        \b6_2ZTGIf[33]\, \b6_2ZTGIf[34]\, \b6_2ZTGIf[35]\, 
        \b6_2ZTGIf[36]\, \b6_2ZTGIf[37]\, \b6_2ZTGIf[38]\, 
        \b6_2ZTGIf[39]\, \b6_2ZTGIf[40]\, \b6_2ZTGIf[41]\, 
        \b6_2ZTGIf[42]\, \b6_2ZTGIf[43]\, \b6_2ZTGIf[44]\, 
        \b6_2ZTGIf[45]\, \b6_2ZTGIf[46]\, \b6_2ZTGIf[47]\, 
        \b6_2ZTGIf[48]\, \b6_2ZTGIf[49]\, \b6_2ZTGIf[50]\, 
        \b6_2ZTGIf[51]\, \b6_2ZTGIf[52]\, \b6_2ZTGIf[53]\, 
        \b6_2ZTGIf[54]\, \b6_2ZTGIf[55]\, \b6_2ZTGIf[56]\, 
        \b6_2ZTGIf[57]\, \b6_2ZTGIf[58]\, \b6_2ZTGIf[59]\, 
        \b6_2ZTGIf[60]\, \b6_2ZTGIf[61]\, \b6_2ZTGIf[62]\, 
        \b6_2ZTGIf[63]\, \b6_2ZTGIf[64]\, \b6_2ZTGIf[65]\, 
        \b6_2ZTGIf[66]\, \b6_2ZTGIf[67]\, \b6_2ZTGIf[68]\, 
        \b6_2ZTGIf[69]\, \b6_2ZTGIf[70]\, \b6_2ZTGIf[71]\, 
        \b6_2ZTGIf[72]\, \b6_2ZTGIf[73]\, \b6_2ZTGIf[74]\, 
        \b6_2ZTGIf[75]\, \b6_2ZTGIf[76]\, \b6_2ZTGIf[77]\, 
        \b6_2ZTGIf[78]\, \b6_2ZTGIf[79]\, \b6_2ZTGIf[80]\, 
        \b6_2ZTGIf[81]\, \b6_2ZTGIf[82]\, \b6_2ZTGIf[83]\, 
        \b6_2ZTGIf[84]\, \b6_2ZTGIf[85]\, \b6_2ZTGIf[86]\, 
        \b6_2ZTGIf[87]\, \b6_2ZTGIf[88]\, \b6_2ZTGIf[89]\, 
        \b6_2ZTGIf[90]\, \b6_2ZTGIf[91]\, \b6_2ZTGIf[92]\, 
        \b6_2ZTGIf[93]\, \b6_2ZTGIf[94]\, \b6_2ZTGIf[95]\, 
        \b6_2ZTGIf[96]\, \b6_2ZTGIf[97]\, \b6_2ZTGIf[98]\, 
        \b6_2ZTGIf[99]\, \b6_2ZTGIf[100]\, \b6_2ZTGIf[101]\, 
        \b6_2ZTGIf[102]\, \b6_2ZTGIf[103]\, \b6_2ZTGIf[104]\, 
        \b6_2ZTGIf[105]\, \b6_2ZTGIf[106]\, \b6_2ZTGIf[107]\, 
        \b6_2ZTGIf[108]\, \b6_2ZTGIf[109]\, \b6_2ZTGIf[110]\, 
        \b6_2ZTGIf[111]\, \b6_2ZTGIf[112]\, \b6_2ZTGIf[113]\, 
        \b6_2ZTGIf[114]\, \b6_2ZTGIf[115]\, \b6_2ZTGIf[116]\, 
        \b6_2ZTGIf[117]\, \b6_2ZTGIf[118]\, \b6_2ZTGIf[119]\, 
        \b6_2ZTGIf[120]\, \b6_2ZTGIf[121]\, \b6_2ZTGIf[122]\, 
        \b6_2ZTGIf[123]\, \b6_2ZTGIf[124]\, \b6_2ZTGIf[125]\, 
        \b6_2ZTGIf[126]\, \b6_2ZTGIf[127]\, \b6_2ZTGIf[128]\, 
        \b6_2ZTGIf[129]\, \b6_2ZTGIf[130]\, \b6_2ZTGIf[131]\, 
        \b6_2ZTGIf[132]\, \b6_2ZTGIf[133]\, \b6_2ZTGIf[134]\, 
        \b6_2ZTGIf[135]\, \b6_2ZTGIf[136]\, \b6_2ZTGIf[137]\, 
        \b6_2ZTGIf[138]\, \b6_2ZTGIf[139]\, \b6_2ZTGIf[140]\, 
        \b6_2ZTGIf[141]\, \b6_2ZTGIf[142]\, \b6_2ZTGIf[143]\, 
        \b6_2ZTGIf[144]\, \b6_2ZTGIf[145]\, \b6_2ZTGIf[146]\, 
        \b6_2ZTGIf[147]\, \b6_2ZTGIf[148]\, \b6_2ZTGIf[149]\, 
        \b6_2ZTGIf[150]\, \b6_2ZTGIf[151]\, \b6_2ZTGIf[152]\, 
        \b6_2ZTGIf[153]\, \b6_2ZTGIf[154]\, \b6_2ZTGIf[155]\, 
        \b6_2ZTGIf[156]\, \b6_2ZTGIf[157]\, \b6_2ZTGIf[158]\, 
        \b6_2ZTGIf[159]\, \b6_2ZTGIf[160]\, \b6_2ZTGIf[161]\, 
        \b6_2ZTGIf[162]\, \b6_2ZTGIf[163]\, \b6_2ZTGIf[164]\, 
        \b6_2ZTGIf[165]\, \b6_2ZTGIf[166]\, \b6_2ZTGIf[167]\, 
        GND_net_1, VCC_net_1 : std_logic;

    for all : b8_1LbcQDr1_x_39_0
	Use entity work.b8_1LbcQDr1_x_39_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_93_0
	Use entity work.b8_1LbcQDr1_x_93_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_16_0
	Use entity work.b8_1LbcQDr1_x_16_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_40_0
	Use entity work.b8_1LbcQDr1_x_40_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_153_0
	Use entity work.b8_1LbcQDr1_x_153_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_96_0
	Use entity work.b8_1LbcQDr1_x_96_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_156_0
	Use entity work.b8_1LbcQDr1_x_156_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_47_0
	Use entity work.b8_1LbcQDr1_x_47_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_97_0
	Use entity work.b8_1LbcQDr1_x_97_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_157_0
	Use entity work.b8_1LbcQDr1_x_157_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_116_0
	Use entity work.b8_1LbcQDr1_x_116_0(DEF_ARCH);
    for all : b16_CRGcTCua_eH4_uaL_x_0
	Use entity work.b16_CRGcTCua_eH4_uaL_x_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_117_0
	Use entity work.b8_1LbcQDr1_x_117_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_85_0
	Use entity work.b8_1LbcQDr1_x_85_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_46_0
	Use entity work.b8_1LbcQDr1_x_46_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_142_0
	Use entity work.b8_1LbcQDr1_x_142_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_102_0
	Use entity work.b8_1LbcQDr1_x_102_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_133_0
	Use entity work.b8_1LbcQDr1_x_133_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_3_0
	Use entity work.b8_1LbcQDr1_x_3_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_1_0
	Use entity work.b8_1LbcQDr1_x_1_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_103_0
	Use entity work.b8_1LbcQDr1_x_103_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_23_0
	Use entity work.b8_1LbcQDr1_x_23_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_21_0
	Use entity work.b8_1LbcQDr1_x_21_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_14_0
	Use entity work.b8_1LbcQDr1_x_14_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_143_0
	Use entity work.b8_1LbcQDr1_x_143_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_145_0
	Use entity work.b8_1LbcQDr1_x_145_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_105_0
	Use entity work.b8_1LbcQDr1_x_105_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_126_0
	Use entity work.b8_1LbcQDr1_x_126_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_89_0
	Use entity work.b8_1LbcQDr1_x_89_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_149_0
	Use entity work.b8_1LbcQDr1_x_149_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_80_0
	Use entity work.b8_1LbcQDr1_x_80_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_127_0
	Use entity work.b8_1LbcQDr1_x_127_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_131_0
	Use entity work.b8_1LbcQDr1_x_131_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_109_0
	Use entity work.b8_1LbcQDr1_x_109_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_44_0
	Use entity work.b8_1LbcQDr1_x_44_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_88_0
	Use entity work.b8_1LbcQDr1_x_88_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_148_0
	Use entity work.b8_1LbcQDr1_x_148_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_33_0
	Use entity work.b8_1LbcQDr1_x_33_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_108_0
	Use entity work.b8_1LbcQDr1_x_108_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_163_0
	Use entity work.b8_1LbcQDr1_x_163_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_31_0
	Use entity work.b8_1LbcQDr1_x_31_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_140_0
	Use entity work.b8_1LbcQDr1_x_140_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_100_0
	Use entity work.b8_1LbcQDr1_x_100_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_53_0
	Use entity work.b8_1LbcQDr1_x_53_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_71_0
	Use entity work.b8_1LbcQDr1_x_71_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_51_0
	Use entity work.b8_1LbcQDr1_x_51_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_63_0
	Use entity work.b8_1LbcQDr1_x_63_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_134_0
	Use entity work.b8_1LbcQDr1_x_134_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_61_0
	Use entity work.b8_1LbcQDr1_x_61_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_119_0
	Use entity work.b8_1LbcQDr1_x_119_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_92_0
	Use entity work.b8_1LbcQDr1_x_92_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_152_0
	Use entity work.b8_1LbcQDr1_x_152_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_160_0
	Use entity work.b8_1LbcQDr1_x_160_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_112_0
	Use entity work.b8_1LbcQDr1_x_112_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_118_0
	Use entity work.b8_1LbcQDr1_x_118_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_136_0
	Use entity work.b8_1LbcQDr1_x_136_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_95_0
	Use entity work.b8_1LbcQDr1_x_95_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_155_0
	Use entity work.b8_1LbcQDr1_x_155_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_137_0
	Use entity work.b8_1LbcQDr1_x_137_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_5_0
	Use entity work.b8_1LbcQDr1_x_5_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_115_0
	Use entity work.b8_1LbcQDr1_x_115_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_25_0
	Use entity work.b8_1LbcQDr1_x_25_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_74_0
	Use entity work.b8_1LbcQDr1_x_74_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_161_0
	Use entity work.b8_1LbcQDr1_x_161_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_2_0
	Use entity work.b8_1LbcQDr1_x_2_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_22_0
	Use entity work.b8_1LbcQDr1_x_22_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_122_0
	Use entity work.b8_1LbcQDr1_x_122_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_18_0
	Use entity work.b8_1LbcQDr1_x_18_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_0_0
	Use entity work.b8_1LbcQDr1_x_0_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_76_0
	Use entity work.b8_1LbcQDr1_x_76_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_162_0
	Use entity work.b8_1LbcQDr1_x_162_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_19_0
	Use entity work.b8_1LbcQDr1_x_19_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_77_0
	Use entity work.b8_1LbcQDr1_x_77_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_7_0
	Use entity work.b8_1LbcQDr1_x_7_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_35_0
	Use entity work.b8_1LbcQDr1_x_35_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_20_0
	Use entity work.b8_1LbcQDr1_x_20_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_90_0
	Use entity work.b8_1LbcQDr1_x_90_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_150_0
	Use entity work.b8_1LbcQDr1_x_150_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_113_0
	Use entity work.b8_1LbcQDr1_x_113_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_165_0
	Use entity work.b8_1LbcQDr1_x_165_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_110_0
	Use entity work.b8_1LbcQDr1_x_110_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_27_0
	Use entity work.b8_1LbcQDr1_x_27_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_129_0
	Use entity work.b8_1LbcQDr1_x_129_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_81_0
	Use entity work.b8_1LbcQDr1_x_81_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_125_0
	Use entity work.b8_1LbcQDr1_x_125_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_6_0
	Use entity work.b8_1LbcQDr1_x_6_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_32_0
	Use entity work.b8_1LbcQDr1_x_32_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_128_0
	Use entity work.b8_1LbcQDr1_x_128_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_26_0
	Use entity work.b8_1LbcQDr1_x_26_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_28_0
	Use entity work.b8_1LbcQDr1_x_28_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_55_0
	Use entity work.b8_1LbcQDr1_x_55_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_13_0
	Use entity work.b8_1LbcQDr1_x_13_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_65_0
	Use entity work.b8_1LbcQDr1_x_65_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_29_0
	Use entity work.b8_1LbcQDr1_x_29_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_11_0
	Use entity work.b8_1LbcQDr1_x_11_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_30_0
	Use entity work.b8_1LbcQDr1_x_30_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_141_0
	Use entity work.b8_1LbcQDr1_x_141_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_167_0
	Use entity work.b8_1LbcQDr1_x_167_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_37_0
	Use entity work.b8_1LbcQDr1_x_37_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_101_0
	Use entity work.b8_1LbcQDr1_x_101_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_52_0
	Use entity work.b8_1LbcQDr1_x_52_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_62_0
	Use entity work.b8_1LbcQDr1_x_62_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_69_0
	Use entity work.b8_1LbcQDr1_x_69_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_84_0
	Use entity work.b8_1LbcQDr1_x_84_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_43_0
	Use entity work.b8_1LbcQDr1_x_43_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_120_0
	Use entity work.b8_1LbcQDr1_x_120_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_48_0
	Use entity work.b8_1LbcQDr1_x_48_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_41_0
	Use entity work.b8_1LbcQDr1_x_41_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_36_0
	Use entity work.b8_1LbcQDr1_x_36_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_58_0
	Use entity work.b8_1LbcQDr1_x_58_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_4_0
	Use entity work.b8_1LbcQDr1_x_4_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_49_0
	Use entity work.b8_1LbcQDr1_x_49_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_68_0
	Use entity work.b8_1LbcQDr1_x_68_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_132_0
	Use entity work.b8_1LbcQDr1_x_132_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_59_0
	Use entity work.b8_1LbcQDr1_x_59_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_164_0
	Use entity work.b8_1LbcQDr1_x_164_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_50_0
	Use entity work.b8_1LbcQDr1_x_50_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_24_0
	Use entity work.b8_1LbcQDr1_x_24_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_60_0
	Use entity work.b8_1LbcQDr1_x_60_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_57_0
	Use entity work.b8_1LbcQDr1_x_57_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_67_0
	Use entity work.b8_1LbcQDr1_x_67_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_86_0
	Use entity work.b8_1LbcQDr1_x_86_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_87_0
	Use entity work.b8_1LbcQDr1_x_87_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_135_0
	Use entity work.b8_1LbcQDr1_x_135_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_56_0
	Use entity work.b8_1LbcQDr1_x_56_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_144_0
	Use entity work.b8_1LbcQDr1_x_144_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_104_0
	Use entity work.b8_1LbcQDr1_x_104_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_66_0
	Use entity work.b8_1LbcQDr1_x_66_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_34_0
	Use entity work.b8_1LbcQDr1_x_34_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_72_0
	Use entity work.b8_1LbcQDr1_x_72_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_159_0
	Use entity work.b8_1LbcQDr1_x_159_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_146_0
	Use entity work.b8_1LbcQDr1_x_146_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_106_0
	Use entity work.b8_1LbcQDr1_x_106_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_147_0
	Use entity work.b8_1LbcQDr1_x_147_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_107_0
	Use entity work.b8_1LbcQDr1_x_107_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_75_0
	Use entity work.b8_1LbcQDr1_x_75_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_91_0
	Use entity work.b8_1LbcQDr1_x_91_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_151_0
	Use entity work.b8_1LbcQDr1_x_151_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_123_0
	Use entity work.b8_1LbcQDr1_x_123_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_130_0
	Use entity work.b8_1LbcQDr1_x_130_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_54_0
	Use entity work.b8_1LbcQDr1_x_54_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_79_0
	Use entity work.b8_1LbcQDr1_x_79_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_64_0
	Use entity work.b8_1LbcQDr1_x_64_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_111_0
	Use entity work.b8_1LbcQDr1_x_111_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_83_0
	Use entity work.b8_1LbcQDr1_x_83_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_15_0
	Use entity work.b8_1LbcQDr1_x_15_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_78_0
	Use entity work.b8_1LbcQDr1_x_78_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_166_0
	Use entity work.b8_1LbcQDr1_x_166_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_12_0
	Use entity work.b8_1LbcQDr1_x_12_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_73_0
	Use entity work.b8_1LbcQDr1_x_73_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_45_0
	Use entity work.b8_1LbcQDr1_x_45_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_158_0
	Use entity work.b8_1LbcQDr1_x_158_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_8_0
	Use entity work.b8_1LbcQDr1_x_8_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_139_0
	Use entity work.b8_1LbcQDr1_x_139_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_9_0
	Use entity work.b8_1LbcQDr1_x_9_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_99_0
	Use entity work.b8_1LbcQDr1_x_99_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_70_0
	Use entity work.b8_1LbcQDr1_x_70_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_94_0
	Use entity work.b8_1LbcQDr1_x_94_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_154_0
	Use entity work.b8_1LbcQDr1_x_154_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_124_0
	Use entity work.b8_1LbcQDr1_x_124_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_10_0
	Use entity work.b8_1LbcQDr1_x_10_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_42_0
	Use entity work.b8_1LbcQDr1_x_42_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_114_0
	Use entity work.b8_1LbcQDr1_x_114_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_138_0
	Use entity work.b8_1LbcQDr1_x_138_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_17_0
	Use entity work.b8_1LbcQDr1_x_17_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_98_0
	Use entity work.b8_1LbcQDr1_x_98_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_121_0
	Use entity work.b8_1LbcQDr1_x_121_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_38_0
	Use entity work.b8_1LbcQDr1_x_38_0(DEF_ARCH);
    for all : b8_1LbcQDr1_x_82_0
	Use entity work.b8_1LbcQDr1_x_82_0(DEF_ARCH);
begin 


    b9_1LbcgKGIS : b8_1LbcQDr1_x_39_0
      port map(b4_nUAi(386) => b4_nUAi(386), b4_nUAi(385) => 
        b4_nUAi(385), b4_nUAi(384) => b4_nUAi(384), b6_2ZTGIf_0
         => \b6_2ZTGIf[128]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(17), mdiclink_reg_0 => mdiclink_reg(150));
    
    b8_1LbcgKxQ0 : b8_1LbcQDr1_x_93_0
      port map(b4_nUAi(224) => b4_nUAi(224), b4_nUAi(223) => 
        b4_nUAi(223), b4_nUAi(222) => b4_nUAi(222), b6_2ZTGIf_0
         => \b6_2ZTGIf[74]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(149), mdiclink_reg_0 => mdiclink_reg(18));
    
    b9_1LbcgKGUn : b8_1LbcQDr1_x_16_0
      port map(b4_nUAi(455) => b4_nUAi(455), b4_nUAi(454) => 
        b4_nUAi(454), b4_nUAi(453) => b4_nUAi(453), b6_2ZTGIf_0
         => \b6_2ZTGIf[151]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(8), mdiclink_reg_0 => mdiclink_reg(159));
    
    b9_1LbcgKGIe : b8_1LbcQDr1_x_40_0
      port map(b4_nUAi(383) => b4_nUAi(383), b4_nUAi(382) => 
        b4_nUAi(382), b4_nUAi(381) => b4_nUAi(381), b6_2ZTGIf_0
         => \b6_2ZTGIf[127]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(18), mdiclink_reg_0 => mdiclink_reg(149));
    
    b8_1LbcgKGQ0 : b8_1LbcQDr1_x_153_0
      port map(b4_nUAi(44) => b4_nUAi(44), b4_nUAi(43) => 
        b4_nUAi(43), b4_nUAi(42) => b4_nUAi(42), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[14]\, b11_OFWNT9L_8tZ_0 => b11_OFWNT9L_8tZ(80), 
        mdiclink_reg_0 => mdiclink_reg(87));
    
    b8_1LbcgKxS : b8_1LbcQDr1_x_96_0
      port map(b4_nUAi(215) => b4_nUAi(215), b4_nUAi(214) => 
        b4_nUAi(214), b4_nUAi(213) => b4_nUAi(213), b6_2ZTGIf_0
         => \b6_2ZTGIf[71]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(152), mdiclink_reg_0 => mdiclink_reg(15));
    
    b8_1LbcgKGS : b8_1LbcQDr1_x_156_0
      port map(b4_nUAi(35) => b4_nUAi(35), b4_nUAi(34) => 
        b4_nUAi(34), b4_nUAi(33) => b4_nUAi(33), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[11]\, b11_OFWNT9L_8tZ_0 => b11_OFWNT9L_8tZ(95), 
        mdiclink_reg_0 => mdiclink_reg(72));
    
    b9_1LbcgKGIm : b8_1LbcQDr1_x_47_0
      port map(b4_nUAi(362) => b4_nUAi(362), b4_nUAi(361) => 
        b4_nUAi(361), b4_nUAi(360) => b4_nUAi(360), b6_2ZTGIf_0
         => \b6_2ZTGIf[120]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(33), mdiclink_reg_0 => mdiclink_reg(134));
    
    b8_1LbcgKxR : b8_1LbcQDr1_x_97_0
      port map(b4_nUAi(212) => b4_nUAi(212), b4_nUAi(211) => 
        b4_nUAi(211), b4_nUAi(210) => b4_nUAi(210), b6_2ZTGIf_0
         => \b6_2ZTGIf[70]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(153), mdiclink_reg_0 => mdiclink_reg(14));
    
    b8_1LbcgKGR : b8_1LbcQDr1_x_157_0
      port map(b4_nUAi(32) => b4_nUAi(32), b4_nUAi(31) => 
        b4_nUAi(31), b4_nUAi(30) => b4_nUAi(30), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[10]\, b11_OFWNT9L_8tZ_0 => b11_OFWNT9L_8tZ(96), 
        mdiclink_reg_0 => mdiclink_reg(71));
    
    b8_1LbcgKIS : b8_1LbcQDr1_x_116_0
      port map(b4_nUAi(155) => b4_nUAi(155), b4_nUAi(154) => 
        b4_nUAi(154), b4_nUAi(153) => b4_nUAi(153), b6_2ZTGIf_0
         => \b6_2ZTGIf[51]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(67), mdiclink_reg_0 => mdiclink_reg(100));
    
    b6_2ZGFQ9 : b16_CRGcTCua_eH4_uaL_x_0
      port map(b6_2ZTGIf(167) => \b6_2ZTGIf[167]\, b6_2ZTGIf(166)
         => \b6_2ZTGIf[166]\, b6_2ZTGIf(165) => \b6_2ZTGIf[165]\, 
        b6_2ZTGIf(164) => \b6_2ZTGIf[164]\, b6_2ZTGIf(163) => 
        \b6_2ZTGIf[163]\, b6_2ZTGIf(162) => \b6_2ZTGIf[162]\, 
        b6_2ZTGIf(161) => \b6_2ZTGIf[161]\, b6_2ZTGIf(160) => 
        \b6_2ZTGIf[160]\, b6_2ZTGIf(159) => \b6_2ZTGIf[159]\, 
        b6_2ZTGIf(158) => \b6_2ZTGIf[158]\, b6_2ZTGIf(157) => 
        \b6_2ZTGIf[157]\, b6_2ZTGIf(156) => \b6_2ZTGIf[156]\, 
        b6_2ZTGIf(155) => \b6_2ZTGIf[155]\, b6_2ZTGIf(154) => 
        \b6_2ZTGIf[154]\, b6_2ZTGIf(153) => \b6_2ZTGIf[153]\, 
        b6_2ZTGIf(152) => \b6_2ZTGIf[152]\, b6_2ZTGIf(151) => 
        \b6_2ZTGIf[151]\, b6_2ZTGIf(150) => \b6_2ZTGIf[150]\, 
        b6_2ZTGIf(149) => \b6_2ZTGIf[149]\, b6_2ZTGIf(148) => 
        \b6_2ZTGIf[148]\, b6_2ZTGIf(147) => \b6_2ZTGIf[147]\, 
        b6_2ZTGIf(146) => \b6_2ZTGIf[146]\, b6_2ZTGIf(145) => 
        \b6_2ZTGIf[145]\, b6_2ZTGIf(144) => \b6_2ZTGIf[144]\, 
        b6_2ZTGIf(143) => \b6_2ZTGIf[143]\, b6_2ZTGIf(142) => 
        \b6_2ZTGIf[142]\, b6_2ZTGIf(141) => \b6_2ZTGIf[141]\, 
        b6_2ZTGIf(140) => \b6_2ZTGIf[140]\, b6_2ZTGIf(139) => 
        \b6_2ZTGIf[139]\, b6_2ZTGIf(138) => \b6_2ZTGIf[138]\, 
        b6_2ZTGIf(137) => \b6_2ZTGIf[137]\, b6_2ZTGIf(136) => 
        \b6_2ZTGIf[136]\, b6_2ZTGIf(135) => \b6_2ZTGIf[135]\, 
        b6_2ZTGIf(134) => \b6_2ZTGIf[134]\, b6_2ZTGIf(133) => 
        \b6_2ZTGIf[133]\, b6_2ZTGIf(132) => \b6_2ZTGIf[132]\, 
        b6_2ZTGIf(131) => \b6_2ZTGIf[131]\, b6_2ZTGIf(130) => 
        \b6_2ZTGIf[130]\, b6_2ZTGIf(129) => \b6_2ZTGIf[129]\, 
        b6_2ZTGIf(128) => \b6_2ZTGIf[128]\, b6_2ZTGIf(127) => 
        \b6_2ZTGIf[127]\, b6_2ZTGIf(126) => \b6_2ZTGIf[126]\, 
        b6_2ZTGIf(125) => \b6_2ZTGIf[125]\, b6_2ZTGIf(124) => 
        \b6_2ZTGIf[124]\, b6_2ZTGIf(123) => \b6_2ZTGIf[123]\, 
        b6_2ZTGIf(122) => \b6_2ZTGIf[122]\, b6_2ZTGIf(121) => 
        \b6_2ZTGIf[121]\, b6_2ZTGIf(120) => \b6_2ZTGIf[120]\, 
        b6_2ZTGIf(119) => \b6_2ZTGIf[119]\, b6_2ZTGIf(118) => 
        \b6_2ZTGIf[118]\, b6_2ZTGIf(117) => \b6_2ZTGIf[117]\, 
        b6_2ZTGIf(116) => \b6_2ZTGIf[116]\, b6_2ZTGIf(115) => 
        \b6_2ZTGIf[115]\, b6_2ZTGIf(114) => \b6_2ZTGIf[114]\, 
        b6_2ZTGIf(113) => \b6_2ZTGIf[113]\, b6_2ZTGIf(112) => 
        \b6_2ZTGIf[112]\, b6_2ZTGIf(111) => \b6_2ZTGIf[111]\, 
        b6_2ZTGIf(110) => \b6_2ZTGIf[110]\, b6_2ZTGIf(109) => 
        \b6_2ZTGIf[109]\, b6_2ZTGIf(108) => \b6_2ZTGIf[108]\, 
        b6_2ZTGIf(107) => \b6_2ZTGIf[107]\, b6_2ZTGIf(106) => 
        \b6_2ZTGIf[106]\, b6_2ZTGIf(105) => \b6_2ZTGIf[105]\, 
        b6_2ZTGIf(104) => \b6_2ZTGIf[104]\, b6_2ZTGIf(103) => 
        \b6_2ZTGIf[103]\, b6_2ZTGIf(102) => \b6_2ZTGIf[102]\, 
        b6_2ZTGIf(101) => \b6_2ZTGIf[101]\, b6_2ZTGIf(100) => 
        \b6_2ZTGIf[100]\, b6_2ZTGIf(99) => \b6_2ZTGIf[99]\, 
        b6_2ZTGIf(98) => \b6_2ZTGIf[98]\, b6_2ZTGIf(97) => 
        \b6_2ZTGIf[97]\, b6_2ZTGIf(96) => \b6_2ZTGIf[96]\, 
        b6_2ZTGIf(95) => \b6_2ZTGIf[95]\, b6_2ZTGIf(94) => 
        \b6_2ZTGIf[94]\, b6_2ZTGIf(93) => \b6_2ZTGIf[93]\, 
        b6_2ZTGIf(92) => \b6_2ZTGIf[92]\, b6_2ZTGIf(91) => 
        \b6_2ZTGIf[91]\, b6_2ZTGIf(90) => \b6_2ZTGIf[90]\, 
        b6_2ZTGIf(89) => \b6_2ZTGIf[89]\, b6_2ZTGIf(88) => 
        \b6_2ZTGIf[88]\, b6_2ZTGIf(87) => \b6_2ZTGIf[87]\, 
        b6_2ZTGIf(86) => \b6_2ZTGIf[86]\, b6_2ZTGIf(85) => 
        \b6_2ZTGIf[85]\, b6_2ZTGIf(84) => \b6_2ZTGIf[84]\, 
        b6_2ZTGIf(83) => \b6_2ZTGIf[83]\, b6_2ZTGIf(82) => 
        \b6_2ZTGIf[82]\, b6_2ZTGIf(81) => \b6_2ZTGIf[81]\, 
        b6_2ZTGIf(80) => \b6_2ZTGIf[80]\, b6_2ZTGIf(79) => 
        \b6_2ZTGIf[79]\, b6_2ZTGIf(78) => \b6_2ZTGIf[78]\, 
        b6_2ZTGIf(77) => \b6_2ZTGIf[77]\, b6_2ZTGIf(76) => 
        \b6_2ZTGIf[76]\, b6_2ZTGIf(75) => \b6_2ZTGIf[75]\, 
        b6_2ZTGIf(74) => \b6_2ZTGIf[74]\, b6_2ZTGIf(73) => 
        \b6_2ZTGIf[73]\, b6_2ZTGIf(72) => \b6_2ZTGIf[72]\, 
        b6_2ZTGIf(71) => \b6_2ZTGIf[71]\, b6_2ZTGIf(70) => 
        \b6_2ZTGIf[70]\, b6_2ZTGIf(69) => \b6_2ZTGIf[69]\, 
        b6_2ZTGIf(68) => \b6_2ZTGIf[68]\, b6_2ZTGIf(67) => 
        \b6_2ZTGIf[67]\, b6_2ZTGIf(66) => \b6_2ZTGIf[66]\, 
        b6_2ZTGIf(65) => \b6_2ZTGIf[65]\, b6_2ZTGIf(64) => 
        \b6_2ZTGIf[64]\, b6_2ZTGIf(63) => \b6_2ZTGIf[63]\, 
        b6_2ZTGIf(62) => \b6_2ZTGIf[62]\, b6_2ZTGIf(61) => 
        \b6_2ZTGIf[61]\, b6_2ZTGIf(60) => \b6_2ZTGIf[60]\, 
        b6_2ZTGIf(59) => \b6_2ZTGIf[59]\, b6_2ZTGIf(58) => 
        \b6_2ZTGIf[58]\, b6_2ZTGIf(57) => \b6_2ZTGIf[57]\, 
        b6_2ZTGIf(56) => \b6_2ZTGIf[56]\, b6_2ZTGIf(55) => 
        \b6_2ZTGIf[55]\, b6_2ZTGIf(54) => \b6_2ZTGIf[54]\, 
        b6_2ZTGIf(53) => \b6_2ZTGIf[53]\, b6_2ZTGIf(52) => 
        \b6_2ZTGIf[52]\, b6_2ZTGIf(51) => \b6_2ZTGIf[51]\, 
        b6_2ZTGIf(50) => \b6_2ZTGIf[50]\, b6_2ZTGIf(49) => 
        \b6_2ZTGIf[49]\, b6_2ZTGIf(48) => \b6_2ZTGIf[48]\, 
        b6_2ZTGIf(47) => \b6_2ZTGIf[47]\, b6_2ZTGIf(46) => 
        \b6_2ZTGIf[46]\, b6_2ZTGIf(45) => \b6_2ZTGIf[45]\, 
        b6_2ZTGIf(44) => \b6_2ZTGIf[44]\, b6_2ZTGIf(43) => 
        \b6_2ZTGIf[43]\, b6_2ZTGIf(42) => \b6_2ZTGIf[42]\, 
        b6_2ZTGIf(41) => \b6_2ZTGIf[41]\, b6_2ZTGIf(40) => 
        \b6_2ZTGIf[40]\, b6_2ZTGIf(39) => \b6_2ZTGIf[39]\, 
        b6_2ZTGIf(38) => \b6_2ZTGIf[38]\, b6_2ZTGIf(37) => 
        \b6_2ZTGIf[37]\, b6_2ZTGIf(36) => \b6_2ZTGIf[36]\, 
        b6_2ZTGIf(35) => \b6_2ZTGIf[35]\, b6_2ZTGIf(34) => 
        \b6_2ZTGIf[34]\, b6_2ZTGIf(33) => \b6_2ZTGIf[33]\, 
        b6_2ZTGIf(32) => \b6_2ZTGIf[32]\, b6_2ZTGIf(31) => 
        \b6_2ZTGIf[31]\, b6_2ZTGIf(30) => \b6_2ZTGIf[30]\, 
        b6_2ZTGIf(29) => \b6_2ZTGIf[29]\, b6_2ZTGIf(28) => 
        \b6_2ZTGIf[28]\, b6_2ZTGIf(27) => \b6_2ZTGIf[27]\, 
        b6_2ZTGIf(26) => \b6_2ZTGIf[26]\, b6_2ZTGIf(25) => 
        \b6_2ZTGIf[25]\, b6_2ZTGIf(24) => \b6_2ZTGIf[24]\, 
        b6_2ZTGIf(23) => \b6_2ZTGIf[23]\, b6_2ZTGIf(22) => 
        \b6_2ZTGIf[22]\, b6_2ZTGIf(21) => \b6_2ZTGIf[21]\, 
        b6_2ZTGIf(20) => \b6_2ZTGIf[20]\, b6_2ZTGIf(19) => 
        \b6_2ZTGIf[19]\, b6_2ZTGIf(18) => \b6_2ZTGIf[18]\, 
        b6_2ZTGIf(17) => \b6_2ZTGIf[17]\, b6_2ZTGIf(16) => 
        \b6_2ZTGIf[16]\, b6_2ZTGIf(15) => \b6_2ZTGIf[15]\, 
        b6_2ZTGIf(14) => \b6_2ZTGIf[14]\, b6_2ZTGIf(13) => 
        \b6_2ZTGIf[13]\, b6_2ZTGIf(12) => \b6_2ZTGIf[12]\, 
        b6_2ZTGIf(11) => \b6_2ZTGIf[11]\, b6_2ZTGIf(10) => 
        \b6_2ZTGIf[10]\, b6_2ZTGIf(9) => \b6_2ZTGIf[9]\, 
        b6_2ZTGIf(8) => \b6_2ZTGIf[8]\, b6_2ZTGIf(7) => 
        \b6_2ZTGIf[7]\, b6_2ZTGIf(6) => \b6_2ZTGIf[6]\, 
        b6_2ZTGIf(5) => \b6_2ZTGIf[5]\, b6_2ZTGIf(4) => 
        \b6_2ZTGIf[4]\, b6_2ZTGIf(3) => \b6_2ZTGIf[3]\, 
        b6_2ZTGIf(2) => \b6_2ZTGIf[2]\, b6_2ZTGIf(1) => 
        \b6_2ZTGIf[1]\, b6_2ZTGIf(0) => \b6_2ZTGIf[0]\, 
        b10_nYBzIXrKbK_0 => b10_nYBzIXrKbK_0, CommsFPGA_CCC_0_GL0
         => CommsFPGA_CCC_0_GL0);
    
    b8_1LbcgKIR : b8_1LbcQDr1_x_117_0
      port map(b4_nUAi(152) => b4_nUAi(152), b4_nUAi(151) => 
        b4_nUAi(151), b4_nUAi(150) => b4_nUAi(150), b6_2ZTGIf_0
         => \b6_2ZTGIf[50]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(68), mdiclink_reg_0 => mdiclink_reg(99));
    
    b8_1LbcgKbI : b8_1LbcQDr1_x_85_0
      port map(b4_nUAi(248) => b4_nUAi(248), b4_nUAi(247) => 
        b4_nUAi(247), b4_nUAi(246) => b4_nUAi(246), b6_2ZTGIf_0
         => \b6_2ZTGIf[82]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(140), mdiclink_reg_0 => mdiclink_reg(27));
    
    b9_1LbcgKGIn : b8_1LbcQDr1_x_46_0
      port map(b4_nUAi(365) => b4_nUAi(365), b4_nUAi(364) => 
        b4_nUAi(364), b4_nUAi(363) => b4_nUAi(363), b6_2ZTGIf_0
         => \b6_2ZTGIf[121]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(32), mdiclink_reg_0 => mdiclink_reg(135));
    
    b8_1LbcgKwU : b8_1LbcQDr1_x_142_0
      port map(b4_nUAi(77) => b4_nUAi(77), b4_nUAi(76) => 
        b4_nUAi(76), b4_nUAi(75) => b4_nUAi(75), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[25]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(163), mdiclink_reg_0 => mdiclink_reg(4));
    
    b8_1LbcgKoU : b8_1LbcQDr1_x_102_0
      port map(b4_nUAi(197) => b4_nUAi(197), b4_nUAi(196) => 
        b4_nUAi(196), b4_nUAi(195) => b4_nUAi(195), b6_2ZTGIf_0
         => \b6_2ZTGIf[65]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(158), mdiclink_reg_0 => mdiclink_reg(9));
    
    b8_1LbcgKeQ0 : b8_1LbcQDr1_x_133_0
      port map(b4_nUAi(104) => b4_nUAi(104), b4_nUAi(103) => 
        b4_nUAi(103), b4_nUAi(102) => b4_nUAi(102), b6_2ZTGIf_0
         => \b6_2ZTGIf[34]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(106), mdiclink_reg_0 => mdiclink_reg(61));
    
    b9_1LbcgKGAl : b8_1LbcQDr1_x_3_0
      port map(b4_nUAi(494) => b4_nUAi(494), b4_nUAi(493) => 
        b4_nUAi(493), b4_nUAi(492) => b4_nUAi(492), b6_2ZTGIf_0
         => \b6_2ZTGIf[164]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(91), mdiclink_reg_0 => mdiclink_reg(76));
    
    b9_1LbcgKGA5 : b8_1LbcQDr1_x_1_0
      port map(b4_nUAi(500) => b4_nUAi(500), b4_nUAi(499) => 
        b4_nUAi(499), b4_nUAi(498) => b4_nUAi(498), b6_2ZTGIf_0
         => \b6_2ZTGIf[166]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(89), mdiclink_reg_0 => mdiclink_reg(78));
    
    b8_1LbcgKoQ0 : b8_1LbcQDr1_x_103_0
      port map(b4_nUAi(194) => b4_nUAi(194), b4_nUAi(193) => 
        b4_nUAi(193), b4_nUAi(192) => b4_nUAi(192), b6_2ZTGIf_0
         => \b6_2ZTGIf[64]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(159), mdiclink_reg_0 => mdiclink_reg(8));
    
    b9_1LbcgKGQl0 : b8_1LbcQDr1_x_23_0
      port map(b4_nUAi(434) => b4_nUAi(434), b4_nUAi(433) => 
        b4_nUAi(433), b4_nUAi(432) => b4_nUAi(432), b6_2ZTGIf_0
         => \b6_2ZTGIf[144]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(43), mdiclink_reg_0 => mdiclink_reg(124));
    
    b9_1LbcgKGQ50 : b8_1LbcQDr1_x_21_0
      port map(b4_nUAi(440) => b4_nUAi(440), b4_nUAi(439) => 
        b4_nUAi(439), b4_nUAi(438) => b4_nUAi(438), b6_2ZTGIf_0
         => \b6_2ZTGIf[146]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(41), mdiclink_reg_0 => mdiclink_reg(126));
    
    b9_1LbcgKGUV : b8_1LbcQDr1_x_14_0
      port map(b4_nUAi(461) => b4_nUAi(461), b4_nUAi(460) => 
        b4_nUAi(460), b4_nUAi(459) => b4_nUAi(459), b6_2ZTGIf_0
         => \b6_2ZTGIf[153]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(134), mdiclink_reg_0 => mdiclink_reg(33));
    
    b8_1LbcgKwQ0 : b8_1LbcQDr1_x_143_0
      port map(b4_nUAi(74) => b4_nUAi(74), b4_nUAi(73) => 
        b4_nUAi(73), b4_nUAi(72) => b4_nUAi(72), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[24]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(164), mdiclink_reg_0 => mdiclink_reg(3));
    
    b8_1LbcgKwI : b8_1LbcQDr1_x_145_0
      port map(b4_nUAi(68) => b4_nUAi(68), b4_nUAi(67) => 
        b4_nUAi(67), b4_nUAi(66) => b4_nUAi(66), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[22]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(166), mdiclink_reg_0 => mdiclink_reg(1));
    
    b8_1LbcgKoI : b8_1LbcQDr1_x_105_0
      port map(b4_nUAi(188) => b4_nUAi(188), b4_nUAi(187) => 
        b4_nUAi(187), b4_nUAi(186) => b4_nUAi(186), b6_2ZTGIf_0
         => \b6_2ZTGIf[62]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(161), mdiclink_reg_0 => mdiclink_reg(6));
    
    b8_1LbcgKES0 : b8_1LbcQDr1_x_126_0
      port map(b4_nUAi(125) => b4_nUAi(125), b4_nUAi(124) => 
        b4_nUAi(124), b4_nUAi(123) => b4_nUAi(123), b6_2ZTGIf_0
         => \b6_2ZTGIf[41]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(21), mdiclink_reg_0 => mdiclink_reg(146));
    
    b8_1LbcgKxn : b8_1LbcQDr1_x_89_0
      port map(b4_nUAi(236) => b4_nUAi(236), b4_nUAi(235) => 
        b4_nUAi(235), b4_nUAi(234) => b4_nUAi(234), b6_2ZTGIf_0
         => \b6_2ZTGIf[78]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(145), mdiclink_reg_0 => mdiclink_reg(22));
    
    b8_1LbcgKGn : b8_1LbcQDr1_x_149_0
      port map(b4_nUAi(56) => b4_nUAi(56), b4_nUAi(55) => 
        b4_nUAi(55), b4_nUAi(54) => b4_nUAi(54), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[18]\, b11_OFWNT9L_8tZ_0 => b11_OFWNT9L_8tZ(76), 
        mdiclink_reg_0 => mdiclink_reg(91));
    
    b8_1LbcgKbJ : b8_1LbcQDr1_x_80_0
      port map(b4_nUAi(263) => b4_nUAi(263), b4_nUAi(262) => 
        b4_nUAi(262), b4_nUAi(261) => b4_nUAi(261), b6_2ZTGIf_0
         => \b6_2ZTGIf[87]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(135), mdiclink_reg_0 => mdiclink_reg(32));
    
    b8_1LbcgKER0 : b8_1LbcQDr1_x_127_0
      port map(b4_nUAi(122) => b4_nUAi(122), b4_nUAi(121) => 
        b4_nUAi(121), b4_nUAi(120) => b4_nUAi(120), b6_2ZTGIf_0
         => \b6_2ZTGIf[40]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(22), mdiclink_reg_0 => mdiclink_reg(145));
    
    b8_1LbcgKeA : b8_1LbcQDr1_x_131_0
      port map(b4_nUAi(110) => b4_nUAi(110), b4_nUAi(109) => 
        b4_nUAi(109), b4_nUAi(108) => b4_nUAi(108), b6_2ZTGIf_0
         => \b6_2ZTGIf[36]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(26), mdiclink_reg_0 => mdiclink_reg(141));
    
    b8_1LbcgKIn : b8_1LbcQDr1_x_109_0
      port map(b4_nUAi(176) => b4_nUAi(176), b4_nUAi(175) => 
        b4_nUAi(175), b4_nUAi(174) => b4_nUAi(174), b6_2ZTGIf_0
         => \b6_2ZTGIf[58]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(84), mdiclink_reg_0 => mdiclink_reg(83));
    
    b9_1LbcgKGIV : b8_1LbcQDr1_x_44_0
      port map(b4_nUAi(371) => b4_nUAi(371), b4_nUAi(370) => 
        b4_nUAi(370), b4_nUAi(369) => b4_nUAi(369), b6_2ZTGIf_0
         => \b6_2ZTGIf[123]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(30), mdiclink_reg_0 => mdiclink_reg(137));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b8_1LbcgKxV : b8_1LbcQDr1_x_88_0
      port map(b4_nUAi(239) => b4_nUAi(239), b4_nUAi(238) => 
        b4_nUAi(238), b4_nUAi(237) => b4_nUAi(237), b6_2ZTGIf_0
         => \b6_2ZTGIf[79]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(143), mdiclink_reg_0 => mdiclink_reg(24));
    
    b8_1LbcgKGV : b8_1LbcQDr1_x_148_0
      port map(b4_nUAi(59) => b4_nUAi(59), b4_nUAi(58) => 
        b4_nUAi(58), b4_nUAi(57) => b4_nUAi(57), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[19]\, b11_OFWNT9L_8tZ_0 => b11_OFWNT9L_8tZ(64), 
        mdiclink_reg_0 => mdiclink_reg(103));
    
    b9_1LbcgKGql : b8_1LbcQDr1_x_33_0
      port map(b4_nUAi(404) => b4_nUAi(404), b4_nUAi(403) => 
        b4_nUAi(403), b4_nUAi(402) => b4_nUAi(402), b6_2ZTGIf_0
         => \b6_2ZTGIf[134]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(6), mdiclink_reg_0 => mdiclink_reg(161));
    
    b8_1LbcgKIV : b8_1LbcQDr1_x_108_0
      port map(b4_nUAi(179) => b4_nUAi(179), b4_nUAi(178) => 
        b4_nUAi(178), b4_nUAi(177) => b4_nUAi(177), b6_2ZTGIf_0
         => \b6_2ZTGIf[59]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(83), mdiclink_reg_0 => mdiclink_reg(84));
    
    b7_1LbcgKE0 : b8_1LbcQDr1_x_163_0
      port map(b4_nUAi(14) => b4_nUAi(14), b4_nUAi(13) => 
        b4_nUAi(13), b4_nUAi(12) => b4_nUAi(12), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[4]\, b11_OFWNT9L_8tZ_0 => b11_OFWNT9L_8tZ(102), 
        mdiclink_reg_0 => mdiclink_reg(65));
    
    b9_1LbcgKGq5 : b8_1LbcQDr1_x_31_0
      port map(b4_nUAi(410) => b4_nUAi(410), b4_nUAi(409) => 
        b4_nUAi(409), b4_nUAi(408) => b4_nUAi(408), b6_2ZTGIf_0
         => \b6_2ZTGIf[136]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(51), mdiclink_reg_0 => mdiclink_reg(116));
    
    b8_1LbcgKwJ : b8_1LbcQDr1_x_140_0
      port map(b4_nUAi(83) => b4_nUAi(83), b4_nUAi(82) => 
        b4_nUAi(82), b4_nUAi(81) => b4_nUAi(81), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[27]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(131), mdiclink_reg_0 => mdiclink_reg(36));
    
    b8_1LbcgKoJ : b8_1LbcQDr1_x_100_0
      port map(b4_nUAi(203) => b4_nUAi(203), b4_nUAi(202) => 
        b4_nUAi(202), b4_nUAi(201) => b4_nUAi(201), b6_2ZTGIf_0
         => \b6_2ZTGIf[67]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(156), mdiclink_reg_0 => mdiclink_reg(11));
    
    b9_1LbcgKGSl : b8_1LbcQDr1_x_53_0
      port map(b4_nUAi(344) => b4_nUAi(344), b4_nUAi(343) => 
        b4_nUAi(343), b4_nUAi(342) => b4_nUAi(342), b6_2ZTGIf_0
         => \b6_2ZTGIf[114]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(110), mdiclink_reg_0 => mdiclink_reg(57));
    
    b8_1LbcgKJA : b8_1LbcQDr1_x_71_0
      port map(b4_nUAi(290) => b4_nUAi(290), b4_nUAi(289) => 
        b4_nUAi(289), b4_nUAi(288) => b4_nUAi(288), b6_2ZTGIf_0
         => \b6_2ZTGIf[96]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(4), mdiclink_reg_0 => mdiclink_reg(163));
    
    b9_1LbcgKGS5 : b8_1LbcQDr1_x_51_0
      port map(b4_nUAi(350) => b4_nUAi(350), b4_nUAi(349) => 
        b4_nUAi(349), b4_nUAi(348) => b4_nUAi(348), b6_2ZTGIf_0
         => \b6_2ZTGIf[116]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(108), mdiclink_reg_0 => mdiclink_reg(59));
    
    b9_1LbcgKGRl : b8_1LbcQDr1_x_63_0
      port map(b4_nUAi(314) => b4_nUAi(314), b4_nUAi(313) => 
        b4_nUAi(313), b4_nUAi(312) => b4_nUAi(312), b6_2ZTGIf_0
         => \b6_2ZTGIf[104]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(123), mdiclink_reg_0 => mdiclink_reg(44));
    
    b8_1LbcgKeq : b8_1LbcQDr1_x_134_0
      port map(b4_nUAi(101) => b4_nUAi(101), b4_nUAi(100) => 
        b4_nUAi(100), b4_nUAi(99) => b4_nUAi(99), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[33]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(116), mdiclink_reg_0 => mdiclink_reg(51));
    
    b9_1LbcgKGR5 : b8_1LbcQDr1_x_61_0
      port map(b4_nUAi(320) => b4_nUAi(320), b4_nUAi(319) => 
        b4_nUAi(319), b4_nUAi(318) => b4_nUAi(318), b6_2ZTGIf_0
         => \b6_2ZTGIf[106]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(121), mdiclink_reg_0 => mdiclink_reg(46));
    
    b8_1LbcgKEn0 : b8_1LbcQDr1_x_119_0
      port map(b4_nUAi(146) => b4_nUAi(146), b4_nUAi(145) => 
        b4_nUAi(145), b4_nUAi(144) => b4_nUAi(144), b6_2ZTGIf_0
         => \b6_2ZTGIf[48]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(70), mdiclink_reg_0 => mdiclink_reg(97));
    
    b8_1LbcgKxU : b8_1LbcQDr1_x_92_0
      port map(b4_nUAi(227) => b4_nUAi(227), b4_nUAi(226) => 
        b4_nUAi(226), b4_nUAi(225) => b4_nUAi(225), b6_2ZTGIf_0
         => \b6_2ZTGIf[75]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(148), mdiclink_reg_0 => mdiclink_reg(19));
    
    b8_1LbcgKGU : b8_1LbcQDr1_x_152_0
      port map(b4_nUAi(47) => b4_nUAi(47), b4_nUAi(46) => 
        b4_nUAi(46), b4_nUAi(45) => b4_nUAi(45), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[15]\, b11_OFWNT9L_8tZ_0 => b11_OFWNT9L_8tZ(79), 
        mdiclink_reg_0 => mdiclink_reg(88));
    
    b7_1LbcgKx : b8_1LbcQDr1_x_160_0
      port map(b4_nUAi(23) => b4_nUAi(23), b4_nUAi(22) => 
        b4_nUAi(22), b4_nUAi(21) => b4_nUAi(21), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[7]\, b11_OFWNT9L_8tZ_0 => b11_OFWNT9L_8tZ(99), 
        mdiclink_reg_0 => mdiclink_reg(68));
    
    b8_1LbcgKIU : b8_1LbcQDr1_x_112_0
      port map(b4_nUAi(167) => b4_nUAi(167), b4_nUAi(166) => 
        b4_nUAi(166), b4_nUAi(165) => b4_nUAi(165), b6_2ZTGIf_0
         => \b6_2ZTGIf[55]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(87), mdiclink_reg_0 => mdiclink_reg(80));
    
    b8_1LbcgKEV0 : b8_1LbcQDr1_x_118_0
      port map(b4_nUAi(149) => b4_nUAi(149), b4_nUAi(148) => 
        b4_nUAi(148), b4_nUAi(147) => b4_nUAi(147), b6_2ZTGIf_0
         => \b6_2ZTGIf[49]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(69), mdiclink_reg_0 => mdiclink_reg(98));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b8_1LbcgKeS : b8_1LbcQDr1_x_136_0
      port map(b4_nUAi(95) => b4_nUAi(95), b4_nUAi(94) => 
        b4_nUAi(94), b4_nUAi(93) => b4_nUAi(93), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[31]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(118), mdiclink_reg_0 => mdiclink_reg(49));
    
    b8_1LbcgKxI : b8_1LbcQDr1_x_95_0
      port map(b4_nUAi(218) => b4_nUAi(218), b4_nUAi(217) => 
        b4_nUAi(217), b4_nUAi(216) => b4_nUAi(216), b6_2ZTGIf_0
         => \b6_2ZTGIf[72]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(151), mdiclink_reg_0 => mdiclink_reg(16));
    
    b8_1LbcgKGI : b8_1LbcQDr1_x_155_0
      port map(b4_nUAi(38) => b4_nUAi(38), b4_nUAi(37) => 
        b4_nUAi(37), b4_nUAi(36) => b4_nUAi(36), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[12]\, b11_OFWNT9L_8tZ_0 => b11_OFWNT9L_8tZ(94), 
        mdiclink_reg_0 => mdiclink_reg(73));
    
    b8_1LbcgKeR : b8_1LbcQDr1_x_137_0
      port map(b4_nUAi(92) => b4_nUAi(92), b4_nUAi(91) => 
        b4_nUAi(91), b4_nUAi(90) => b4_nUAi(90), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[30]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(128), mdiclink_reg_0 => mdiclink_reg(39));
    
    b9_1LbcgKGAd : b8_1LbcQDr1_x_5_0
      port map(b4_nUAi(488) => b4_nUAi(488), b4_nUAi(487) => 
        b4_nUAi(487), b4_nUAi(486) => b4_nUAi(486), b6_2ZTGIf_0
         => \b6_2ZTGIf[162]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(53), mdiclink_reg_0 => mdiclink_reg(114));
    
    b8_1LbcgKII : b8_1LbcQDr1_x_115_0
      port map(b4_nUAi(158) => b4_nUAi(158), b4_nUAi(157) => 
        b4_nUAi(157), b4_nUAi(156) => b4_nUAi(156), b6_2ZTGIf_0
         => \b6_2ZTGIf[52]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(66), mdiclink_reg_0 => mdiclink_reg(101));
    
    b9_1LbcgKGQd0 : b8_1LbcQDr1_x_25_0
      port map(b4_nUAi(428) => b4_nUAi(428), b4_nUAi(427) => 
        b4_nUAi(427), b4_nUAi(426) => b4_nUAi(426), b6_2ZTGIf_0
         => \b6_2ZTGIf[142]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(45), mdiclink_reg_0 => mdiclink_reg(122));
    
    b8_1LbcgKJq : b8_1LbcQDr1_x_74_0
      port map(b4_nUAi(281) => b4_nUAi(281), b4_nUAi(280) => 
        b4_nUAi(280), b4_nUAi(279) => b4_nUAi(279), b6_2ZTGIf_0
         => \b6_2ZTGIf[93]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(40), mdiclink_reg_0 => mdiclink_reg(127));
    
    b7_1LbcgKo : b8_1LbcQDr1_x_161_0
      port map(b4_nUAi(20) => b4_nUAi(20), b4_nUAi(19) => 
        b4_nUAi(19), b4_nUAi(18) => b4_nUAi(18), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[6]\, b11_OFWNT9L_8tZ_0 => b11_OFWNT9L_8tZ(100), 
        mdiclink_reg_0 => mdiclink_reg(67));
    
    b9_1LbcgKGAp : b8_1LbcQDr1_x_2_0
      port map(b4_nUAi(497) => b4_nUAi(497), b4_nUAi(496) => 
        b4_nUAi(496), b4_nUAi(495) => b4_nUAi(495), b6_2ZTGIf_0
         => \b6_2ZTGIf[165]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(90), mdiclink_reg_0 => mdiclink_reg(77));
    
    b9_1LbcgKGQp0 : b8_1LbcQDr1_x_22_0
      port map(b4_nUAi(437) => b4_nUAi(437), b4_nUAi(436) => 
        b4_nUAi(436), b4_nUAi(435) => b4_nUAi(435), b6_2ZTGIf_0
         => \b6_2ZTGIf[145]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(42), mdiclink_reg_0 => mdiclink_reg(125));
    
    b8_1LbcgKEU0 : b8_1LbcQDr1_x_122_0
      port map(b4_nUAi(137) => b4_nUAi(137), b4_nUAi(136) => 
        b4_nUAi(136), b4_nUAi(135) => b4_nUAi(135), b6_2ZTGIf_0
         => \b6_2ZTGIf[45]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(73), mdiclink_reg_0 => mdiclink_reg(94));
    
    b9_1LbcgKGQq0 : b8_1LbcQDr1_x_18_0
      port map(b4_nUAi(449) => b4_nUAi(449), b4_nUAi(448) => 
        b4_nUAi(448), b4_nUAi(447) => b4_nUAi(447), b6_2ZTGIf_0
         => \b6_2ZTGIf[149]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(10), mdiclink_reg_0 => mdiclink_reg(157));
    
    b9_1LbcgKGAe : b8_1LbcQDr1_x_0_0
      port map(b4_nUAi(502) => b4_nUAi(502), b4_nUAi(501) => 
        b4_nUAi(501), b6_2ZTGIf_0 => \b6_2ZTGIf[167]\, 
        b11_OFWNT9L_8tZ_0 => b11_OFWNT9L_8tZ(11), mdiclink_reg_0
         => mdiclink_reg(156), b12_PSyi_XlK_qHv => 
        b12_PSyi_XlK_qHv);
    
    b8_1LbcgKJS : b8_1LbcQDr1_x_76_0
      port map(b4_nUAi(275) => b4_nUAi(275), b4_nUAi(274) => 
        b4_nUAi(274), b4_nUAi(273) => b4_nUAi(273), b6_2ZTGIf_0
         => \b6_2ZTGIf[91]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(93), mdiclink_reg_0 => mdiclink_reg(74));
    
    b7_1LbcgKI : b8_1LbcQDr1_x_162_0
      port map(b4_nUAi(17) => b4_nUAi(17), b4_nUAi(16) => 
        b4_nUAi(16), b4_nUAi(15) => b4_nUAi(15), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[5]\, b11_OFWNT9L_8tZ_0 => b11_OFWNT9L_8tZ(101), 
        mdiclink_reg_0 => mdiclink_reg(66));
    
    b9_1LbcgKGQS0 : b8_1LbcQDr1_x_19_0
      port map(b4_nUAi(446) => b4_nUAi(446), b4_nUAi(445) => 
        b4_nUAi(445), b4_nUAi(444) => b4_nUAi(444), b6_2ZTGIf_0
         => \b6_2ZTGIf[148]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(37), mdiclink_reg_0 => mdiclink_reg(130));
    
    b8_1LbcgKJR : b8_1LbcQDr1_x_77_0
      port map(b4_nUAi(272) => b4_nUAi(272), b4_nUAi(271) => 
        b4_nUAi(271), b4_nUAi(270) => b4_nUAi(270), b6_2ZTGIf_0
         => \b6_2ZTGIf[90]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(107), mdiclink_reg_0 => mdiclink_reg(60));
    
    b9_1LbcgKGAm : b8_1LbcQDr1_x_7_0
      port map(b4_nUAi(482) => b4_nUAi(482), b4_nUAi(481) => 
        b4_nUAi(481), b4_nUAi(480) => b4_nUAi(480), b6_2ZTGIf_0
         => \b6_2ZTGIf[160]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(55), mdiclink_reg_0 => mdiclink_reg(112));
    
    b9_1LbcgKGqd : b8_1LbcQDr1_x_35_0
      port map(b4_nUAi(398) => b4_nUAi(398), b4_nUAi(397) => 
        b4_nUAi(397), b4_nUAi(396) => b4_nUAi(396), b6_2ZTGIf_0
         => \b6_2ZTGIf[132]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(13), mdiclink_reg_0 => mdiclink_reg(154));
    
    b9_1LbcgKGQe0 : b8_1LbcQDr1_x_20_0
      port map(b4_nUAi(443) => b4_nUAi(443), b4_nUAi(442) => 
        b4_nUAi(442), b4_nUAi(441) => b4_nUAi(441), b6_2ZTGIf_0
         => \b6_2ZTGIf[147]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(39), mdiclink_reg_0 => mdiclink_reg(128));
    
    b8_1LbcgKxJ : b8_1LbcQDr1_x_90_0
      port map(b4_nUAi(233) => b4_nUAi(233), b4_nUAi(232) => 
        b4_nUAi(232), b4_nUAi(231) => b4_nUAi(231), b6_2ZTGIf_0
         => \b6_2ZTGIf[77]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(146), mdiclink_reg_0 => mdiclink_reg(21));
    
    b8_1LbcgKGJ : b8_1LbcQDr1_x_150_0
      port map(b4_nUAi(53) => b4_nUAi(53), b4_nUAi(52) => 
        b4_nUAi(52), b4_nUAi(51) => b4_nUAi(51), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[17]\, b11_OFWNT9L_8tZ_0 => b11_OFWNT9L_8tZ(77), 
        mdiclink_reg_0 => mdiclink_reg(90));
    
    b8_1LbcgKIQ0 : b8_1LbcQDr1_x_113_0
      port map(b4_nUAi(164) => b4_nUAi(164), b4_nUAi(163) => 
        b4_nUAi(163), b4_nUAi(162) => b4_nUAi(162), b6_2ZTGIf_0
         => \b6_2ZTGIf[54]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(88), mdiclink_reg_0 => mdiclink_reg(79));
    
    b7_1LbcgKw : b8_1LbcQDr1_x_165_0
      port map(b4_nUAi(8) => b4_nUAi(8), b4_nUAi(7) => b4_nUAi(7), 
        b4_nUAi(6) => b4_nUAi(6), b6_2ZTGIf_0 => \b6_2ZTGIf[2]\, 
        b11_OFWNT9L_8tZ_0 => b11_OFWNT9L_8tZ(104), mdiclink_reg_0
         => mdiclink_reg(63));
    
    b8_1LbcgKIJ : b8_1LbcQDr1_x_110_0
      port map(b4_nUAi(173) => b4_nUAi(173), b4_nUAi(172) => 
        b4_nUAi(172), b4_nUAi(171) => b4_nUAi(171), b6_2ZTGIf_0
         => \b6_2ZTGIf[57]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(85), mdiclink_reg_0 => mdiclink_reg(82));
    
    b9_1LbcgKGQm0 : b8_1LbcQDr1_x_27_0
      port map(b4_nUAi(422) => b4_nUAi(422), b4_nUAi(421) => 
        b4_nUAi(421), b4_nUAi(420) => b4_nUAi(420), b6_2ZTGIf_0
         => \b6_2ZTGIf[140]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(47), mdiclink_reg_0 => mdiclink_reg(120));
    
    b8_1LbcgKen : b8_1LbcQDr1_x_129_0
      port map(b4_nUAi(116) => b4_nUAi(116), b4_nUAi(115) => 
        b4_nUAi(115), b4_nUAi(114) => b4_nUAi(114), b6_2ZTGIf_0
         => \b6_2ZTGIf[38]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(24), mdiclink_reg_0 => mdiclink_reg(143));
    
    b8_1LbcgKbA : b8_1LbcQDr1_x_81_0
      port map(b4_nUAi(260) => b4_nUAi(260), b4_nUAi(259) => 
        b4_nUAi(259), b4_nUAi(258) => b4_nUAi(258), b6_2ZTGIf_0
         => \b6_2ZTGIf[86]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(136), mdiclink_reg_0 => mdiclink_reg(31));
    
    b8_1LbcgKEI0 : b8_1LbcQDr1_x_125_0
      port map(b4_nUAi(128) => b4_nUAi(128), b4_nUAi(127) => 
        b4_nUAi(127), b4_nUAi(126) => b4_nUAi(126), b6_2ZTGIf_0
         => \b6_2ZTGIf[42]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(20), mdiclink_reg_0 => mdiclink_reg(147));
    
    b9_1LbcgKGAn : b8_1LbcQDr1_x_6_0
      port map(b4_nUAi(485) => b4_nUAi(485), b4_nUAi(484) => 
        b4_nUAi(484), b4_nUAi(483) => b4_nUAi(483), b6_2ZTGIf_0
         => \b6_2ZTGIf[161]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(54), mdiclink_reg_0 => mdiclink_reg(113));
    
    b9_1LbcgKGqp : b8_1LbcQDr1_x_32_0
      port map(b4_nUAi(407) => b4_nUAi(407), b4_nUAi(406) => 
        b4_nUAi(406), b4_nUAi(405) => b4_nUAi(405), b6_2ZTGIf_0
         => \b6_2ZTGIf[135]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(127), mdiclink_reg_0 => mdiclink_reg(40));
    
    b8_1LbcgKeV : b8_1LbcQDr1_x_128_0
      port map(b4_nUAi(119) => b4_nUAi(119), b4_nUAi(118) => 
        b4_nUAi(118), b4_nUAi(117) => b4_nUAi(117), b6_2ZTGIf_0
         => \b6_2ZTGIf[39]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(23), mdiclink_reg_0 => mdiclink_reg(144));
    
    b9_1LbcgKGQn0 : b8_1LbcQDr1_x_26_0
      port map(b4_nUAi(425) => b4_nUAi(425), b4_nUAi(424) => 
        b4_nUAi(424), b4_nUAi(423) => b4_nUAi(423), b6_2ZTGIf_0
         => \b6_2ZTGIf[141]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(46), mdiclink_reg_0 => mdiclink_reg(121));
    
    b9_1LbcgKGqq : b8_1LbcQDr1_x_28_0
      port map(b4_nUAi(419) => b4_nUAi(419), b4_nUAi(418) => 
        b4_nUAi(418), b4_nUAi(417) => b4_nUAi(417), b6_2ZTGIf_0
         => \b6_2ZTGIf[139]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(48), mdiclink_reg_0 => mdiclink_reg(119));
    
    b9_1LbcgKGSd : b8_1LbcQDr1_x_55_0
      port map(b4_nUAi(338) => b4_nUAi(338), b4_nUAi(337) => 
        b4_nUAi(337), b4_nUAi(336) => b4_nUAi(336), b6_2ZTGIf_0
         => \b6_2ZTGIf[112]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(112), mdiclink_reg_0 => mdiclink_reg(55));
    
    b9_1LbcgKGUl : b8_1LbcQDr1_x_13_0
      port map(b4_nUAi(464) => b4_nUAi(464), b4_nUAi(463) => 
        b4_nUAi(463), b4_nUAi(462) => b4_nUAi(462), b6_2ZTGIf_0
         => \b6_2ZTGIf[154]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(62), mdiclink_reg_0 => mdiclink_reg(105));
    
    b9_1LbcgKGRd : b8_1LbcQDr1_x_65_0
      port map(b4_nUAi(308) => b4_nUAi(308), b4_nUAi(307) => 
        b4_nUAi(307), b4_nUAi(306) => b4_nUAi(306), b6_2ZTGIf_0
         => \b6_2ZTGIf[102]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(125), mdiclink_reg_0 => mdiclink_reg(42));
    
    b9_1LbcgKGqS : b8_1LbcQDr1_x_29_0
      port map(b4_nUAi(416) => b4_nUAi(416), b4_nUAi(415) => 
        b4_nUAi(415), b4_nUAi(414) => b4_nUAi(414), b6_2ZTGIf_0
         => \b6_2ZTGIf[138]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(49), mdiclink_reg_0 => mdiclink_reg(118));
    
    b9_1LbcgKGU5 : b8_1LbcQDr1_x_11_0
      port map(b4_nUAi(470) => b4_nUAi(470), b4_nUAi(469) => 
        b4_nUAi(469), b4_nUAi(468) => b4_nUAi(468), b6_2ZTGIf_0
         => \b6_2ZTGIf[156]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(59), mdiclink_reg_0 => mdiclink_reg(108));
    
    b9_1LbcgKGqe : b8_1LbcQDr1_x_30_0
      port map(b4_nUAi(413) => b4_nUAi(413), b4_nUAi(412) => 
        b4_nUAi(412), b4_nUAi(411) => b4_nUAi(411), b6_2ZTGIf_0
         => \b6_2ZTGIf[137]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(50), mdiclink_reg_0 => mdiclink_reg(117));
    
    b8_1LbcgKwA : b8_1LbcQDr1_x_141_0
      port map(b4_nUAi(80) => b4_nUAi(80), b4_nUAi(79) => 
        b4_nUAi(79), b4_nUAi(78) => b4_nUAi(78), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[26]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(162), mdiclink_reg_0 => mdiclink_reg(5));
    
    b7_1LbcgKF : b8_1LbcQDr1_x_167_0
      port map(b4_nUAi(2) => b4_nUAi(2), b4_nUAi(1) => b4_nUAi(1), 
        b4_nUAi(0) => b4_nUAi(0), b6_2ZTGIf_0 => \b6_2ZTGIf[0]\, 
        b11_OFWNT9L_8tZ_0 => b11_OFWNT9L_8tZ(133), mdiclink_reg_0
         => mdiclink_reg(34));
    
    b9_1LbcgKGqm : b8_1LbcQDr1_x_37_0
      port map(b4_nUAi(392) => b4_nUAi(392), b4_nUAi(391) => 
        b4_nUAi(391), b4_nUAi(390) => b4_nUAi(390), b6_2ZTGIf_0
         => \b6_2ZTGIf[130]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(15), mdiclink_reg_0 => mdiclink_reg(152));
    
    b8_1LbcgKoA : b8_1LbcQDr1_x_101_0
      port map(b4_nUAi(200) => b4_nUAi(200), b4_nUAi(199) => 
        b4_nUAi(199), b4_nUAi(198) => b4_nUAi(198), b6_2ZTGIf_0
         => \b6_2ZTGIf[66]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(157), mdiclink_reg_0 => mdiclink_reg(10));
    
    b9_1LbcgKGSp : b8_1LbcQDr1_x_52_0
      port map(b4_nUAi(347) => b4_nUAi(347), b4_nUAi(346) => 
        b4_nUAi(346), b4_nUAi(345) => b4_nUAi(345), b6_2ZTGIf_0
         => \b6_2ZTGIf[115]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(109), mdiclink_reg_0 => mdiclink_reg(58));
    
    b9_1LbcgKGRp : b8_1LbcQDr1_x_62_0
      port map(b4_nUAi(317) => b4_nUAi(317), b4_nUAi(316) => 
        b4_nUAi(316), b4_nUAi(315) => b4_nUAi(315), b6_2ZTGIf_0
         => \b6_2ZTGIf[105]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(122), mdiclink_reg_0 => mdiclink_reg(45));
    
    b8_1LbcgKJn : b8_1LbcQDr1_x_69_0
      port map(b4_nUAi(296) => b4_nUAi(296), b4_nUAi(295) => 
        b4_nUAi(295), b4_nUAi(294) => b4_nUAi(294), b6_2ZTGIf_0
         => \b6_2ZTGIf[98]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(2), mdiclink_reg_0 => mdiclink_reg(165));
    
    b8_1LbcgKbq : b8_1LbcQDr1_x_84_0
      port map(b4_nUAi(251) => b4_nUAi(251), b4_nUAi(250) => 
        b4_nUAi(250), b4_nUAi(249) => b4_nUAi(249), b6_2ZTGIf_0
         => \b6_2ZTGIf[83]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(139), mdiclink_reg_0 => mdiclink_reg(28));
    
    b9_1LbcgKGIl : b8_1LbcQDr1_x_43_0
      port map(b4_nUAi(374) => b4_nUAi(374), b4_nUAi(373) => 
        b4_nUAi(373), b4_nUAi(372) => b4_nUAi(372), b6_2ZTGIf_0
         => \b6_2ZTGIf[124]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(29), mdiclink_reg_0 => mdiclink_reg(138));
    
    b8_1LbcgKEJ0 : b8_1LbcQDr1_x_120_0
      port map(b4_nUAi(143) => b4_nUAi(143), b4_nUAi(142) => 
        b4_nUAi(142), b4_nUAi(141) => b4_nUAi(141), b6_2ZTGIf_0
         => \b6_2ZTGIf[47]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(71), mdiclink_reg_0 => mdiclink_reg(96));
    
    b9_1LbcgKGSq : b8_1LbcQDr1_x_48_0
      port map(b4_nUAi(359) => b4_nUAi(359), b4_nUAi(358) => 
        b4_nUAi(358), b4_nUAi(357) => b4_nUAi(357), b6_2ZTGIf_0
         => \b6_2ZTGIf[119]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(34), mdiclink_reg_0 => mdiclink_reg(133));
    
    b9_1LbcgKGI5 : b8_1LbcQDr1_x_41_0
      port map(b4_nUAi(380) => b4_nUAi(380), b4_nUAi(379) => 
        b4_nUAi(379), b4_nUAi(378) => b4_nUAi(378), b6_2ZTGIf_0
         => \b6_2ZTGIf[126]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(19), mdiclink_reg_0 => mdiclink_reg(148));
    
    b9_1LbcgKGqn : b8_1LbcQDr1_x_36_0
      port map(b4_nUAi(395) => b4_nUAi(395), b4_nUAi(394) => 
        b4_nUAi(394), b4_nUAi(393) => b4_nUAi(393), b6_2ZTGIf_0
         => \b6_2ZTGIf[131]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(14), mdiclink_reg_0 => mdiclink_reg(153));
    
    b9_1LbcgKGRq : b8_1LbcQDr1_x_58_0
      port map(b4_nUAi(329) => b4_nUAi(329), b4_nUAi(328) => 
        b4_nUAi(328), b4_nUAi(327) => b4_nUAi(327), b6_2ZTGIf_0
         => \b6_2ZTGIf[109]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(115), mdiclink_reg_0 => mdiclink_reg(52));
    
    b9_1LbcgKGAV : b8_1LbcQDr1_x_4_0
      port map(b4_nUAi(491) => b4_nUAi(491), b4_nUAi(490) => 
        b4_nUAi(490), b4_nUAi(489) => b4_nUAi(489), b6_2ZTGIf_0
         => \b6_2ZTGIf[163]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(52), mdiclink_reg_0 => mdiclink_reg(115));
    
    b9_1LbcgKGSS : b8_1LbcQDr1_x_49_0
      port map(b4_nUAi(356) => b4_nUAi(356), b4_nUAi(355) => 
        b4_nUAi(355), b4_nUAi(354) => b4_nUAi(354), b6_2ZTGIf_0
         => \b6_2ZTGIf[118]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(35), mdiclink_reg_0 => mdiclink_reg(132));
    
    b8_1LbcgKJV : b8_1LbcQDr1_x_68_0
      port map(b4_nUAi(299) => b4_nUAi(299), b4_nUAi(298) => 
        b4_nUAi(298), b4_nUAi(297) => b4_nUAi(297), b6_2ZTGIf_0
         => \b6_2ZTGIf[99]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(1), mdiclink_reg_0 => mdiclink_reg(166));
    
    b8_1LbcgKeU : b8_1LbcQDr1_x_132_0
      port map(b4_nUAi(107) => b4_nUAi(107), b4_nUAi(106) => 
        b4_nUAi(106), b4_nUAi(105) => b4_nUAi(105), b6_2ZTGIf_0
         => \b6_2ZTGIf[35]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(27), mdiclink_reg_0 => mdiclink_reg(140));
    
    b9_1LbcgKGRS : b8_1LbcQDr1_x_59_0
      port map(b4_nUAi(326) => b4_nUAi(326), b4_nUAi(325) => 
        b4_nUAi(325), b4_nUAi(324) => b4_nUAi(324), b6_2ZTGIf_0
         => \b6_2ZTGIf[108]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(119), mdiclink_reg_0 => mdiclink_reg(48));
    
    b7_1LbcgKe : b8_1LbcQDr1_x_164_0
      port map(b4_nUAi(11) => b4_nUAi(11), b4_nUAi(10) => 
        b4_nUAi(10), b4_nUAi(9) => b4_nUAi(9), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[3]\, b11_OFWNT9L_8tZ_0 => b11_OFWNT9L_8tZ(103), 
        mdiclink_reg_0 => mdiclink_reg(64));
    
    b9_1LbcgKGSe : b8_1LbcQDr1_x_50_0
      port map(b4_nUAi(353) => b4_nUAi(353), b4_nUAi(352) => 
        b4_nUAi(352), b4_nUAi(351) => b4_nUAi(351), b6_2ZTGIf_0
         => \b6_2ZTGIf[117]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(36), mdiclink_reg_0 => mdiclink_reg(131));
    
    b9_1LbcgKGQV0 : b8_1LbcQDr1_x_24_0
      port map(b4_nUAi(431) => b4_nUAi(431), b4_nUAi(430) => 
        b4_nUAi(430), b4_nUAi(429) => b4_nUAi(429), b6_2ZTGIf_0
         => \b6_2ZTGIf[143]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(44), mdiclink_reg_0 => mdiclink_reg(123));
    
    b9_1LbcgKGRe : b8_1LbcQDr1_x_60_0
      port map(b4_nUAi(323) => b4_nUAi(323), b4_nUAi(322) => 
        b4_nUAi(322), b4_nUAi(321) => b4_nUAi(321), b6_2ZTGIf_0
         => \b6_2ZTGIf[107]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(120), mdiclink_reg_0 => mdiclink_reg(47));
    
    b9_1LbcgKGSm : b8_1LbcQDr1_x_57_0
      port map(b4_nUAi(332) => b4_nUAi(332), b4_nUAi(331) => 
        b4_nUAi(331), b4_nUAi(330) => b4_nUAi(330), b6_2ZTGIf_0
         => \b6_2ZTGIf[110]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(114), mdiclink_reg_0 => mdiclink_reg(53));
    
    b9_1LbcgKGRm : b8_1LbcQDr1_x_67_0
      port map(b4_nUAi(302) => b4_nUAi(302), b4_nUAi(301) => 
        b4_nUAi(301), b4_nUAi(300) => b4_nUAi(300), b6_2ZTGIf_0
         => \b6_2ZTGIf[100]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(0), mdiclink_reg_0 => mdiclink_reg(167));
    
    b8_1LbcgKbS : b8_1LbcQDr1_x_86_0
      port map(b4_nUAi(245) => b4_nUAi(245), b4_nUAi(244) => 
        b4_nUAi(244), b4_nUAi(243) => b4_nUAi(243), b6_2ZTGIf_0
         => \b6_2ZTGIf[81]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(141), mdiclink_reg_0 => mdiclink_reg(26));
    
    b8_1LbcgKbR : b8_1LbcQDr1_x_87_0
      port map(b4_nUAi(242) => b4_nUAi(242), b4_nUAi(241) => 
        b4_nUAi(241), b4_nUAi(240) => b4_nUAi(240), b6_2ZTGIf_0
         => \b6_2ZTGIf[80]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(142), mdiclink_reg_0 => mdiclink_reg(25));
    
    b8_1LbcgKeI : b8_1LbcQDr1_x_135_0
      port map(b4_nUAi(98) => b4_nUAi(98), b4_nUAi(97) => 
        b4_nUAi(97), b4_nUAi(96) => b4_nUAi(96), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[32]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(117), mdiclink_reg_0 => mdiclink_reg(50));
    
    b9_1LbcgKGSn : b8_1LbcQDr1_x_56_0
      port map(b4_nUAi(335) => b4_nUAi(335), b4_nUAi(334) => 
        b4_nUAi(334), b4_nUAi(333) => b4_nUAi(333), b6_2ZTGIf_0
         => \b6_2ZTGIf[111]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(113), mdiclink_reg_0 => mdiclink_reg(54));
    
    b8_1LbcgKwq : b8_1LbcQDr1_x_144_0
      port map(b4_nUAi(71) => b4_nUAi(71), b4_nUAi(70) => 
        b4_nUAi(70), b4_nUAi(69) => b4_nUAi(69), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[23]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(165), mdiclink_reg_0 => mdiclink_reg(2));
    
    b8_1LbcgKoq : b8_1LbcQDr1_x_104_0
      port map(b4_nUAi(191) => b4_nUAi(191), b4_nUAi(190) => 
        b4_nUAi(190), b4_nUAi(189) => b4_nUAi(189), b6_2ZTGIf_0
         => \b6_2ZTGIf[63]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(160), mdiclink_reg_0 => mdiclink_reg(7));
    
    b9_1LbcgKGRn : b8_1LbcQDr1_x_66_0
      port map(b4_nUAi(305) => b4_nUAi(305), b4_nUAi(304) => 
        b4_nUAi(304), b4_nUAi(303) => b4_nUAi(303), b6_2ZTGIf_0
         => \b6_2ZTGIf[101]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(126), mdiclink_reg_0 => mdiclink_reg(41));
    
    b9_1LbcgKGqV : b8_1LbcQDr1_x_34_0
      port map(b4_nUAi(401) => b4_nUAi(401), b4_nUAi(400) => 
        b4_nUAi(400), b4_nUAi(399) => b4_nUAi(399), b6_2ZTGIf_0
         => \b6_2ZTGIf[133]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(12), mdiclink_reg_0 => mdiclink_reg(155));
    
    b8_1LbcgKJU : b8_1LbcQDr1_x_72_0
      port map(b4_nUAi(287) => b4_nUAi(287), b4_nUAi(286) => 
        b4_nUAi(286), b4_nUAi(285) => b4_nUAi(285), b6_2ZTGIf_0
         => \b6_2ZTGIf[95]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(5), mdiclink_reg_0 => mdiclink_reg(162));
    
    b7_1LbcgKb : b8_1LbcQDr1_x_159_0
      port map(b4_nUAi(26) => b4_nUAi(26), b4_nUAi(25) => 
        b4_nUAi(25), b4_nUAi(24) => b4_nUAi(24), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[8]\, b11_OFWNT9L_8tZ_0 => b11_OFWNT9L_8tZ(98), 
        mdiclink_reg_0 => mdiclink_reg(69));
    
    b8_1LbcgKwS : b8_1LbcQDr1_x_146_0
      port map(b4_nUAi(65) => b4_nUAi(65), b4_nUAi(64) => 
        b4_nUAi(64), b4_nUAi(63) => b4_nUAi(63), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[21]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(167), mdiclink_reg_0 => mdiclink_reg(0));
    
    b8_1LbcgKoS : b8_1LbcQDr1_x_106_0
      port map(b4_nUAi(185) => b4_nUAi(185), b4_nUAi(184) => 
        b4_nUAi(184), b4_nUAi(183) => b4_nUAi(183), b6_2ZTGIf_0
         => \b6_2ZTGIf[61]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(81), mdiclink_reg_0 => mdiclink_reg(86));
    
    b8_1LbcgKwR : b8_1LbcQDr1_x_147_0
      port map(b4_nUAi(62) => b4_nUAi(62), b4_nUAi(61) => 
        b4_nUAi(61), b4_nUAi(60) => b4_nUAi(60), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[20]\, b11_OFWNT9L_8tZ_0 => b11_OFWNT9L_8tZ(63), 
        mdiclink_reg_0 => mdiclink_reg(104));
    
    b8_1LbcgKoR : b8_1LbcQDr1_x_107_0
      port map(b4_nUAi(182) => b4_nUAi(182), b4_nUAi(181) => 
        b4_nUAi(181), b4_nUAi(180) => b4_nUAi(180), b6_2ZTGIf_0
         => \b6_2ZTGIf[60]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(82), mdiclink_reg_0 => mdiclink_reg(85));
    
    b8_1LbcgKJI : b8_1LbcQDr1_x_75_0
      port map(b4_nUAi(278) => b4_nUAi(278), b4_nUAi(277) => 
        b4_nUAi(277), b4_nUAi(276) => b4_nUAi(276), b6_2ZTGIf_0
         => \b6_2ZTGIf[92]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(61), mdiclink_reg_0 => mdiclink_reg(106));
    
    b8_1LbcgKxA : b8_1LbcQDr1_x_91_0
      port map(b4_nUAi(230) => b4_nUAi(230), b4_nUAi(229) => 
        b4_nUAi(229), b4_nUAi(228) => b4_nUAi(228), b6_2ZTGIf_0
         => \b6_2ZTGIf[76]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(147), mdiclink_reg_0 => mdiclink_reg(20));
    
    b8_1LbcgKGA : b8_1LbcQDr1_x_151_0
      port map(b4_nUAi(50) => b4_nUAi(50), b4_nUAi(49) => 
        b4_nUAi(49), b4_nUAi(48) => b4_nUAi(48), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[16]\, b11_OFWNT9L_8tZ_0 => b11_OFWNT9L_8tZ(78), 
        mdiclink_reg_0 => mdiclink_reg(89));
    
    \b8_1LbcgKEQ0\ : b8_1LbcQDr1_x_123_0
      port map(b4_nUAi(134) => b4_nUAi(134), b4_nUAi(133) => 
        b4_nUAi(133), b4_nUAi(132) => b4_nUAi(132), b6_2ZTGIf_0
         => \b6_2ZTGIf[44]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(74), mdiclink_reg_0 => mdiclink_reg(93));
    
    b8_1LbcgKeJ : b8_1LbcQDr1_x_130_0
      port map(b4_nUAi(113) => b4_nUAi(113), b4_nUAi(112) => 
        b4_nUAi(112), b4_nUAi(111) => b4_nUAi(111), b6_2ZTGIf_0
         => \b6_2ZTGIf[37]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(25), mdiclink_reg_0 => mdiclink_reg(142));
    
    b9_1LbcgKGSV : b8_1LbcQDr1_x_54_0
      port map(b4_nUAi(341) => b4_nUAi(341), b4_nUAi(340) => 
        b4_nUAi(340), b4_nUAi(339) => b4_nUAi(339), b6_2ZTGIf_0
         => \b6_2ZTGIf[113]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(111), mdiclink_reg_0 => mdiclink_reg(56));
    
    b8_1LbcgKbn : b8_1LbcQDr1_x_79_0
      port map(b4_nUAi(266) => b4_nUAi(266), b4_nUAi(265) => 
        b4_nUAi(265), b4_nUAi(264) => b4_nUAi(264), b6_2ZTGIf_0
         => \b6_2ZTGIf[88]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(144), mdiclink_reg_0 => mdiclink_reg(23));
    
    b9_1LbcgKGRV : b8_1LbcQDr1_x_64_0
      port map(b4_nUAi(311) => b4_nUAi(311), b4_nUAi(310) => 
        b4_nUAi(310), b4_nUAi(309) => b4_nUAi(309), b6_2ZTGIf_0
         => \b6_2ZTGIf[103]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(124), mdiclink_reg_0 => mdiclink_reg(43));
    
    b8_1LbcgKIA : b8_1LbcQDr1_x_111_0
      port map(b4_nUAi(170) => b4_nUAi(170), b4_nUAi(169) => 
        b4_nUAi(169), b4_nUAi(168) => b4_nUAi(168), b6_2ZTGIf_0
         => \b6_2ZTGIf[56]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(86), mdiclink_reg_0 => mdiclink_reg(81));
    
    b8_1LbcgKbQ0 : b8_1LbcQDr1_x_83_0
      port map(b4_nUAi(254) => b4_nUAi(254), b4_nUAi(253) => 
        b4_nUAi(253), b4_nUAi(252) => b4_nUAi(252), b6_2ZTGIf_0
         => \b6_2ZTGIf[84]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(138), mdiclink_reg_0 => mdiclink_reg(29));
    
    b9_1LbcgKGUd : b8_1LbcQDr1_x_15_0
      port map(b4_nUAi(458) => b4_nUAi(458), b4_nUAi(457) => 
        b4_nUAi(457), b4_nUAi(456) => b4_nUAi(456), b6_2ZTGIf_0
         => \b6_2ZTGIf[152]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(7), mdiclink_reg_0 => mdiclink_reg(160));
    
    b8_1LbcgKbV : b8_1LbcQDr1_x_78_0
      port map(b4_nUAi(269) => b4_nUAi(269), b4_nUAi(268) => 
        b4_nUAi(268), b4_nUAi(267) => b4_nUAi(267), b6_2ZTGIf_0
         => \b6_2ZTGIf[89]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(132), mdiclink_reg_0 => mdiclink_reg(35));
    
    b7_1LbcgKG : b8_1LbcQDr1_x_166_0
      port map(b4_nUAi(5) => b4_nUAi(5), b4_nUAi(4) => b4_nUAi(4), 
        b4_nUAi(3) => b4_nUAi(3), b6_2ZTGIf_0 => \b6_2ZTGIf[1]\, 
        b11_OFWNT9L_8tZ_0 => b11_OFWNT9L_8tZ(105), mdiclink_reg_0
         => mdiclink_reg(62));
    
    b9_1LbcgKGUp : b8_1LbcQDr1_x_12_0
      port map(b4_nUAi(467) => b4_nUAi(467), b4_nUAi(466) => 
        b4_nUAi(466), b4_nUAi(465) => b4_nUAi(465), b6_2ZTGIf_0
         => \b6_2ZTGIf[155]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(60), mdiclink_reg_0 => mdiclink_reg(107));
    
    b8_1LbcgKJQ0 : b8_1LbcQDr1_x_73_0
      port map(b4_nUAi(284) => b4_nUAi(284), b4_nUAi(283) => 
        b4_nUAi(283), b4_nUAi(282) => b4_nUAi(282), b6_2ZTGIf_0
         => \b6_2ZTGIf[94]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(38), mdiclink_reg_0 => mdiclink_reg(129));
    
    b9_1LbcgKGId : b8_1LbcQDr1_x_45_0
      port map(b4_nUAi(368) => b4_nUAi(368), b4_nUAi(367) => 
        b4_nUAi(367), b4_nUAi(366) => b4_nUAi(366), b6_2ZTGIf_0
         => \b6_2ZTGIf[122]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(31), mdiclink_reg_0 => mdiclink_reg(136));
    
    b7_1LbcgKJ : b8_1LbcQDr1_x_158_0
      port map(b4_nUAi(29) => b4_nUAi(29), b4_nUAi(28) => 
        b4_nUAi(28), b4_nUAi(27) => b4_nUAi(27), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[9]\, b11_OFWNT9L_8tZ_0 => b11_OFWNT9L_8tZ(97), 
        mdiclink_reg_0 => mdiclink_reg(70));
    
    b9_1LbcgKGUq : b8_1LbcQDr1_x_8_0
      port map(b4_nUAi(479) => b4_nUAi(479), b4_nUAi(478) => 
        b4_nUAi(478), b4_nUAi(477) => b4_nUAi(477), b6_2ZTGIf_0
         => \b6_2ZTGIf[159]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(56), mdiclink_reg_0 => mdiclink_reg(111));
    
    b8_1LbcgKwn : b8_1LbcQDr1_x_139_0
      port map(b4_nUAi(86) => b4_nUAi(86), b4_nUAi(85) => 
        b4_nUAi(85), b4_nUAi(84) => b4_nUAi(84), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[28]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(130), mdiclink_reg_0 => mdiclink_reg(37));
    
    b9_1LbcgKGUS : b8_1LbcQDr1_x_9_0
      port map(b4_nUAi(476) => b4_nUAi(476), b4_nUAi(475) => 
        b4_nUAi(475), b4_nUAi(474) => b4_nUAi(474), b6_2ZTGIf_0
         => \b6_2ZTGIf[158]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(57), mdiclink_reg_0 => mdiclink_reg(110));
    
    b8_1LbcgKon : b8_1LbcQDr1_x_99_0
      port map(b4_nUAi(206) => b4_nUAi(206), b4_nUAi(205) => 
        b4_nUAi(205), b4_nUAi(204) => b4_nUAi(204), b6_2ZTGIf_0
         => \b6_2ZTGIf[68]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(155), mdiclink_reg_0 => mdiclink_reg(12));
    
    b8_1LbcgKJJ : b8_1LbcQDr1_x_70_0
      port map(b4_nUAi(293) => b4_nUAi(293), b4_nUAi(292) => 
        b4_nUAi(292), b4_nUAi(291) => b4_nUAi(291), b6_2ZTGIf_0
         => \b6_2ZTGIf[97]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(3), mdiclink_reg_0 => mdiclink_reg(164));
    
    b8_1LbcgKxq : b8_1LbcQDr1_x_94_0
      port map(b4_nUAi(221) => b4_nUAi(221), b4_nUAi(220) => 
        b4_nUAi(220), b4_nUAi(219) => b4_nUAi(219), b6_2ZTGIf_0
         => \b6_2ZTGIf[73]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(150), mdiclink_reg_0 => mdiclink_reg(17));
    
    b8_1LbcgKGq : b8_1LbcQDr1_x_154_0
      port map(b4_nUAi(41) => b4_nUAi(41), b4_nUAi(40) => 
        b4_nUAi(40), b4_nUAi(39) => b4_nUAi(39), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[13]\, b11_OFWNT9L_8tZ_0 => b11_OFWNT9L_8tZ(92), 
        mdiclink_reg_0 => mdiclink_reg(75));
    
    \b8_1LbcgKEq0\ : b8_1LbcQDr1_x_124_0
      port map(b4_nUAi(131) => b4_nUAi(131), b4_nUAi(130) => 
        b4_nUAi(130), b4_nUAi(129) => b4_nUAi(129), b6_2ZTGIf_0
         => \b6_2ZTGIf[43]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(75), mdiclink_reg_0 => mdiclink_reg(92));
    
    b9_1LbcgKGUe : b8_1LbcQDr1_x_10_0
      port map(b4_nUAi(473) => b4_nUAi(473), b4_nUAi(472) => 
        b4_nUAi(472), b4_nUAi(471) => b4_nUAi(471), b6_2ZTGIf_0
         => \b6_2ZTGIf[157]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(58), mdiclink_reg_0 => mdiclink_reg(109));
    
    b9_1LbcgKGIp : b8_1LbcQDr1_x_42_0
      port map(b4_nUAi(377) => b4_nUAi(377), b4_nUAi(376) => 
        b4_nUAi(376), b4_nUAi(375) => b4_nUAi(375), b6_2ZTGIf_0
         => \b6_2ZTGIf[125]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(28), mdiclink_reg_0 => mdiclink_reg(139));
    
    b8_1LbcgKIq : b8_1LbcQDr1_x_114_0
      port map(b4_nUAi(161) => b4_nUAi(161), b4_nUAi(160) => 
        b4_nUAi(160), b4_nUAi(159) => b4_nUAi(159), b6_2ZTGIf_0
         => \b6_2ZTGIf[53]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(65), mdiclink_reg_0 => mdiclink_reg(102));
    
    b8_1LbcgKwV : b8_1LbcQDr1_x_138_0
      port map(b4_nUAi(89) => b4_nUAi(89), b4_nUAi(88) => 
        b4_nUAi(88), b4_nUAi(87) => b4_nUAi(87), b6_2ZTGIf_0 => 
        \b6_2ZTGIf[29]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(129), mdiclink_reg_0 => mdiclink_reg(38));
    
    b9_1LbcgKGUm : b8_1LbcQDr1_x_17_0
      port map(b4_nUAi(452) => b4_nUAi(452), b4_nUAi(451) => 
        b4_nUAi(451), b4_nUAi(450) => b4_nUAi(450), b6_2ZTGIf_0
         => \b6_2ZTGIf[150]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(9), mdiclink_reg_0 => mdiclink_reg(158));
    
    b8_1LbcgKoV : b8_1LbcQDr1_x_98_0
      port map(b4_nUAi(209) => b4_nUAi(209), b4_nUAi(208) => 
        b4_nUAi(208), b4_nUAi(207) => b4_nUAi(207), b6_2ZTGIf_0
         => \b6_2ZTGIf[69]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(154), mdiclink_reg_0 => mdiclink_reg(13));
    
    b8_1LbcgKEA0 : b8_1LbcQDr1_x_121_0
      port map(b4_nUAi(140) => b4_nUAi(140), b4_nUAi(139) => 
        b4_nUAi(139), b4_nUAi(138) => b4_nUAi(138), b6_2ZTGIf_0
         => \b6_2ZTGIf[46]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(72), mdiclink_reg_0 => mdiclink_reg(95));
    
    b9_1LbcgKGIq : b8_1LbcQDr1_x_38_0
      port map(b4_nUAi(389) => b4_nUAi(389), b4_nUAi(388) => 
        b4_nUAi(388), b4_nUAi(387) => b4_nUAi(387), b6_2ZTGIf_0
         => \b6_2ZTGIf[129]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(16), mdiclink_reg_0 => mdiclink_reg(151));
    
    b8_1LbcgKbU : b8_1LbcQDr1_x_82_0
      port map(b4_nUAi(257) => b4_nUAi(257), b4_nUAi(256) => 
        b4_nUAi(256), b4_nUAi(255) => b4_nUAi(255), b6_2ZTGIf_0
         => \b6_2ZTGIf[85]\, b11_OFWNT9L_8tZ_0 => 
        b11_OFWNT9L_8tZ(137), mdiclink_reg_0 => mdiclink_reg(30));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_PfFzrNYI_x is

    port( b11_OFWNT9L_8tZ     : in    std_logic_vector(167 downto 0);
          mdiclink_reg        : in    std_logic_vector(167 downto 0);
          IICE_comm2iice_4    : in    std_logic;
          IICE_comm2iice_0    : in    std_logic;
          IICE_comm2iice_3    : in    std_logic;
          b10_nYBzIXrKbK_0    : out   std_logic;
          b7_PSyi_9u          : in    std_logic;
          b12_PSyi_XlK_qHv    : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic
        );

end b8_PfFzrNYI_x;

architecture DEF_ARCH of b8_PfFzrNYI_x is 

  component b5_nvmFL_504s_x_0
    port( b4_nUAi          : out   std_logic_vector(502 downto 0);
          IICE_comm2iice_4 : in    std_logic := 'U';
          IICE_comm2iice_0 : in    std_logic := 'U';
          IICE_comm2iice_3 : in    std_logic := 'U';
          b7_PSyi_9u       : in    std_logic := 'U';
          b12_PSyi_XlK_qHv : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component b13_PSyil9s1fkJ_L_x
    port( mdiclink_reg        : in    std_logic_vector(167 downto 0) := (others => 'U');
          b11_OFWNT9L_8tZ     : in    std_logic_vector(167 downto 0) := (others => 'U');
          b4_nUAi             : in    std_logic_vector(502 downto 0) := (others => 'U');
          b10_nYBzIXrKbK_0    : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          b12_PSyi_XlK_qHv    : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \b4_nUAi[0]\, \b4_nUAi[1]\, \b4_nUAi[2]\, 
        \b4_nUAi[3]\, \b4_nUAi[4]\, \b4_nUAi[5]\, \b4_nUAi[6]\, 
        \b4_nUAi[7]\, \b4_nUAi[8]\, \b4_nUAi[9]\, \b4_nUAi[10]\, 
        \b4_nUAi[11]\, \b4_nUAi[12]\, \b4_nUAi[13]\, 
        \b4_nUAi[14]\, \b4_nUAi[15]\, \b4_nUAi[16]\, 
        \b4_nUAi[17]\, \b4_nUAi[18]\, \b4_nUAi[19]\, 
        \b4_nUAi[20]\, \b4_nUAi[21]\, \b4_nUAi[22]\, 
        \b4_nUAi[23]\, \b4_nUAi[24]\, \b4_nUAi[25]\, 
        \b4_nUAi[26]\, \b4_nUAi[27]\, \b4_nUAi[28]\, 
        \b4_nUAi[29]\, \b4_nUAi[30]\, \b4_nUAi[31]\, 
        \b4_nUAi[32]\, \b4_nUAi[33]\, \b4_nUAi[34]\, 
        \b4_nUAi[35]\, \b4_nUAi[36]\, \b4_nUAi[37]\, 
        \b4_nUAi[38]\, \b4_nUAi[39]\, \b4_nUAi[40]\, 
        \b4_nUAi[41]\, \b4_nUAi[42]\, \b4_nUAi[43]\, 
        \b4_nUAi[44]\, \b4_nUAi[45]\, \b4_nUAi[46]\, 
        \b4_nUAi[47]\, \b4_nUAi[48]\, \b4_nUAi[49]\, 
        \b4_nUAi[50]\, \b4_nUAi[51]\, \b4_nUAi[52]\, 
        \b4_nUAi[53]\, \b4_nUAi[54]\, \b4_nUAi[55]\, 
        \b4_nUAi[56]\, \b4_nUAi[57]\, \b4_nUAi[58]\, 
        \b4_nUAi[59]\, \b4_nUAi[60]\, \b4_nUAi[61]\, 
        \b4_nUAi[62]\, \b4_nUAi[63]\, \b4_nUAi[64]\, 
        \b4_nUAi[65]\, \b4_nUAi[66]\, \b4_nUAi[67]\, 
        \b4_nUAi[68]\, \b4_nUAi[69]\, \b4_nUAi[70]\, 
        \b4_nUAi[71]\, \b4_nUAi[72]\, \b4_nUAi[73]\, 
        \b4_nUAi[74]\, \b4_nUAi[75]\, \b4_nUAi[76]\, 
        \b4_nUAi[77]\, \b4_nUAi[78]\, \b4_nUAi[79]\, 
        \b4_nUAi[80]\, \b4_nUAi[81]\, \b4_nUAi[82]\, 
        \b4_nUAi[83]\, \b4_nUAi[84]\, \b4_nUAi[85]\, 
        \b4_nUAi[86]\, \b4_nUAi[87]\, \b4_nUAi[88]\, 
        \b4_nUAi[89]\, \b4_nUAi[90]\, \b4_nUAi[91]\, 
        \b4_nUAi[92]\, \b4_nUAi[93]\, \b4_nUAi[94]\, 
        \b4_nUAi[95]\, \b4_nUAi[96]\, \b4_nUAi[97]\, 
        \b4_nUAi[98]\, \b4_nUAi[99]\, \b4_nUAi[100]\, 
        \b4_nUAi[101]\, \b4_nUAi[102]\, \b4_nUAi[103]\, 
        \b4_nUAi[104]\, \b4_nUAi[105]\, \b4_nUAi[106]\, 
        \b4_nUAi[107]\, \b4_nUAi[108]\, \b4_nUAi[109]\, 
        \b4_nUAi[110]\, \b4_nUAi[111]\, \b4_nUAi[112]\, 
        \b4_nUAi[113]\, \b4_nUAi[114]\, \b4_nUAi[115]\, 
        \b4_nUAi[116]\, \b4_nUAi[117]\, \b4_nUAi[118]\, 
        \b4_nUAi[119]\, \b4_nUAi[120]\, \b4_nUAi[121]\, 
        \b4_nUAi[122]\, \b4_nUAi[123]\, \b4_nUAi[124]\, 
        \b4_nUAi[125]\, \b4_nUAi[126]\, \b4_nUAi[127]\, 
        \b4_nUAi[128]\, \b4_nUAi[129]\, \b4_nUAi[130]\, 
        \b4_nUAi[131]\, \b4_nUAi[132]\, \b4_nUAi[133]\, 
        \b4_nUAi[134]\, \b4_nUAi[135]\, \b4_nUAi[136]\, 
        \b4_nUAi[137]\, \b4_nUAi[138]\, \b4_nUAi[139]\, 
        \b4_nUAi[140]\, \b4_nUAi[141]\, \b4_nUAi[142]\, 
        \b4_nUAi[143]\, \b4_nUAi[144]\, \b4_nUAi[145]\, 
        \b4_nUAi[146]\, \b4_nUAi[147]\, \b4_nUAi[148]\, 
        \b4_nUAi[149]\, \b4_nUAi[150]\, \b4_nUAi[151]\, 
        \b4_nUAi[152]\, \b4_nUAi[153]\, \b4_nUAi[154]\, 
        \b4_nUAi[155]\, \b4_nUAi[156]\, \b4_nUAi[157]\, 
        \b4_nUAi[158]\, \b4_nUAi[159]\, \b4_nUAi[160]\, 
        \b4_nUAi[161]\, \b4_nUAi[162]\, \b4_nUAi[163]\, 
        \b4_nUAi[164]\, \b4_nUAi[165]\, \b4_nUAi[166]\, 
        \b4_nUAi[167]\, \b4_nUAi[168]\, \b4_nUAi[169]\, 
        \b4_nUAi[170]\, \b4_nUAi[171]\, \b4_nUAi[172]\, 
        \b4_nUAi[173]\, \b4_nUAi[174]\, \b4_nUAi[175]\, 
        \b4_nUAi[176]\, \b4_nUAi[177]\, \b4_nUAi[178]\, 
        \b4_nUAi[179]\, \b4_nUAi[180]\, \b4_nUAi[181]\, 
        \b4_nUAi[182]\, \b4_nUAi[183]\, \b4_nUAi[184]\, 
        \b4_nUAi[185]\, \b4_nUAi[186]\, \b4_nUAi[187]\, 
        \b4_nUAi[188]\, \b4_nUAi[189]\, \b4_nUAi[190]\, 
        \b4_nUAi[191]\, \b4_nUAi[192]\, \b4_nUAi[193]\, 
        \b4_nUAi[194]\, \b4_nUAi[195]\, \b4_nUAi[196]\, 
        \b4_nUAi[197]\, \b4_nUAi[198]\, \b4_nUAi[199]\, 
        \b4_nUAi[200]\, \b4_nUAi[201]\, \b4_nUAi[202]\, 
        \b4_nUAi[203]\, \b4_nUAi[204]\, \b4_nUAi[205]\, 
        \b4_nUAi[206]\, \b4_nUAi[207]\, \b4_nUAi[208]\, 
        \b4_nUAi[209]\, \b4_nUAi[210]\, \b4_nUAi[211]\, 
        \b4_nUAi[212]\, \b4_nUAi[213]\, \b4_nUAi[214]\, 
        \b4_nUAi[215]\, \b4_nUAi[216]\, \b4_nUAi[217]\, 
        \b4_nUAi[218]\, \b4_nUAi[219]\, \b4_nUAi[220]\, 
        \b4_nUAi[221]\, \b4_nUAi[222]\, \b4_nUAi[223]\, 
        \b4_nUAi[224]\, \b4_nUAi[225]\, \b4_nUAi[226]\, 
        \b4_nUAi[227]\, \b4_nUAi[228]\, \b4_nUAi[229]\, 
        \b4_nUAi[230]\, \b4_nUAi[231]\, \b4_nUAi[232]\, 
        \b4_nUAi[233]\, \b4_nUAi[234]\, \b4_nUAi[235]\, 
        \b4_nUAi[236]\, \b4_nUAi[237]\, \b4_nUAi[238]\, 
        \b4_nUAi[239]\, \b4_nUAi[240]\, \b4_nUAi[241]\, 
        \b4_nUAi[242]\, \b4_nUAi[243]\, \b4_nUAi[244]\, 
        \b4_nUAi[245]\, \b4_nUAi[246]\, \b4_nUAi[247]\, 
        \b4_nUAi[248]\, \b4_nUAi[249]\, \b4_nUAi[250]\, 
        \b4_nUAi[251]\, \b4_nUAi[252]\, \b4_nUAi[253]\, 
        \b4_nUAi[254]\, \b4_nUAi[255]\, \b4_nUAi[256]\, 
        \b4_nUAi[257]\, \b4_nUAi[258]\, \b4_nUAi[259]\, 
        \b4_nUAi[260]\, \b4_nUAi[261]\, \b4_nUAi[262]\, 
        \b4_nUAi[263]\, \b4_nUAi[264]\, \b4_nUAi[265]\, 
        \b4_nUAi[266]\, \b4_nUAi[267]\, \b4_nUAi[268]\, 
        \b4_nUAi[269]\, \b4_nUAi[270]\, \b4_nUAi[271]\, 
        \b4_nUAi[272]\, \b4_nUAi[273]\, \b4_nUAi[274]\, 
        \b4_nUAi[275]\, \b4_nUAi[276]\, \b4_nUAi[277]\, 
        \b4_nUAi[278]\, \b4_nUAi[279]\, \b4_nUAi[280]\, 
        \b4_nUAi[281]\, \b4_nUAi[282]\, \b4_nUAi[283]\, 
        \b4_nUAi[284]\, \b4_nUAi[285]\, \b4_nUAi[286]\, 
        \b4_nUAi[287]\, \b4_nUAi[288]\, \b4_nUAi[289]\, 
        \b4_nUAi[290]\, \b4_nUAi[291]\, \b4_nUAi[292]\, 
        \b4_nUAi[293]\, \b4_nUAi[294]\, \b4_nUAi[295]\, 
        \b4_nUAi[296]\, \b4_nUAi[297]\, \b4_nUAi[298]\, 
        \b4_nUAi[299]\, \b4_nUAi[300]\, \b4_nUAi[301]\, 
        \b4_nUAi[302]\, \b4_nUAi[303]\, \b4_nUAi[304]\, 
        \b4_nUAi[305]\, \b4_nUAi[306]\, \b4_nUAi[307]\, 
        \b4_nUAi[308]\, \b4_nUAi[309]\, \b4_nUAi[310]\, 
        \b4_nUAi[311]\, \b4_nUAi[312]\, \b4_nUAi[313]\, 
        \b4_nUAi[314]\, \b4_nUAi[315]\, \b4_nUAi[316]\, 
        \b4_nUAi[317]\, \b4_nUAi[318]\, \b4_nUAi[319]\, 
        \b4_nUAi[320]\, \b4_nUAi[321]\, \b4_nUAi[322]\, 
        \b4_nUAi[323]\, \b4_nUAi[324]\, \b4_nUAi[325]\, 
        \b4_nUAi[326]\, \b4_nUAi[327]\, \b4_nUAi[328]\, 
        \b4_nUAi[329]\, \b4_nUAi[330]\, \b4_nUAi[331]\, 
        \b4_nUAi[332]\, \b4_nUAi[333]\, \b4_nUAi[334]\, 
        \b4_nUAi[335]\, \b4_nUAi[336]\, \b4_nUAi[337]\, 
        \b4_nUAi[338]\, \b4_nUAi[339]\, \b4_nUAi[340]\, 
        \b4_nUAi[341]\, \b4_nUAi[342]\, \b4_nUAi[343]\, 
        \b4_nUAi[344]\, \b4_nUAi[345]\, \b4_nUAi[346]\, 
        \b4_nUAi[347]\, \b4_nUAi[348]\, \b4_nUAi[349]\, 
        \b4_nUAi[350]\, \b4_nUAi[351]\, \b4_nUAi[352]\, 
        \b4_nUAi[353]\, \b4_nUAi[354]\, \b4_nUAi[355]\, 
        \b4_nUAi[356]\, \b4_nUAi[357]\, \b4_nUAi[358]\, 
        \b4_nUAi[359]\, \b4_nUAi[360]\, \b4_nUAi[361]\, 
        \b4_nUAi[362]\, \b4_nUAi[363]\, \b4_nUAi[364]\, 
        \b4_nUAi[365]\, \b4_nUAi[366]\, \b4_nUAi[367]\, 
        \b4_nUAi[368]\, \b4_nUAi[369]\, \b4_nUAi[370]\, 
        \b4_nUAi[371]\, \b4_nUAi[372]\, \b4_nUAi[373]\, 
        \b4_nUAi[374]\, \b4_nUAi[375]\, \b4_nUAi[376]\, 
        \b4_nUAi[377]\, \b4_nUAi[378]\, \b4_nUAi[379]\, 
        \b4_nUAi[380]\, \b4_nUAi[381]\, \b4_nUAi[382]\, 
        \b4_nUAi[383]\, \b4_nUAi[384]\, \b4_nUAi[385]\, 
        \b4_nUAi[386]\, \b4_nUAi[387]\, \b4_nUAi[388]\, 
        \b4_nUAi[389]\, \b4_nUAi[390]\, \b4_nUAi[391]\, 
        \b4_nUAi[392]\, \b4_nUAi[393]\, \b4_nUAi[394]\, 
        \b4_nUAi[395]\, \b4_nUAi[396]\, \b4_nUAi[397]\, 
        \b4_nUAi[398]\, \b4_nUAi[399]\, \b4_nUAi[400]\, 
        \b4_nUAi[401]\, \b4_nUAi[402]\, \b4_nUAi[403]\, 
        \b4_nUAi[404]\, \b4_nUAi[405]\, \b4_nUAi[406]\, 
        \b4_nUAi[407]\, \b4_nUAi[408]\, \b4_nUAi[409]\, 
        \b4_nUAi[410]\, \b4_nUAi[411]\, \b4_nUAi[412]\, 
        \b4_nUAi[413]\, \b4_nUAi[414]\, \b4_nUAi[415]\, 
        \b4_nUAi[416]\, \b4_nUAi[417]\, \b4_nUAi[418]\, 
        \b4_nUAi[419]\, \b4_nUAi[420]\, \b4_nUAi[421]\, 
        \b4_nUAi[422]\, \b4_nUAi[423]\, \b4_nUAi[424]\, 
        \b4_nUAi[425]\, \b4_nUAi[426]\, \b4_nUAi[427]\, 
        \b4_nUAi[428]\, \b4_nUAi[429]\, \b4_nUAi[430]\, 
        \b4_nUAi[431]\, \b4_nUAi[432]\, \b4_nUAi[433]\, 
        \b4_nUAi[434]\, \b4_nUAi[435]\, \b4_nUAi[436]\, 
        \b4_nUAi[437]\, \b4_nUAi[438]\, \b4_nUAi[439]\, 
        \b4_nUAi[440]\, \b4_nUAi[441]\, \b4_nUAi[442]\, 
        \b4_nUAi[443]\, \b4_nUAi[444]\, \b4_nUAi[445]\, 
        \b4_nUAi[446]\, \b4_nUAi[447]\, \b4_nUAi[448]\, 
        \b4_nUAi[449]\, \b4_nUAi[450]\, \b4_nUAi[451]\, 
        \b4_nUAi[452]\, \b4_nUAi[453]\, \b4_nUAi[454]\, 
        \b4_nUAi[455]\, \b4_nUAi[456]\, \b4_nUAi[457]\, 
        \b4_nUAi[458]\, \b4_nUAi[459]\, \b4_nUAi[460]\, 
        \b4_nUAi[461]\, \b4_nUAi[462]\, \b4_nUAi[463]\, 
        \b4_nUAi[464]\, \b4_nUAi[465]\, \b4_nUAi[466]\, 
        \b4_nUAi[467]\, \b4_nUAi[468]\, \b4_nUAi[469]\, 
        \b4_nUAi[470]\, \b4_nUAi[471]\, \b4_nUAi[472]\, 
        \b4_nUAi[473]\, \b4_nUAi[474]\, \b4_nUAi[475]\, 
        \b4_nUAi[476]\, \b4_nUAi[477]\, \b4_nUAi[478]\, 
        \b4_nUAi[479]\, \b4_nUAi[480]\, \b4_nUAi[481]\, 
        \b4_nUAi[482]\, \b4_nUAi[483]\, \b4_nUAi[484]\, 
        \b4_nUAi[485]\, \b4_nUAi[486]\, \b4_nUAi[487]\, 
        \b4_nUAi[488]\, \b4_nUAi[489]\, \b4_nUAi[490]\, 
        \b4_nUAi[491]\, \b4_nUAi[492]\, \b4_nUAi[493]\, 
        \b4_nUAi[494]\, \b4_nUAi[495]\, \b4_nUAi[496]\, 
        \b4_nUAi[497]\, \b4_nUAi[498]\, \b4_nUAi[499]\, 
        \b4_nUAi[500]\, \b4_nUAi[501]\, \b4_nUAi[502]\, 
        \b12_PSyi_XlK_qHv\, GND_net_1, VCC_net_1 : std_logic;

    for all : b5_nvmFL_504s_x_0
	Use entity work.b5_nvmFL_504s_x_0(DEF_ARCH);
    for all : b13_PSyil9s1fkJ_L_x
	Use entity work.b13_PSyil9s1fkJ_L_x(DEF_ARCH);
begin 

    b12_PSyi_XlK_qHv <= \b12_PSyi_XlK_qHv\;

    b5_PbrtL : b5_nvmFL_504s_x_0
      port map(b4_nUAi(502) => \b4_nUAi[502]\, b4_nUAi(501) => 
        \b4_nUAi[501]\, b4_nUAi(500) => \b4_nUAi[500]\, 
        b4_nUAi(499) => \b4_nUAi[499]\, b4_nUAi(498) => 
        \b4_nUAi[498]\, b4_nUAi(497) => \b4_nUAi[497]\, 
        b4_nUAi(496) => \b4_nUAi[496]\, b4_nUAi(495) => 
        \b4_nUAi[495]\, b4_nUAi(494) => \b4_nUAi[494]\, 
        b4_nUAi(493) => \b4_nUAi[493]\, b4_nUAi(492) => 
        \b4_nUAi[492]\, b4_nUAi(491) => \b4_nUAi[491]\, 
        b4_nUAi(490) => \b4_nUAi[490]\, b4_nUAi(489) => 
        \b4_nUAi[489]\, b4_nUAi(488) => \b4_nUAi[488]\, 
        b4_nUAi(487) => \b4_nUAi[487]\, b4_nUAi(486) => 
        \b4_nUAi[486]\, b4_nUAi(485) => \b4_nUAi[485]\, 
        b4_nUAi(484) => \b4_nUAi[484]\, b4_nUAi(483) => 
        \b4_nUAi[483]\, b4_nUAi(482) => \b4_nUAi[482]\, 
        b4_nUAi(481) => \b4_nUAi[481]\, b4_nUAi(480) => 
        \b4_nUAi[480]\, b4_nUAi(479) => \b4_nUAi[479]\, 
        b4_nUAi(478) => \b4_nUAi[478]\, b4_nUAi(477) => 
        \b4_nUAi[477]\, b4_nUAi(476) => \b4_nUAi[476]\, 
        b4_nUAi(475) => \b4_nUAi[475]\, b4_nUAi(474) => 
        \b4_nUAi[474]\, b4_nUAi(473) => \b4_nUAi[473]\, 
        b4_nUAi(472) => \b4_nUAi[472]\, b4_nUAi(471) => 
        \b4_nUAi[471]\, b4_nUAi(470) => \b4_nUAi[470]\, 
        b4_nUAi(469) => \b4_nUAi[469]\, b4_nUAi(468) => 
        \b4_nUAi[468]\, b4_nUAi(467) => \b4_nUAi[467]\, 
        b4_nUAi(466) => \b4_nUAi[466]\, b4_nUAi(465) => 
        \b4_nUAi[465]\, b4_nUAi(464) => \b4_nUAi[464]\, 
        b4_nUAi(463) => \b4_nUAi[463]\, b4_nUAi(462) => 
        \b4_nUAi[462]\, b4_nUAi(461) => \b4_nUAi[461]\, 
        b4_nUAi(460) => \b4_nUAi[460]\, b4_nUAi(459) => 
        \b4_nUAi[459]\, b4_nUAi(458) => \b4_nUAi[458]\, 
        b4_nUAi(457) => \b4_nUAi[457]\, b4_nUAi(456) => 
        \b4_nUAi[456]\, b4_nUAi(455) => \b4_nUAi[455]\, 
        b4_nUAi(454) => \b4_nUAi[454]\, b4_nUAi(453) => 
        \b4_nUAi[453]\, b4_nUAi(452) => \b4_nUAi[452]\, 
        b4_nUAi(451) => \b4_nUAi[451]\, b4_nUAi(450) => 
        \b4_nUAi[450]\, b4_nUAi(449) => \b4_nUAi[449]\, 
        b4_nUAi(448) => \b4_nUAi[448]\, b4_nUAi(447) => 
        \b4_nUAi[447]\, b4_nUAi(446) => \b4_nUAi[446]\, 
        b4_nUAi(445) => \b4_nUAi[445]\, b4_nUAi(444) => 
        \b4_nUAi[444]\, b4_nUAi(443) => \b4_nUAi[443]\, 
        b4_nUAi(442) => \b4_nUAi[442]\, b4_nUAi(441) => 
        \b4_nUAi[441]\, b4_nUAi(440) => \b4_nUAi[440]\, 
        b4_nUAi(439) => \b4_nUAi[439]\, b4_nUAi(438) => 
        \b4_nUAi[438]\, b4_nUAi(437) => \b4_nUAi[437]\, 
        b4_nUAi(436) => \b4_nUAi[436]\, b4_nUAi(435) => 
        \b4_nUAi[435]\, b4_nUAi(434) => \b4_nUAi[434]\, 
        b4_nUAi(433) => \b4_nUAi[433]\, b4_nUAi(432) => 
        \b4_nUAi[432]\, b4_nUAi(431) => \b4_nUAi[431]\, 
        b4_nUAi(430) => \b4_nUAi[430]\, b4_nUAi(429) => 
        \b4_nUAi[429]\, b4_nUAi(428) => \b4_nUAi[428]\, 
        b4_nUAi(427) => \b4_nUAi[427]\, b4_nUAi(426) => 
        \b4_nUAi[426]\, b4_nUAi(425) => \b4_nUAi[425]\, 
        b4_nUAi(424) => \b4_nUAi[424]\, b4_nUAi(423) => 
        \b4_nUAi[423]\, b4_nUAi(422) => \b4_nUAi[422]\, 
        b4_nUAi(421) => \b4_nUAi[421]\, b4_nUAi(420) => 
        \b4_nUAi[420]\, b4_nUAi(419) => \b4_nUAi[419]\, 
        b4_nUAi(418) => \b4_nUAi[418]\, b4_nUAi(417) => 
        \b4_nUAi[417]\, b4_nUAi(416) => \b4_nUAi[416]\, 
        b4_nUAi(415) => \b4_nUAi[415]\, b4_nUAi(414) => 
        \b4_nUAi[414]\, b4_nUAi(413) => \b4_nUAi[413]\, 
        b4_nUAi(412) => \b4_nUAi[412]\, b4_nUAi(411) => 
        \b4_nUAi[411]\, b4_nUAi(410) => \b4_nUAi[410]\, 
        b4_nUAi(409) => \b4_nUAi[409]\, b4_nUAi(408) => 
        \b4_nUAi[408]\, b4_nUAi(407) => \b4_nUAi[407]\, 
        b4_nUAi(406) => \b4_nUAi[406]\, b4_nUAi(405) => 
        \b4_nUAi[405]\, b4_nUAi(404) => \b4_nUAi[404]\, 
        b4_nUAi(403) => \b4_nUAi[403]\, b4_nUAi(402) => 
        \b4_nUAi[402]\, b4_nUAi(401) => \b4_nUAi[401]\, 
        b4_nUAi(400) => \b4_nUAi[400]\, b4_nUAi(399) => 
        \b4_nUAi[399]\, b4_nUAi(398) => \b4_nUAi[398]\, 
        b4_nUAi(397) => \b4_nUAi[397]\, b4_nUAi(396) => 
        \b4_nUAi[396]\, b4_nUAi(395) => \b4_nUAi[395]\, 
        b4_nUAi(394) => \b4_nUAi[394]\, b4_nUAi(393) => 
        \b4_nUAi[393]\, b4_nUAi(392) => \b4_nUAi[392]\, 
        b4_nUAi(391) => \b4_nUAi[391]\, b4_nUAi(390) => 
        \b4_nUAi[390]\, b4_nUAi(389) => \b4_nUAi[389]\, 
        b4_nUAi(388) => \b4_nUAi[388]\, b4_nUAi(387) => 
        \b4_nUAi[387]\, b4_nUAi(386) => \b4_nUAi[386]\, 
        b4_nUAi(385) => \b4_nUAi[385]\, b4_nUAi(384) => 
        \b4_nUAi[384]\, b4_nUAi(383) => \b4_nUAi[383]\, 
        b4_nUAi(382) => \b4_nUAi[382]\, b4_nUAi(381) => 
        \b4_nUAi[381]\, b4_nUAi(380) => \b4_nUAi[380]\, 
        b4_nUAi(379) => \b4_nUAi[379]\, b4_nUAi(378) => 
        \b4_nUAi[378]\, b4_nUAi(377) => \b4_nUAi[377]\, 
        b4_nUAi(376) => \b4_nUAi[376]\, b4_nUAi(375) => 
        \b4_nUAi[375]\, b4_nUAi(374) => \b4_nUAi[374]\, 
        b4_nUAi(373) => \b4_nUAi[373]\, b4_nUAi(372) => 
        \b4_nUAi[372]\, b4_nUAi(371) => \b4_nUAi[371]\, 
        b4_nUAi(370) => \b4_nUAi[370]\, b4_nUAi(369) => 
        \b4_nUAi[369]\, b4_nUAi(368) => \b4_nUAi[368]\, 
        b4_nUAi(367) => \b4_nUAi[367]\, b4_nUAi(366) => 
        \b4_nUAi[366]\, b4_nUAi(365) => \b4_nUAi[365]\, 
        b4_nUAi(364) => \b4_nUAi[364]\, b4_nUAi(363) => 
        \b4_nUAi[363]\, b4_nUAi(362) => \b4_nUAi[362]\, 
        b4_nUAi(361) => \b4_nUAi[361]\, b4_nUAi(360) => 
        \b4_nUAi[360]\, b4_nUAi(359) => \b4_nUAi[359]\, 
        b4_nUAi(358) => \b4_nUAi[358]\, b4_nUAi(357) => 
        \b4_nUAi[357]\, b4_nUAi(356) => \b4_nUAi[356]\, 
        b4_nUAi(355) => \b4_nUAi[355]\, b4_nUAi(354) => 
        \b4_nUAi[354]\, b4_nUAi(353) => \b4_nUAi[353]\, 
        b4_nUAi(352) => \b4_nUAi[352]\, b4_nUAi(351) => 
        \b4_nUAi[351]\, b4_nUAi(350) => \b4_nUAi[350]\, 
        b4_nUAi(349) => \b4_nUAi[349]\, b4_nUAi(348) => 
        \b4_nUAi[348]\, b4_nUAi(347) => \b4_nUAi[347]\, 
        b4_nUAi(346) => \b4_nUAi[346]\, b4_nUAi(345) => 
        \b4_nUAi[345]\, b4_nUAi(344) => \b4_nUAi[344]\, 
        b4_nUAi(343) => \b4_nUAi[343]\, b4_nUAi(342) => 
        \b4_nUAi[342]\, b4_nUAi(341) => \b4_nUAi[341]\, 
        b4_nUAi(340) => \b4_nUAi[340]\, b4_nUAi(339) => 
        \b4_nUAi[339]\, b4_nUAi(338) => \b4_nUAi[338]\, 
        b4_nUAi(337) => \b4_nUAi[337]\, b4_nUAi(336) => 
        \b4_nUAi[336]\, b4_nUAi(335) => \b4_nUAi[335]\, 
        b4_nUAi(334) => \b4_nUAi[334]\, b4_nUAi(333) => 
        \b4_nUAi[333]\, b4_nUAi(332) => \b4_nUAi[332]\, 
        b4_nUAi(331) => \b4_nUAi[331]\, b4_nUAi(330) => 
        \b4_nUAi[330]\, b4_nUAi(329) => \b4_nUAi[329]\, 
        b4_nUAi(328) => \b4_nUAi[328]\, b4_nUAi(327) => 
        \b4_nUAi[327]\, b4_nUAi(326) => \b4_nUAi[326]\, 
        b4_nUAi(325) => \b4_nUAi[325]\, b4_nUAi(324) => 
        \b4_nUAi[324]\, b4_nUAi(323) => \b4_nUAi[323]\, 
        b4_nUAi(322) => \b4_nUAi[322]\, b4_nUAi(321) => 
        \b4_nUAi[321]\, b4_nUAi(320) => \b4_nUAi[320]\, 
        b4_nUAi(319) => \b4_nUAi[319]\, b4_nUAi(318) => 
        \b4_nUAi[318]\, b4_nUAi(317) => \b4_nUAi[317]\, 
        b4_nUAi(316) => \b4_nUAi[316]\, b4_nUAi(315) => 
        \b4_nUAi[315]\, b4_nUAi(314) => \b4_nUAi[314]\, 
        b4_nUAi(313) => \b4_nUAi[313]\, b4_nUAi(312) => 
        \b4_nUAi[312]\, b4_nUAi(311) => \b4_nUAi[311]\, 
        b4_nUAi(310) => \b4_nUAi[310]\, b4_nUAi(309) => 
        \b4_nUAi[309]\, b4_nUAi(308) => \b4_nUAi[308]\, 
        b4_nUAi(307) => \b4_nUAi[307]\, b4_nUAi(306) => 
        \b4_nUAi[306]\, b4_nUAi(305) => \b4_nUAi[305]\, 
        b4_nUAi(304) => \b4_nUAi[304]\, b4_nUAi(303) => 
        \b4_nUAi[303]\, b4_nUAi(302) => \b4_nUAi[302]\, 
        b4_nUAi(301) => \b4_nUAi[301]\, b4_nUAi(300) => 
        \b4_nUAi[300]\, b4_nUAi(299) => \b4_nUAi[299]\, 
        b4_nUAi(298) => \b4_nUAi[298]\, b4_nUAi(297) => 
        \b4_nUAi[297]\, b4_nUAi(296) => \b4_nUAi[296]\, 
        b4_nUAi(295) => \b4_nUAi[295]\, b4_nUAi(294) => 
        \b4_nUAi[294]\, b4_nUAi(293) => \b4_nUAi[293]\, 
        b4_nUAi(292) => \b4_nUAi[292]\, b4_nUAi(291) => 
        \b4_nUAi[291]\, b4_nUAi(290) => \b4_nUAi[290]\, 
        b4_nUAi(289) => \b4_nUAi[289]\, b4_nUAi(288) => 
        \b4_nUAi[288]\, b4_nUAi(287) => \b4_nUAi[287]\, 
        b4_nUAi(286) => \b4_nUAi[286]\, b4_nUAi(285) => 
        \b4_nUAi[285]\, b4_nUAi(284) => \b4_nUAi[284]\, 
        b4_nUAi(283) => \b4_nUAi[283]\, b4_nUAi(282) => 
        \b4_nUAi[282]\, b4_nUAi(281) => \b4_nUAi[281]\, 
        b4_nUAi(280) => \b4_nUAi[280]\, b4_nUAi(279) => 
        \b4_nUAi[279]\, b4_nUAi(278) => \b4_nUAi[278]\, 
        b4_nUAi(277) => \b4_nUAi[277]\, b4_nUAi(276) => 
        \b4_nUAi[276]\, b4_nUAi(275) => \b4_nUAi[275]\, 
        b4_nUAi(274) => \b4_nUAi[274]\, b4_nUAi(273) => 
        \b4_nUAi[273]\, b4_nUAi(272) => \b4_nUAi[272]\, 
        b4_nUAi(271) => \b4_nUAi[271]\, b4_nUAi(270) => 
        \b4_nUAi[270]\, b4_nUAi(269) => \b4_nUAi[269]\, 
        b4_nUAi(268) => \b4_nUAi[268]\, b4_nUAi(267) => 
        \b4_nUAi[267]\, b4_nUAi(266) => \b4_nUAi[266]\, 
        b4_nUAi(265) => \b4_nUAi[265]\, b4_nUAi(264) => 
        \b4_nUAi[264]\, b4_nUAi(263) => \b4_nUAi[263]\, 
        b4_nUAi(262) => \b4_nUAi[262]\, b4_nUAi(261) => 
        \b4_nUAi[261]\, b4_nUAi(260) => \b4_nUAi[260]\, 
        b4_nUAi(259) => \b4_nUAi[259]\, b4_nUAi(258) => 
        \b4_nUAi[258]\, b4_nUAi(257) => \b4_nUAi[257]\, 
        b4_nUAi(256) => \b4_nUAi[256]\, b4_nUAi(255) => 
        \b4_nUAi[255]\, b4_nUAi(254) => \b4_nUAi[254]\, 
        b4_nUAi(253) => \b4_nUAi[253]\, b4_nUAi(252) => 
        \b4_nUAi[252]\, b4_nUAi(251) => \b4_nUAi[251]\, 
        b4_nUAi(250) => \b4_nUAi[250]\, b4_nUAi(249) => 
        \b4_nUAi[249]\, b4_nUAi(248) => \b4_nUAi[248]\, 
        b4_nUAi(247) => \b4_nUAi[247]\, b4_nUAi(246) => 
        \b4_nUAi[246]\, b4_nUAi(245) => \b4_nUAi[245]\, 
        b4_nUAi(244) => \b4_nUAi[244]\, b4_nUAi(243) => 
        \b4_nUAi[243]\, b4_nUAi(242) => \b4_nUAi[242]\, 
        b4_nUAi(241) => \b4_nUAi[241]\, b4_nUAi(240) => 
        \b4_nUAi[240]\, b4_nUAi(239) => \b4_nUAi[239]\, 
        b4_nUAi(238) => \b4_nUAi[238]\, b4_nUAi(237) => 
        \b4_nUAi[237]\, b4_nUAi(236) => \b4_nUAi[236]\, 
        b4_nUAi(235) => \b4_nUAi[235]\, b4_nUAi(234) => 
        \b4_nUAi[234]\, b4_nUAi(233) => \b4_nUAi[233]\, 
        b4_nUAi(232) => \b4_nUAi[232]\, b4_nUAi(231) => 
        \b4_nUAi[231]\, b4_nUAi(230) => \b4_nUAi[230]\, 
        b4_nUAi(229) => \b4_nUAi[229]\, b4_nUAi(228) => 
        \b4_nUAi[228]\, b4_nUAi(227) => \b4_nUAi[227]\, 
        b4_nUAi(226) => \b4_nUAi[226]\, b4_nUAi(225) => 
        \b4_nUAi[225]\, b4_nUAi(224) => \b4_nUAi[224]\, 
        b4_nUAi(223) => \b4_nUAi[223]\, b4_nUAi(222) => 
        \b4_nUAi[222]\, b4_nUAi(221) => \b4_nUAi[221]\, 
        b4_nUAi(220) => \b4_nUAi[220]\, b4_nUAi(219) => 
        \b4_nUAi[219]\, b4_nUAi(218) => \b4_nUAi[218]\, 
        b4_nUAi(217) => \b4_nUAi[217]\, b4_nUAi(216) => 
        \b4_nUAi[216]\, b4_nUAi(215) => \b4_nUAi[215]\, 
        b4_nUAi(214) => \b4_nUAi[214]\, b4_nUAi(213) => 
        \b4_nUAi[213]\, b4_nUAi(212) => \b4_nUAi[212]\, 
        b4_nUAi(211) => \b4_nUAi[211]\, b4_nUAi(210) => 
        \b4_nUAi[210]\, b4_nUAi(209) => \b4_nUAi[209]\, 
        b4_nUAi(208) => \b4_nUAi[208]\, b4_nUAi(207) => 
        \b4_nUAi[207]\, b4_nUAi(206) => \b4_nUAi[206]\, 
        b4_nUAi(205) => \b4_nUAi[205]\, b4_nUAi(204) => 
        \b4_nUAi[204]\, b4_nUAi(203) => \b4_nUAi[203]\, 
        b4_nUAi(202) => \b4_nUAi[202]\, b4_nUAi(201) => 
        \b4_nUAi[201]\, b4_nUAi(200) => \b4_nUAi[200]\, 
        b4_nUAi(199) => \b4_nUAi[199]\, b4_nUAi(198) => 
        \b4_nUAi[198]\, b4_nUAi(197) => \b4_nUAi[197]\, 
        b4_nUAi(196) => \b4_nUAi[196]\, b4_nUAi(195) => 
        \b4_nUAi[195]\, b4_nUAi(194) => \b4_nUAi[194]\, 
        b4_nUAi(193) => \b4_nUAi[193]\, b4_nUAi(192) => 
        \b4_nUAi[192]\, b4_nUAi(191) => \b4_nUAi[191]\, 
        b4_nUAi(190) => \b4_nUAi[190]\, b4_nUAi(189) => 
        \b4_nUAi[189]\, b4_nUAi(188) => \b4_nUAi[188]\, 
        b4_nUAi(187) => \b4_nUAi[187]\, b4_nUAi(186) => 
        \b4_nUAi[186]\, b4_nUAi(185) => \b4_nUAi[185]\, 
        b4_nUAi(184) => \b4_nUAi[184]\, b4_nUAi(183) => 
        \b4_nUAi[183]\, b4_nUAi(182) => \b4_nUAi[182]\, 
        b4_nUAi(181) => \b4_nUAi[181]\, b4_nUAi(180) => 
        \b4_nUAi[180]\, b4_nUAi(179) => \b4_nUAi[179]\, 
        b4_nUAi(178) => \b4_nUAi[178]\, b4_nUAi(177) => 
        \b4_nUAi[177]\, b4_nUAi(176) => \b4_nUAi[176]\, 
        b4_nUAi(175) => \b4_nUAi[175]\, b4_nUAi(174) => 
        \b4_nUAi[174]\, b4_nUAi(173) => \b4_nUAi[173]\, 
        b4_nUAi(172) => \b4_nUAi[172]\, b4_nUAi(171) => 
        \b4_nUAi[171]\, b4_nUAi(170) => \b4_nUAi[170]\, 
        b4_nUAi(169) => \b4_nUAi[169]\, b4_nUAi(168) => 
        \b4_nUAi[168]\, b4_nUAi(167) => \b4_nUAi[167]\, 
        b4_nUAi(166) => \b4_nUAi[166]\, b4_nUAi(165) => 
        \b4_nUAi[165]\, b4_nUAi(164) => \b4_nUAi[164]\, 
        b4_nUAi(163) => \b4_nUAi[163]\, b4_nUAi(162) => 
        \b4_nUAi[162]\, b4_nUAi(161) => \b4_nUAi[161]\, 
        b4_nUAi(160) => \b4_nUAi[160]\, b4_nUAi(159) => 
        \b4_nUAi[159]\, b4_nUAi(158) => \b4_nUAi[158]\, 
        b4_nUAi(157) => \b4_nUAi[157]\, b4_nUAi(156) => 
        \b4_nUAi[156]\, b4_nUAi(155) => \b4_nUAi[155]\, 
        b4_nUAi(154) => \b4_nUAi[154]\, b4_nUAi(153) => 
        \b4_nUAi[153]\, b4_nUAi(152) => \b4_nUAi[152]\, 
        b4_nUAi(151) => \b4_nUAi[151]\, b4_nUAi(150) => 
        \b4_nUAi[150]\, b4_nUAi(149) => \b4_nUAi[149]\, 
        b4_nUAi(148) => \b4_nUAi[148]\, b4_nUAi(147) => 
        \b4_nUAi[147]\, b4_nUAi(146) => \b4_nUAi[146]\, 
        b4_nUAi(145) => \b4_nUAi[145]\, b4_nUAi(144) => 
        \b4_nUAi[144]\, b4_nUAi(143) => \b4_nUAi[143]\, 
        b4_nUAi(142) => \b4_nUAi[142]\, b4_nUAi(141) => 
        \b4_nUAi[141]\, b4_nUAi(140) => \b4_nUAi[140]\, 
        b4_nUAi(139) => \b4_nUAi[139]\, b4_nUAi(138) => 
        \b4_nUAi[138]\, b4_nUAi(137) => \b4_nUAi[137]\, 
        b4_nUAi(136) => \b4_nUAi[136]\, b4_nUAi(135) => 
        \b4_nUAi[135]\, b4_nUAi(134) => \b4_nUAi[134]\, 
        b4_nUAi(133) => \b4_nUAi[133]\, b4_nUAi(132) => 
        \b4_nUAi[132]\, b4_nUAi(131) => \b4_nUAi[131]\, 
        b4_nUAi(130) => \b4_nUAi[130]\, b4_nUAi(129) => 
        \b4_nUAi[129]\, b4_nUAi(128) => \b4_nUAi[128]\, 
        b4_nUAi(127) => \b4_nUAi[127]\, b4_nUAi(126) => 
        \b4_nUAi[126]\, b4_nUAi(125) => \b4_nUAi[125]\, 
        b4_nUAi(124) => \b4_nUAi[124]\, b4_nUAi(123) => 
        \b4_nUAi[123]\, b4_nUAi(122) => \b4_nUAi[122]\, 
        b4_nUAi(121) => \b4_nUAi[121]\, b4_nUAi(120) => 
        \b4_nUAi[120]\, b4_nUAi(119) => \b4_nUAi[119]\, 
        b4_nUAi(118) => \b4_nUAi[118]\, b4_nUAi(117) => 
        \b4_nUAi[117]\, b4_nUAi(116) => \b4_nUAi[116]\, 
        b4_nUAi(115) => \b4_nUAi[115]\, b4_nUAi(114) => 
        \b4_nUAi[114]\, b4_nUAi(113) => \b4_nUAi[113]\, 
        b4_nUAi(112) => \b4_nUAi[112]\, b4_nUAi(111) => 
        \b4_nUAi[111]\, b4_nUAi(110) => \b4_nUAi[110]\, 
        b4_nUAi(109) => \b4_nUAi[109]\, b4_nUAi(108) => 
        \b4_nUAi[108]\, b4_nUAi(107) => \b4_nUAi[107]\, 
        b4_nUAi(106) => \b4_nUAi[106]\, b4_nUAi(105) => 
        \b4_nUAi[105]\, b4_nUAi(104) => \b4_nUAi[104]\, 
        b4_nUAi(103) => \b4_nUAi[103]\, b4_nUAi(102) => 
        \b4_nUAi[102]\, b4_nUAi(101) => \b4_nUAi[101]\, 
        b4_nUAi(100) => \b4_nUAi[100]\, b4_nUAi(99) => 
        \b4_nUAi[99]\, b4_nUAi(98) => \b4_nUAi[98]\, b4_nUAi(97)
         => \b4_nUAi[97]\, b4_nUAi(96) => \b4_nUAi[96]\, 
        b4_nUAi(95) => \b4_nUAi[95]\, b4_nUAi(94) => 
        \b4_nUAi[94]\, b4_nUAi(93) => \b4_nUAi[93]\, b4_nUAi(92)
         => \b4_nUAi[92]\, b4_nUAi(91) => \b4_nUAi[91]\, 
        b4_nUAi(90) => \b4_nUAi[90]\, b4_nUAi(89) => 
        \b4_nUAi[89]\, b4_nUAi(88) => \b4_nUAi[88]\, b4_nUAi(87)
         => \b4_nUAi[87]\, b4_nUAi(86) => \b4_nUAi[86]\, 
        b4_nUAi(85) => \b4_nUAi[85]\, b4_nUAi(84) => 
        \b4_nUAi[84]\, b4_nUAi(83) => \b4_nUAi[83]\, b4_nUAi(82)
         => \b4_nUAi[82]\, b4_nUAi(81) => \b4_nUAi[81]\, 
        b4_nUAi(80) => \b4_nUAi[80]\, b4_nUAi(79) => 
        \b4_nUAi[79]\, b4_nUAi(78) => \b4_nUAi[78]\, b4_nUAi(77)
         => \b4_nUAi[77]\, b4_nUAi(76) => \b4_nUAi[76]\, 
        b4_nUAi(75) => \b4_nUAi[75]\, b4_nUAi(74) => 
        \b4_nUAi[74]\, b4_nUAi(73) => \b4_nUAi[73]\, b4_nUAi(72)
         => \b4_nUAi[72]\, b4_nUAi(71) => \b4_nUAi[71]\, 
        b4_nUAi(70) => \b4_nUAi[70]\, b4_nUAi(69) => 
        \b4_nUAi[69]\, b4_nUAi(68) => \b4_nUAi[68]\, b4_nUAi(67)
         => \b4_nUAi[67]\, b4_nUAi(66) => \b4_nUAi[66]\, 
        b4_nUAi(65) => \b4_nUAi[65]\, b4_nUAi(64) => 
        \b4_nUAi[64]\, b4_nUAi(63) => \b4_nUAi[63]\, b4_nUAi(62)
         => \b4_nUAi[62]\, b4_nUAi(61) => \b4_nUAi[61]\, 
        b4_nUAi(60) => \b4_nUAi[60]\, b4_nUAi(59) => 
        \b4_nUAi[59]\, b4_nUAi(58) => \b4_nUAi[58]\, b4_nUAi(57)
         => \b4_nUAi[57]\, b4_nUAi(56) => \b4_nUAi[56]\, 
        b4_nUAi(55) => \b4_nUAi[55]\, b4_nUAi(54) => 
        \b4_nUAi[54]\, b4_nUAi(53) => \b4_nUAi[53]\, b4_nUAi(52)
         => \b4_nUAi[52]\, b4_nUAi(51) => \b4_nUAi[51]\, 
        b4_nUAi(50) => \b4_nUAi[50]\, b4_nUAi(49) => 
        \b4_nUAi[49]\, b4_nUAi(48) => \b4_nUAi[48]\, b4_nUAi(47)
         => \b4_nUAi[47]\, b4_nUAi(46) => \b4_nUAi[46]\, 
        b4_nUAi(45) => \b4_nUAi[45]\, b4_nUAi(44) => 
        \b4_nUAi[44]\, b4_nUAi(43) => \b4_nUAi[43]\, b4_nUAi(42)
         => \b4_nUAi[42]\, b4_nUAi(41) => \b4_nUAi[41]\, 
        b4_nUAi(40) => \b4_nUAi[40]\, b4_nUAi(39) => 
        \b4_nUAi[39]\, b4_nUAi(38) => \b4_nUAi[38]\, b4_nUAi(37)
         => \b4_nUAi[37]\, b4_nUAi(36) => \b4_nUAi[36]\, 
        b4_nUAi(35) => \b4_nUAi[35]\, b4_nUAi(34) => 
        \b4_nUAi[34]\, b4_nUAi(33) => \b4_nUAi[33]\, b4_nUAi(32)
         => \b4_nUAi[32]\, b4_nUAi(31) => \b4_nUAi[31]\, 
        b4_nUAi(30) => \b4_nUAi[30]\, b4_nUAi(29) => 
        \b4_nUAi[29]\, b4_nUAi(28) => \b4_nUAi[28]\, b4_nUAi(27)
         => \b4_nUAi[27]\, b4_nUAi(26) => \b4_nUAi[26]\, 
        b4_nUAi(25) => \b4_nUAi[25]\, b4_nUAi(24) => 
        \b4_nUAi[24]\, b4_nUAi(23) => \b4_nUAi[23]\, b4_nUAi(22)
         => \b4_nUAi[22]\, b4_nUAi(21) => \b4_nUAi[21]\, 
        b4_nUAi(20) => \b4_nUAi[20]\, b4_nUAi(19) => 
        \b4_nUAi[19]\, b4_nUAi(18) => \b4_nUAi[18]\, b4_nUAi(17)
         => \b4_nUAi[17]\, b4_nUAi(16) => \b4_nUAi[16]\, 
        b4_nUAi(15) => \b4_nUAi[15]\, b4_nUAi(14) => 
        \b4_nUAi[14]\, b4_nUAi(13) => \b4_nUAi[13]\, b4_nUAi(12)
         => \b4_nUAi[12]\, b4_nUAi(11) => \b4_nUAi[11]\, 
        b4_nUAi(10) => \b4_nUAi[10]\, b4_nUAi(9) => \b4_nUAi[9]\, 
        b4_nUAi(8) => \b4_nUAi[8]\, b4_nUAi(7) => \b4_nUAi[7]\, 
        b4_nUAi(6) => \b4_nUAi[6]\, b4_nUAi(5) => \b4_nUAi[5]\, 
        b4_nUAi(4) => \b4_nUAi[4]\, b4_nUAi(3) => \b4_nUAi[3]\, 
        b4_nUAi(2) => \b4_nUAi[2]\, b4_nUAi(1) => \b4_nUAi[1]\, 
        b4_nUAi(0) => \b4_nUAi[0]\, IICE_comm2iice_4 => 
        IICE_comm2iice_4, IICE_comm2iice_0 => IICE_comm2iice_0, 
        IICE_comm2iice_3 => IICE_comm2iice_3, b7_PSyi_9u => 
        b7_PSyi_9u, b12_PSyi_XlK_qHv => \b12_PSyi_XlK_qHv\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b7_PbTtl9G : b13_PSyil9s1fkJ_L_x
      port map(mdiclink_reg(167) => mdiclink_reg(167), 
        mdiclink_reg(166) => mdiclink_reg(166), mdiclink_reg(165)
         => mdiclink_reg(165), mdiclink_reg(164) => 
        mdiclink_reg(164), mdiclink_reg(163) => mdiclink_reg(163), 
        mdiclink_reg(162) => mdiclink_reg(162), mdiclink_reg(161)
         => mdiclink_reg(161), mdiclink_reg(160) => 
        mdiclink_reg(160), mdiclink_reg(159) => mdiclink_reg(159), 
        mdiclink_reg(158) => mdiclink_reg(158), mdiclink_reg(157)
         => mdiclink_reg(157), mdiclink_reg(156) => 
        mdiclink_reg(156), mdiclink_reg(155) => mdiclink_reg(155), 
        mdiclink_reg(154) => mdiclink_reg(154), mdiclink_reg(153)
         => mdiclink_reg(153), mdiclink_reg(152) => 
        mdiclink_reg(152), mdiclink_reg(151) => mdiclink_reg(151), 
        mdiclink_reg(150) => mdiclink_reg(150), mdiclink_reg(149)
         => mdiclink_reg(149), mdiclink_reg(148) => 
        mdiclink_reg(148), mdiclink_reg(147) => mdiclink_reg(147), 
        mdiclink_reg(146) => mdiclink_reg(146), mdiclink_reg(145)
         => mdiclink_reg(145), mdiclink_reg(144) => 
        mdiclink_reg(144), mdiclink_reg(143) => mdiclink_reg(143), 
        mdiclink_reg(142) => mdiclink_reg(142), mdiclink_reg(141)
         => mdiclink_reg(141), mdiclink_reg(140) => 
        mdiclink_reg(140), mdiclink_reg(139) => mdiclink_reg(139), 
        mdiclink_reg(138) => mdiclink_reg(138), mdiclink_reg(137)
         => mdiclink_reg(137), mdiclink_reg(136) => 
        mdiclink_reg(136), mdiclink_reg(135) => mdiclink_reg(135), 
        mdiclink_reg(134) => mdiclink_reg(134), mdiclink_reg(133)
         => mdiclink_reg(133), mdiclink_reg(132) => 
        mdiclink_reg(132), mdiclink_reg(131) => mdiclink_reg(131), 
        mdiclink_reg(130) => mdiclink_reg(130), mdiclink_reg(129)
         => mdiclink_reg(129), mdiclink_reg(128) => 
        mdiclink_reg(128), mdiclink_reg(127) => mdiclink_reg(127), 
        mdiclink_reg(126) => mdiclink_reg(126), mdiclink_reg(125)
         => mdiclink_reg(125), mdiclink_reg(124) => 
        mdiclink_reg(124), mdiclink_reg(123) => mdiclink_reg(123), 
        mdiclink_reg(122) => mdiclink_reg(122), mdiclink_reg(121)
         => mdiclink_reg(121), mdiclink_reg(120) => 
        mdiclink_reg(120), mdiclink_reg(119) => mdiclink_reg(119), 
        mdiclink_reg(118) => mdiclink_reg(118), mdiclink_reg(117)
         => mdiclink_reg(117), mdiclink_reg(116) => 
        mdiclink_reg(116), mdiclink_reg(115) => mdiclink_reg(115), 
        mdiclink_reg(114) => mdiclink_reg(114), mdiclink_reg(113)
         => mdiclink_reg(113), mdiclink_reg(112) => 
        mdiclink_reg(112), mdiclink_reg(111) => mdiclink_reg(111), 
        mdiclink_reg(110) => mdiclink_reg(110), mdiclink_reg(109)
         => mdiclink_reg(109), mdiclink_reg(108) => 
        mdiclink_reg(108), mdiclink_reg(107) => mdiclink_reg(107), 
        mdiclink_reg(106) => mdiclink_reg(106), mdiclink_reg(105)
         => mdiclink_reg(105), mdiclink_reg(104) => 
        mdiclink_reg(104), mdiclink_reg(103) => mdiclink_reg(103), 
        mdiclink_reg(102) => mdiclink_reg(102), mdiclink_reg(101)
         => mdiclink_reg(101), mdiclink_reg(100) => 
        mdiclink_reg(100), mdiclink_reg(99) => mdiclink_reg(99), 
        mdiclink_reg(98) => mdiclink_reg(98), mdiclink_reg(97)
         => mdiclink_reg(97), mdiclink_reg(96) => 
        mdiclink_reg(96), mdiclink_reg(95) => mdiclink_reg(95), 
        mdiclink_reg(94) => mdiclink_reg(94), mdiclink_reg(93)
         => mdiclink_reg(93), mdiclink_reg(92) => 
        mdiclink_reg(92), mdiclink_reg(91) => mdiclink_reg(91), 
        mdiclink_reg(90) => mdiclink_reg(90), mdiclink_reg(89)
         => mdiclink_reg(89), mdiclink_reg(88) => 
        mdiclink_reg(88), mdiclink_reg(87) => mdiclink_reg(87), 
        mdiclink_reg(86) => mdiclink_reg(86), mdiclink_reg(85)
         => mdiclink_reg(85), mdiclink_reg(84) => 
        mdiclink_reg(84), mdiclink_reg(83) => mdiclink_reg(83), 
        mdiclink_reg(82) => mdiclink_reg(82), mdiclink_reg(81)
         => mdiclink_reg(81), mdiclink_reg(80) => 
        mdiclink_reg(80), mdiclink_reg(79) => mdiclink_reg(79), 
        mdiclink_reg(78) => mdiclink_reg(78), mdiclink_reg(77)
         => mdiclink_reg(77), mdiclink_reg(76) => 
        mdiclink_reg(76), mdiclink_reg(75) => mdiclink_reg(75), 
        mdiclink_reg(74) => mdiclink_reg(74), mdiclink_reg(73)
         => mdiclink_reg(73), mdiclink_reg(72) => 
        mdiclink_reg(72), mdiclink_reg(71) => mdiclink_reg(71), 
        mdiclink_reg(70) => mdiclink_reg(70), mdiclink_reg(69)
         => mdiclink_reg(69), mdiclink_reg(68) => 
        mdiclink_reg(68), mdiclink_reg(67) => mdiclink_reg(67), 
        mdiclink_reg(66) => mdiclink_reg(66), mdiclink_reg(65)
         => mdiclink_reg(65), mdiclink_reg(64) => 
        mdiclink_reg(64), mdiclink_reg(63) => mdiclink_reg(63), 
        mdiclink_reg(62) => mdiclink_reg(62), mdiclink_reg(61)
         => mdiclink_reg(61), mdiclink_reg(60) => 
        mdiclink_reg(60), mdiclink_reg(59) => mdiclink_reg(59), 
        mdiclink_reg(58) => mdiclink_reg(58), mdiclink_reg(57)
         => mdiclink_reg(57), mdiclink_reg(56) => 
        mdiclink_reg(56), mdiclink_reg(55) => mdiclink_reg(55), 
        mdiclink_reg(54) => mdiclink_reg(54), mdiclink_reg(53)
         => mdiclink_reg(53), mdiclink_reg(52) => 
        mdiclink_reg(52), mdiclink_reg(51) => mdiclink_reg(51), 
        mdiclink_reg(50) => mdiclink_reg(50), mdiclink_reg(49)
         => mdiclink_reg(49), mdiclink_reg(48) => 
        mdiclink_reg(48), mdiclink_reg(47) => mdiclink_reg(47), 
        mdiclink_reg(46) => mdiclink_reg(46), mdiclink_reg(45)
         => mdiclink_reg(45), mdiclink_reg(44) => 
        mdiclink_reg(44), mdiclink_reg(43) => mdiclink_reg(43), 
        mdiclink_reg(42) => mdiclink_reg(42), mdiclink_reg(41)
         => mdiclink_reg(41), mdiclink_reg(40) => 
        mdiclink_reg(40), mdiclink_reg(39) => mdiclink_reg(39), 
        mdiclink_reg(38) => mdiclink_reg(38), mdiclink_reg(37)
         => mdiclink_reg(37), mdiclink_reg(36) => 
        mdiclink_reg(36), mdiclink_reg(35) => mdiclink_reg(35), 
        mdiclink_reg(34) => mdiclink_reg(34), mdiclink_reg(33)
         => mdiclink_reg(33), mdiclink_reg(32) => 
        mdiclink_reg(32), mdiclink_reg(31) => mdiclink_reg(31), 
        mdiclink_reg(30) => mdiclink_reg(30), mdiclink_reg(29)
         => mdiclink_reg(29), mdiclink_reg(28) => 
        mdiclink_reg(28), mdiclink_reg(27) => mdiclink_reg(27), 
        mdiclink_reg(26) => mdiclink_reg(26), mdiclink_reg(25)
         => mdiclink_reg(25), mdiclink_reg(24) => 
        mdiclink_reg(24), mdiclink_reg(23) => mdiclink_reg(23), 
        mdiclink_reg(22) => mdiclink_reg(22), mdiclink_reg(21)
         => mdiclink_reg(21), mdiclink_reg(20) => 
        mdiclink_reg(20), mdiclink_reg(19) => mdiclink_reg(19), 
        mdiclink_reg(18) => mdiclink_reg(18), mdiclink_reg(17)
         => mdiclink_reg(17), mdiclink_reg(16) => 
        mdiclink_reg(16), mdiclink_reg(15) => mdiclink_reg(15), 
        mdiclink_reg(14) => mdiclink_reg(14), mdiclink_reg(13)
         => mdiclink_reg(13), mdiclink_reg(12) => 
        mdiclink_reg(12), mdiclink_reg(11) => mdiclink_reg(11), 
        mdiclink_reg(10) => mdiclink_reg(10), mdiclink_reg(9) => 
        mdiclink_reg(9), mdiclink_reg(8) => mdiclink_reg(8), 
        mdiclink_reg(7) => mdiclink_reg(7), mdiclink_reg(6) => 
        mdiclink_reg(6), mdiclink_reg(5) => mdiclink_reg(5), 
        mdiclink_reg(4) => mdiclink_reg(4), mdiclink_reg(3) => 
        mdiclink_reg(3), mdiclink_reg(2) => mdiclink_reg(2), 
        mdiclink_reg(1) => mdiclink_reg(1), mdiclink_reg(0) => 
        mdiclink_reg(0), b11_OFWNT9L_8tZ(167) => 
        b11_OFWNT9L_8tZ(167), b11_OFWNT9L_8tZ(166) => 
        b11_OFWNT9L_8tZ(166), b11_OFWNT9L_8tZ(165) => 
        b11_OFWNT9L_8tZ(165), b11_OFWNT9L_8tZ(164) => 
        b11_OFWNT9L_8tZ(164), b11_OFWNT9L_8tZ(163) => 
        b11_OFWNT9L_8tZ(163), b11_OFWNT9L_8tZ(162) => 
        b11_OFWNT9L_8tZ(162), b11_OFWNT9L_8tZ(161) => 
        b11_OFWNT9L_8tZ(161), b11_OFWNT9L_8tZ(160) => 
        b11_OFWNT9L_8tZ(160), b11_OFWNT9L_8tZ(159) => 
        b11_OFWNT9L_8tZ(159), b11_OFWNT9L_8tZ(158) => 
        b11_OFWNT9L_8tZ(158), b11_OFWNT9L_8tZ(157) => 
        b11_OFWNT9L_8tZ(157), b11_OFWNT9L_8tZ(156) => 
        b11_OFWNT9L_8tZ(156), b11_OFWNT9L_8tZ(155) => 
        b11_OFWNT9L_8tZ(155), b11_OFWNT9L_8tZ(154) => 
        b11_OFWNT9L_8tZ(154), b11_OFWNT9L_8tZ(153) => 
        b11_OFWNT9L_8tZ(153), b11_OFWNT9L_8tZ(152) => 
        b11_OFWNT9L_8tZ(152), b11_OFWNT9L_8tZ(151) => 
        b11_OFWNT9L_8tZ(151), b11_OFWNT9L_8tZ(150) => 
        b11_OFWNT9L_8tZ(150), b11_OFWNT9L_8tZ(149) => 
        b11_OFWNT9L_8tZ(149), b11_OFWNT9L_8tZ(148) => 
        b11_OFWNT9L_8tZ(148), b11_OFWNT9L_8tZ(147) => 
        b11_OFWNT9L_8tZ(147), b11_OFWNT9L_8tZ(146) => 
        b11_OFWNT9L_8tZ(146), b11_OFWNT9L_8tZ(145) => 
        b11_OFWNT9L_8tZ(145), b11_OFWNT9L_8tZ(144) => 
        b11_OFWNT9L_8tZ(144), b11_OFWNT9L_8tZ(143) => 
        b11_OFWNT9L_8tZ(143), b11_OFWNT9L_8tZ(142) => 
        b11_OFWNT9L_8tZ(142), b11_OFWNT9L_8tZ(141) => 
        b11_OFWNT9L_8tZ(141), b11_OFWNT9L_8tZ(140) => 
        b11_OFWNT9L_8tZ(140), b11_OFWNT9L_8tZ(139) => 
        b11_OFWNT9L_8tZ(139), b11_OFWNT9L_8tZ(138) => 
        b11_OFWNT9L_8tZ(138), b11_OFWNT9L_8tZ(137) => 
        b11_OFWNT9L_8tZ(137), b11_OFWNT9L_8tZ(136) => 
        b11_OFWNT9L_8tZ(136), b11_OFWNT9L_8tZ(135) => 
        b11_OFWNT9L_8tZ(135), b11_OFWNT9L_8tZ(134) => 
        b11_OFWNT9L_8tZ(134), b11_OFWNT9L_8tZ(133) => 
        b11_OFWNT9L_8tZ(133), b11_OFWNT9L_8tZ(132) => 
        b11_OFWNT9L_8tZ(132), b11_OFWNT9L_8tZ(131) => 
        b11_OFWNT9L_8tZ(131), b11_OFWNT9L_8tZ(130) => 
        b11_OFWNT9L_8tZ(130), b11_OFWNT9L_8tZ(129) => 
        b11_OFWNT9L_8tZ(129), b11_OFWNT9L_8tZ(128) => 
        b11_OFWNT9L_8tZ(128), b11_OFWNT9L_8tZ(127) => 
        b11_OFWNT9L_8tZ(127), b11_OFWNT9L_8tZ(126) => 
        b11_OFWNT9L_8tZ(126), b11_OFWNT9L_8tZ(125) => 
        b11_OFWNT9L_8tZ(125), b11_OFWNT9L_8tZ(124) => 
        b11_OFWNT9L_8tZ(124), b11_OFWNT9L_8tZ(123) => 
        b11_OFWNT9L_8tZ(123), b11_OFWNT9L_8tZ(122) => 
        b11_OFWNT9L_8tZ(122), b11_OFWNT9L_8tZ(121) => 
        b11_OFWNT9L_8tZ(121), b11_OFWNT9L_8tZ(120) => 
        b11_OFWNT9L_8tZ(120), b11_OFWNT9L_8tZ(119) => 
        b11_OFWNT9L_8tZ(119), b11_OFWNT9L_8tZ(118) => 
        b11_OFWNT9L_8tZ(118), b11_OFWNT9L_8tZ(117) => 
        b11_OFWNT9L_8tZ(117), b11_OFWNT9L_8tZ(116) => 
        b11_OFWNT9L_8tZ(116), b11_OFWNT9L_8tZ(115) => 
        b11_OFWNT9L_8tZ(115), b11_OFWNT9L_8tZ(114) => 
        b11_OFWNT9L_8tZ(114), b11_OFWNT9L_8tZ(113) => 
        b11_OFWNT9L_8tZ(113), b11_OFWNT9L_8tZ(112) => 
        b11_OFWNT9L_8tZ(112), b11_OFWNT9L_8tZ(111) => 
        b11_OFWNT9L_8tZ(111), b11_OFWNT9L_8tZ(110) => 
        b11_OFWNT9L_8tZ(110), b11_OFWNT9L_8tZ(109) => 
        b11_OFWNT9L_8tZ(109), b11_OFWNT9L_8tZ(108) => 
        b11_OFWNT9L_8tZ(108), b11_OFWNT9L_8tZ(107) => 
        b11_OFWNT9L_8tZ(107), b11_OFWNT9L_8tZ(106) => 
        b11_OFWNT9L_8tZ(106), b11_OFWNT9L_8tZ(105) => 
        b11_OFWNT9L_8tZ(105), b11_OFWNT9L_8tZ(104) => 
        b11_OFWNT9L_8tZ(104), b11_OFWNT9L_8tZ(103) => 
        b11_OFWNT9L_8tZ(103), b11_OFWNT9L_8tZ(102) => 
        b11_OFWNT9L_8tZ(102), b11_OFWNT9L_8tZ(101) => 
        b11_OFWNT9L_8tZ(101), b11_OFWNT9L_8tZ(100) => 
        b11_OFWNT9L_8tZ(100), b11_OFWNT9L_8tZ(99) => 
        b11_OFWNT9L_8tZ(99), b11_OFWNT9L_8tZ(98) => 
        b11_OFWNT9L_8tZ(98), b11_OFWNT9L_8tZ(97) => 
        b11_OFWNT9L_8tZ(97), b11_OFWNT9L_8tZ(96) => 
        b11_OFWNT9L_8tZ(96), b11_OFWNT9L_8tZ(95) => 
        b11_OFWNT9L_8tZ(95), b11_OFWNT9L_8tZ(94) => 
        b11_OFWNT9L_8tZ(94), b11_OFWNT9L_8tZ(93) => 
        b11_OFWNT9L_8tZ(93), b11_OFWNT9L_8tZ(92) => 
        b11_OFWNT9L_8tZ(92), b11_OFWNT9L_8tZ(91) => 
        b11_OFWNT9L_8tZ(91), b11_OFWNT9L_8tZ(90) => 
        b11_OFWNT9L_8tZ(90), b11_OFWNT9L_8tZ(89) => 
        b11_OFWNT9L_8tZ(89), b11_OFWNT9L_8tZ(88) => 
        b11_OFWNT9L_8tZ(88), b11_OFWNT9L_8tZ(87) => 
        b11_OFWNT9L_8tZ(87), b11_OFWNT9L_8tZ(86) => 
        b11_OFWNT9L_8tZ(86), b11_OFWNT9L_8tZ(85) => 
        b11_OFWNT9L_8tZ(85), b11_OFWNT9L_8tZ(84) => 
        b11_OFWNT9L_8tZ(84), b11_OFWNT9L_8tZ(83) => 
        b11_OFWNT9L_8tZ(83), b11_OFWNT9L_8tZ(82) => 
        b11_OFWNT9L_8tZ(82), b11_OFWNT9L_8tZ(81) => 
        b11_OFWNT9L_8tZ(81), b11_OFWNT9L_8tZ(80) => 
        b11_OFWNT9L_8tZ(80), b11_OFWNT9L_8tZ(79) => 
        b11_OFWNT9L_8tZ(79), b11_OFWNT9L_8tZ(78) => 
        b11_OFWNT9L_8tZ(78), b11_OFWNT9L_8tZ(77) => 
        b11_OFWNT9L_8tZ(77), b11_OFWNT9L_8tZ(76) => 
        b11_OFWNT9L_8tZ(76), b11_OFWNT9L_8tZ(75) => 
        b11_OFWNT9L_8tZ(75), b11_OFWNT9L_8tZ(74) => 
        b11_OFWNT9L_8tZ(74), b11_OFWNT9L_8tZ(73) => 
        b11_OFWNT9L_8tZ(73), b11_OFWNT9L_8tZ(72) => 
        b11_OFWNT9L_8tZ(72), b11_OFWNT9L_8tZ(71) => 
        b11_OFWNT9L_8tZ(71), b11_OFWNT9L_8tZ(70) => 
        b11_OFWNT9L_8tZ(70), b11_OFWNT9L_8tZ(69) => 
        b11_OFWNT9L_8tZ(69), b11_OFWNT9L_8tZ(68) => 
        b11_OFWNT9L_8tZ(68), b11_OFWNT9L_8tZ(67) => 
        b11_OFWNT9L_8tZ(67), b11_OFWNT9L_8tZ(66) => 
        b11_OFWNT9L_8tZ(66), b11_OFWNT9L_8tZ(65) => 
        b11_OFWNT9L_8tZ(65), b11_OFWNT9L_8tZ(64) => 
        b11_OFWNT9L_8tZ(64), b11_OFWNT9L_8tZ(63) => 
        b11_OFWNT9L_8tZ(63), b11_OFWNT9L_8tZ(62) => 
        b11_OFWNT9L_8tZ(62), b11_OFWNT9L_8tZ(61) => 
        b11_OFWNT9L_8tZ(61), b11_OFWNT9L_8tZ(60) => 
        b11_OFWNT9L_8tZ(60), b11_OFWNT9L_8tZ(59) => 
        b11_OFWNT9L_8tZ(59), b11_OFWNT9L_8tZ(58) => 
        b11_OFWNT9L_8tZ(58), b11_OFWNT9L_8tZ(57) => 
        b11_OFWNT9L_8tZ(57), b11_OFWNT9L_8tZ(56) => 
        b11_OFWNT9L_8tZ(56), b11_OFWNT9L_8tZ(55) => 
        b11_OFWNT9L_8tZ(55), b11_OFWNT9L_8tZ(54) => 
        b11_OFWNT9L_8tZ(54), b11_OFWNT9L_8tZ(53) => 
        b11_OFWNT9L_8tZ(53), b11_OFWNT9L_8tZ(52) => 
        b11_OFWNT9L_8tZ(52), b11_OFWNT9L_8tZ(51) => 
        b11_OFWNT9L_8tZ(51), b11_OFWNT9L_8tZ(50) => 
        b11_OFWNT9L_8tZ(50), b11_OFWNT9L_8tZ(49) => 
        b11_OFWNT9L_8tZ(49), b11_OFWNT9L_8tZ(48) => 
        b11_OFWNT9L_8tZ(48), b11_OFWNT9L_8tZ(47) => 
        b11_OFWNT9L_8tZ(47), b11_OFWNT9L_8tZ(46) => 
        b11_OFWNT9L_8tZ(46), b11_OFWNT9L_8tZ(45) => 
        b11_OFWNT9L_8tZ(45), b11_OFWNT9L_8tZ(44) => 
        b11_OFWNT9L_8tZ(44), b11_OFWNT9L_8tZ(43) => 
        b11_OFWNT9L_8tZ(43), b11_OFWNT9L_8tZ(42) => 
        b11_OFWNT9L_8tZ(42), b11_OFWNT9L_8tZ(41) => 
        b11_OFWNT9L_8tZ(41), b11_OFWNT9L_8tZ(40) => 
        b11_OFWNT9L_8tZ(40), b11_OFWNT9L_8tZ(39) => 
        b11_OFWNT9L_8tZ(39), b11_OFWNT9L_8tZ(38) => 
        b11_OFWNT9L_8tZ(38), b11_OFWNT9L_8tZ(37) => 
        b11_OFWNT9L_8tZ(37), b11_OFWNT9L_8tZ(36) => 
        b11_OFWNT9L_8tZ(36), b11_OFWNT9L_8tZ(35) => 
        b11_OFWNT9L_8tZ(35), b11_OFWNT9L_8tZ(34) => 
        b11_OFWNT9L_8tZ(34), b11_OFWNT9L_8tZ(33) => 
        b11_OFWNT9L_8tZ(33), b11_OFWNT9L_8tZ(32) => 
        b11_OFWNT9L_8tZ(32), b11_OFWNT9L_8tZ(31) => 
        b11_OFWNT9L_8tZ(31), b11_OFWNT9L_8tZ(30) => 
        b11_OFWNT9L_8tZ(30), b11_OFWNT9L_8tZ(29) => 
        b11_OFWNT9L_8tZ(29), b11_OFWNT9L_8tZ(28) => 
        b11_OFWNT9L_8tZ(28), b11_OFWNT9L_8tZ(27) => 
        b11_OFWNT9L_8tZ(27), b11_OFWNT9L_8tZ(26) => 
        b11_OFWNT9L_8tZ(26), b11_OFWNT9L_8tZ(25) => 
        b11_OFWNT9L_8tZ(25), b11_OFWNT9L_8tZ(24) => 
        b11_OFWNT9L_8tZ(24), b11_OFWNT9L_8tZ(23) => 
        b11_OFWNT9L_8tZ(23), b11_OFWNT9L_8tZ(22) => 
        b11_OFWNT9L_8tZ(22), b11_OFWNT9L_8tZ(21) => 
        b11_OFWNT9L_8tZ(21), b11_OFWNT9L_8tZ(20) => 
        b11_OFWNT9L_8tZ(20), b11_OFWNT9L_8tZ(19) => 
        b11_OFWNT9L_8tZ(19), b11_OFWNT9L_8tZ(18) => 
        b11_OFWNT9L_8tZ(18), b11_OFWNT9L_8tZ(17) => 
        b11_OFWNT9L_8tZ(17), b11_OFWNT9L_8tZ(16) => 
        b11_OFWNT9L_8tZ(16), b11_OFWNT9L_8tZ(15) => 
        b11_OFWNT9L_8tZ(15), b11_OFWNT9L_8tZ(14) => 
        b11_OFWNT9L_8tZ(14), b11_OFWNT9L_8tZ(13) => 
        b11_OFWNT9L_8tZ(13), b11_OFWNT9L_8tZ(12) => 
        b11_OFWNT9L_8tZ(12), b11_OFWNT9L_8tZ(11) => 
        b11_OFWNT9L_8tZ(11), b11_OFWNT9L_8tZ(10) => 
        b11_OFWNT9L_8tZ(10), b11_OFWNT9L_8tZ(9) => 
        b11_OFWNT9L_8tZ(9), b11_OFWNT9L_8tZ(8) => 
        b11_OFWNT9L_8tZ(8), b11_OFWNT9L_8tZ(7) => 
        b11_OFWNT9L_8tZ(7), b11_OFWNT9L_8tZ(6) => 
        b11_OFWNT9L_8tZ(6), b11_OFWNT9L_8tZ(5) => 
        b11_OFWNT9L_8tZ(5), b11_OFWNT9L_8tZ(4) => 
        b11_OFWNT9L_8tZ(4), b11_OFWNT9L_8tZ(3) => 
        b11_OFWNT9L_8tZ(3), b11_OFWNT9L_8tZ(2) => 
        b11_OFWNT9L_8tZ(2), b11_OFWNT9L_8tZ(1) => 
        b11_OFWNT9L_8tZ(1), b11_OFWNT9L_8tZ(0) => 
        b11_OFWNT9L_8tZ(0), b4_nUAi(502) => \b4_nUAi[502]\, 
        b4_nUAi(501) => \b4_nUAi[501]\, b4_nUAi(500) => 
        \b4_nUAi[500]\, b4_nUAi(499) => \b4_nUAi[499]\, 
        b4_nUAi(498) => \b4_nUAi[498]\, b4_nUAi(497) => 
        \b4_nUAi[497]\, b4_nUAi(496) => \b4_nUAi[496]\, 
        b4_nUAi(495) => \b4_nUAi[495]\, b4_nUAi(494) => 
        \b4_nUAi[494]\, b4_nUAi(493) => \b4_nUAi[493]\, 
        b4_nUAi(492) => \b4_nUAi[492]\, b4_nUAi(491) => 
        \b4_nUAi[491]\, b4_nUAi(490) => \b4_nUAi[490]\, 
        b4_nUAi(489) => \b4_nUAi[489]\, b4_nUAi(488) => 
        \b4_nUAi[488]\, b4_nUAi(487) => \b4_nUAi[487]\, 
        b4_nUAi(486) => \b4_nUAi[486]\, b4_nUAi(485) => 
        \b4_nUAi[485]\, b4_nUAi(484) => \b4_nUAi[484]\, 
        b4_nUAi(483) => \b4_nUAi[483]\, b4_nUAi(482) => 
        \b4_nUAi[482]\, b4_nUAi(481) => \b4_nUAi[481]\, 
        b4_nUAi(480) => \b4_nUAi[480]\, b4_nUAi(479) => 
        \b4_nUAi[479]\, b4_nUAi(478) => \b4_nUAi[478]\, 
        b4_nUAi(477) => \b4_nUAi[477]\, b4_nUAi(476) => 
        \b4_nUAi[476]\, b4_nUAi(475) => \b4_nUAi[475]\, 
        b4_nUAi(474) => \b4_nUAi[474]\, b4_nUAi(473) => 
        \b4_nUAi[473]\, b4_nUAi(472) => \b4_nUAi[472]\, 
        b4_nUAi(471) => \b4_nUAi[471]\, b4_nUAi(470) => 
        \b4_nUAi[470]\, b4_nUAi(469) => \b4_nUAi[469]\, 
        b4_nUAi(468) => \b4_nUAi[468]\, b4_nUAi(467) => 
        \b4_nUAi[467]\, b4_nUAi(466) => \b4_nUAi[466]\, 
        b4_nUAi(465) => \b4_nUAi[465]\, b4_nUAi(464) => 
        \b4_nUAi[464]\, b4_nUAi(463) => \b4_nUAi[463]\, 
        b4_nUAi(462) => \b4_nUAi[462]\, b4_nUAi(461) => 
        \b4_nUAi[461]\, b4_nUAi(460) => \b4_nUAi[460]\, 
        b4_nUAi(459) => \b4_nUAi[459]\, b4_nUAi(458) => 
        \b4_nUAi[458]\, b4_nUAi(457) => \b4_nUAi[457]\, 
        b4_nUAi(456) => \b4_nUAi[456]\, b4_nUAi(455) => 
        \b4_nUAi[455]\, b4_nUAi(454) => \b4_nUAi[454]\, 
        b4_nUAi(453) => \b4_nUAi[453]\, b4_nUAi(452) => 
        \b4_nUAi[452]\, b4_nUAi(451) => \b4_nUAi[451]\, 
        b4_nUAi(450) => \b4_nUAi[450]\, b4_nUAi(449) => 
        \b4_nUAi[449]\, b4_nUAi(448) => \b4_nUAi[448]\, 
        b4_nUAi(447) => \b4_nUAi[447]\, b4_nUAi(446) => 
        \b4_nUAi[446]\, b4_nUAi(445) => \b4_nUAi[445]\, 
        b4_nUAi(444) => \b4_nUAi[444]\, b4_nUAi(443) => 
        \b4_nUAi[443]\, b4_nUAi(442) => \b4_nUAi[442]\, 
        b4_nUAi(441) => \b4_nUAi[441]\, b4_nUAi(440) => 
        \b4_nUAi[440]\, b4_nUAi(439) => \b4_nUAi[439]\, 
        b4_nUAi(438) => \b4_nUAi[438]\, b4_nUAi(437) => 
        \b4_nUAi[437]\, b4_nUAi(436) => \b4_nUAi[436]\, 
        b4_nUAi(435) => \b4_nUAi[435]\, b4_nUAi(434) => 
        \b4_nUAi[434]\, b4_nUAi(433) => \b4_nUAi[433]\, 
        b4_nUAi(432) => \b4_nUAi[432]\, b4_nUAi(431) => 
        \b4_nUAi[431]\, b4_nUAi(430) => \b4_nUAi[430]\, 
        b4_nUAi(429) => \b4_nUAi[429]\, b4_nUAi(428) => 
        \b4_nUAi[428]\, b4_nUAi(427) => \b4_nUAi[427]\, 
        b4_nUAi(426) => \b4_nUAi[426]\, b4_nUAi(425) => 
        \b4_nUAi[425]\, b4_nUAi(424) => \b4_nUAi[424]\, 
        b4_nUAi(423) => \b4_nUAi[423]\, b4_nUAi(422) => 
        \b4_nUAi[422]\, b4_nUAi(421) => \b4_nUAi[421]\, 
        b4_nUAi(420) => \b4_nUAi[420]\, b4_nUAi(419) => 
        \b4_nUAi[419]\, b4_nUAi(418) => \b4_nUAi[418]\, 
        b4_nUAi(417) => \b4_nUAi[417]\, b4_nUAi(416) => 
        \b4_nUAi[416]\, b4_nUAi(415) => \b4_nUAi[415]\, 
        b4_nUAi(414) => \b4_nUAi[414]\, b4_nUAi(413) => 
        \b4_nUAi[413]\, b4_nUAi(412) => \b4_nUAi[412]\, 
        b4_nUAi(411) => \b4_nUAi[411]\, b4_nUAi(410) => 
        \b4_nUAi[410]\, b4_nUAi(409) => \b4_nUAi[409]\, 
        b4_nUAi(408) => \b4_nUAi[408]\, b4_nUAi(407) => 
        \b4_nUAi[407]\, b4_nUAi(406) => \b4_nUAi[406]\, 
        b4_nUAi(405) => \b4_nUAi[405]\, b4_nUAi(404) => 
        \b4_nUAi[404]\, b4_nUAi(403) => \b4_nUAi[403]\, 
        b4_nUAi(402) => \b4_nUAi[402]\, b4_nUAi(401) => 
        \b4_nUAi[401]\, b4_nUAi(400) => \b4_nUAi[400]\, 
        b4_nUAi(399) => \b4_nUAi[399]\, b4_nUAi(398) => 
        \b4_nUAi[398]\, b4_nUAi(397) => \b4_nUAi[397]\, 
        b4_nUAi(396) => \b4_nUAi[396]\, b4_nUAi(395) => 
        \b4_nUAi[395]\, b4_nUAi(394) => \b4_nUAi[394]\, 
        b4_nUAi(393) => \b4_nUAi[393]\, b4_nUAi(392) => 
        \b4_nUAi[392]\, b4_nUAi(391) => \b4_nUAi[391]\, 
        b4_nUAi(390) => \b4_nUAi[390]\, b4_nUAi(389) => 
        \b4_nUAi[389]\, b4_nUAi(388) => \b4_nUAi[388]\, 
        b4_nUAi(387) => \b4_nUAi[387]\, b4_nUAi(386) => 
        \b4_nUAi[386]\, b4_nUAi(385) => \b4_nUAi[385]\, 
        b4_nUAi(384) => \b4_nUAi[384]\, b4_nUAi(383) => 
        \b4_nUAi[383]\, b4_nUAi(382) => \b4_nUAi[382]\, 
        b4_nUAi(381) => \b4_nUAi[381]\, b4_nUAi(380) => 
        \b4_nUAi[380]\, b4_nUAi(379) => \b4_nUAi[379]\, 
        b4_nUAi(378) => \b4_nUAi[378]\, b4_nUAi(377) => 
        \b4_nUAi[377]\, b4_nUAi(376) => \b4_nUAi[376]\, 
        b4_nUAi(375) => \b4_nUAi[375]\, b4_nUAi(374) => 
        \b4_nUAi[374]\, b4_nUAi(373) => \b4_nUAi[373]\, 
        b4_nUAi(372) => \b4_nUAi[372]\, b4_nUAi(371) => 
        \b4_nUAi[371]\, b4_nUAi(370) => \b4_nUAi[370]\, 
        b4_nUAi(369) => \b4_nUAi[369]\, b4_nUAi(368) => 
        \b4_nUAi[368]\, b4_nUAi(367) => \b4_nUAi[367]\, 
        b4_nUAi(366) => \b4_nUAi[366]\, b4_nUAi(365) => 
        \b4_nUAi[365]\, b4_nUAi(364) => \b4_nUAi[364]\, 
        b4_nUAi(363) => \b4_nUAi[363]\, b4_nUAi(362) => 
        \b4_nUAi[362]\, b4_nUAi(361) => \b4_nUAi[361]\, 
        b4_nUAi(360) => \b4_nUAi[360]\, b4_nUAi(359) => 
        \b4_nUAi[359]\, b4_nUAi(358) => \b4_nUAi[358]\, 
        b4_nUAi(357) => \b4_nUAi[357]\, b4_nUAi(356) => 
        \b4_nUAi[356]\, b4_nUAi(355) => \b4_nUAi[355]\, 
        b4_nUAi(354) => \b4_nUAi[354]\, b4_nUAi(353) => 
        \b4_nUAi[353]\, b4_nUAi(352) => \b4_nUAi[352]\, 
        b4_nUAi(351) => \b4_nUAi[351]\, b4_nUAi(350) => 
        \b4_nUAi[350]\, b4_nUAi(349) => \b4_nUAi[349]\, 
        b4_nUAi(348) => \b4_nUAi[348]\, b4_nUAi(347) => 
        \b4_nUAi[347]\, b4_nUAi(346) => \b4_nUAi[346]\, 
        b4_nUAi(345) => \b4_nUAi[345]\, b4_nUAi(344) => 
        \b4_nUAi[344]\, b4_nUAi(343) => \b4_nUAi[343]\, 
        b4_nUAi(342) => \b4_nUAi[342]\, b4_nUAi(341) => 
        \b4_nUAi[341]\, b4_nUAi(340) => \b4_nUAi[340]\, 
        b4_nUAi(339) => \b4_nUAi[339]\, b4_nUAi(338) => 
        \b4_nUAi[338]\, b4_nUAi(337) => \b4_nUAi[337]\, 
        b4_nUAi(336) => \b4_nUAi[336]\, b4_nUAi(335) => 
        \b4_nUAi[335]\, b4_nUAi(334) => \b4_nUAi[334]\, 
        b4_nUAi(333) => \b4_nUAi[333]\, b4_nUAi(332) => 
        \b4_nUAi[332]\, b4_nUAi(331) => \b4_nUAi[331]\, 
        b4_nUAi(330) => \b4_nUAi[330]\, b4_nUAi(329) => 
        \b4_nUAi[329]\, b4_nUAi(328) => \b4_nUAi[328]\, 
        b4_nUAi(327) => \b4_nUAi[327]\, b4_nUAi(326) => 
        \b4_nUAi[326]\, b4_nUAi(325) => \b4_nUAi[325]\, 
        b4_nUAi(324) => \b4_nUAi[324]\, b4_nUAi(323) => 
        \b4_nUAi[323]\, b4_nUAi(322) => \b4_nUAi[322]\, 
        b4_nUAi(321) => \b4_nUAi[321]\, b4_nUAi(320) => 
        \b4_nUAi[320]\, b4_nUAi(319) => \b4_nUAi[319]\, 
        b4_nUAi(318) => \b4_nUAi[318]\, b4_nUAi(317) => 
        \b4_nUAi[317]\, b4_nUAi(316) => \b4_nUAi[316]\, 
        b4_nUAi(315) => \b4_nUAi[315]\, b4_nUAi(314) => 
        \b4_nUAi[314]\, b4_nUAi(313) => \b4_nUAi[313]\, 
        b4_nUAi(312) => \b4_nUAi[312]\, b4_nUAi(311) => 
        \b4_nUAi[311]\, b4_nUAi(310) => \b4_nUAi[310]\, 
        b4_nUAi(309) => \b4_nUAi[309]\, b4_nUAi(308) => 
        \b4_nUAi[308]\, b4_nUAi(307) => \b4_nUAi[307]\, 
        b4_nUAi(306) => \b4_nUAi[306]\, b4_nUAi(305) => 
        \b4_nUAi[305]\, b4_nUAi(304) => \b4_nUAi[304]\, 
        b4_nUAi(303) => \b4_nUAi[303]\, b4_nUAi(302) => 
        \b4_nUAi[302]\, b4_nUAi(301) => \b4_nUAi[301]\, 
        b4_nUAi(300) => \b4_nUAi[300]\, b4_nUAi(299) => 
        \b4_nUAi[299]\, b4_nUAi(298) => \b4_nUAi[298]\, 
        b4_nUAi(297) => \b4_nUAi[297]\, b4_nUAi(296) => 
        \b4_nUAi[296]\, b4_nUAi(295) => \b4_nUAi[295]\, 
        b4_nUAi(294) => \b4_nUAi[294]\, b4_nUAi(293) => 
        \b4_nUAi[293]\, b4_nUAi(292) => \b4_nUAi[292]\, 
        b4_nUAi(291) => \b4_nUAi[291]\, b4_nUAi(290) => 
        \b4_nUAi[290]\, b4_nUAi(289) => \b4_nUAi[289]\, 
        b4_nUAi(288) => \b4_nUAi[288]\, b4_nUAi(287) => 
        \b4_nUAi[287]\, b4_nUAi(286) => \b4_nUAi[286]\, 
        b4_nUAi(285) => \b4_nUAi[285]\, b4_nUAi(284) => 
        \b4_nUAi[284]\, b4_nUAi(283) => \b4_nUAi[283]\, 
        b4_nUAi(282) => \b4_nUAi[282]\, b4_nUAi(281) => 
        \b4_nUAi[281]\, b4_nUAi(280) => \b4_nUAi[280]\, 
        b4_nUAi(279) => \b4_nUAi[279]\, b4_nUAi(278) => 
        \b4_nUAi[278]\, b4_nUAi(277) => \b4_nUAi[277]\, 
        b4_nUAi(276) => \b4_nUAi[276]\, b4_nUAi(275) => 
        \b4_nUAi[275]\, b4_nUAi(274) => \b4_nUAi[274]\, 
        b4_nUAi(273) => \b4_nUAi[273]\, b4_nUAi(272) => 
        \b4_nUAi[272]\, b4_nUAi(271) => \b4_nUAi[271]\, 
        b4_nUAi(270) => \b4_nUAi[270]\, b4_nUAi(269) => 
        \b4_nUAi[269]\, b4_nUAi(268) => \b4_nUAi[268]\, 
        b4_nUAi(267) => \b4_nUAi[267]\, b4_nUAi(266) => 
        \b4_nUAi[266]\, b4_nUAi(265) => \b4_nUAi[265]\, 
        b4_nUAi(264) => \b4_nUAi[264]\, b4_nUAi(263) => 
        \b4_nUAi[263]\, b4_nUAi(262) => \b4_nUAi[262]\, 
        b4_nUAi(261) => \b4_nUAi[261]\, b4_nUAi(260) => 
        \b4_nUAi[260]\, b4_nUAi(259) => \b4_nUAi[259]\, 
        b4_nUAi(258) => \b4_nUAi[258]\, b4_nUAi(257) => 
        \b4_nUAi[257]\, b4_nUAi(256) => \b4_nUAi[256]\, 
        b4_nUAi(255) => \b4_nUAi[255]\, b4_nUAi(254) => 
        \b4_nUAi[254]\, b4_nUAi(253) => \b4_nUAi[253]\, 
        b4_nUAi(252) => \b4_nUAi[252]\, b4_nUAi(251) => 
        \b4_nUAi[251]\, b4_nUAi(250) => \b4_nUAi[250]\, 
        b4_nUAi(249) => \b4_nUAi[249]\, b4_nUAi(248) => 
        \b4_nUAi[248]\, b4_nUAi(247) => \b4_nUAi[247]\, 
        b4_nUAi(246) => \b4_nUAi[246]\, b4_nUAi(245) => 
        \b4_nUAi[245]\, b4_nUAi(244) => \b4_nUAi[244]\, 
        b4_nUAi(243) => \b4_nUAi[243]\, b4_nUAi(242) => 
        \b4_nUAi[242]\, b4_nUAi(241) => \b4_nUAi[241]\, 
        b4_nUAi(240) => \b4_nUAi[240]\, b4_nUAi(239) => 
        \b4_nUAi[239]\, b4_nUAi(238) => \b4_nUAi[238]\, 
        b4_nUAi(237) => \b4_nUAi[237]\, b4_nUAi(236) => 
        \b4_nUAi[236]\, b4_nUAi(235) => \b4_nUAi[235]\, 
        b4_nUAi(234) => \b4_nUAi[234]\, b4_nUAi(233) => 
        \b4_nUAi[233]\, b4_nUAi(232) => \b4_nUAi[232]\, 
        b4_nUAi(231) => \b4_nUAi[231]\, b4_nUAi(230) => 
        \b4_nUAi[230]\, b4_nUAi(229) => \b4_nUAi[229]\, 
        b4_nUAi(228) => \b4_nUAi[228]\, b4_nUAi(227) => 
        \b4_nUAi[227]\, b4_nUAi(226) => \b4_nUAi[226]\, 
        b4_nUAi(225) => \b4_nUAi[225]\, b4_nUAi(224) => 
        \b4_nUAi[224]\, b4_nUAi(223) => \b4_nUAi[223]\, 
        b4_nUAi(222) => \b4_nUAi[222]\, b4_nUAi(221) => 
        \b4_nUAi[221]\, b4_nUAi(220) => \b4_nUAi[220]\, 
        b4_nUAi(219) => \b4_nUAi[219]\, b4_nUAi(218) => 
        \b4_nUAi[218]\, b4_nUAi(217) => \b4_nUAi[217]\, 
        b4_nUAi(216) => \b4_nUAi[216]\, b4_nUAi(215) => 
        \b4_nUAi[215]\, b4_nUAi(214) => \b4_nUAi[214]\, 
        b4_nUAi(213) => \b4_nUAi[213]\, b4_nUAi(212) => 
        \b4_nUAi[212]\, b4_nUAi(211) => \b4_nUAi[211]\, 
        b4_nUAi(210) => \b4_nUAi[210]\, b4_nUAi(209) => 
        \b4_nUAi[209]\, b4_nUAi(208) => \b4_nUAi[208]\, 
        b4_nUAi(207) => \b4_nUAi[207]\, b4_nUAi(206) => 
        \b4_nUAi[206]\, b4_nUAi(205) => \b4_nUAi[205]\, 
        b4_nUAi(204) => \b4_nUAi[204]\, b4_nUAi(203) => 
        \b4_nUAi[203]\, b4_nUAi(202) => \b4_nUAi[202]\, 
        b4_nUAi(201) => \b4_nUAi[201]\, b4_nUAi(200) => 
        \b4_nUAi[200]\, b4_nUAi(199) => \b4_nUAi[199]\, 
        b4_nUAi(198) => \b4_nUAi[198]\, b4_nUAi(197) => 
        \b4_nUAi[197]\, b4_nUAi(196) => \b4_nUAi[196]\, 
        b4_nUAi(195) => \b4_nUAi[195]\, b4_nUAi(194) => 
        \b4_nUAi[194]\, b4_nUAi(193) => \b4_nUAi[193]\, 
        b4_nUAi(192) => \b4_nUAi[192]\, b4_nUAi(191) => 
        \b4_nUAi[191]\, b4_nUAi(190) => \b4_nUAi[190]\, 
        b4_nUAi(189) => \b4_nUAi[189]\, b4_nUAi(188) => 
        \b4_nUAi[188]\, b4_nUAi(187) => \b4_nUAi[187]\, 
        b4_nUAi(186) => \b4_nUAi[186]\, b4_nUAi(185) => 
        \b4_nUAi[185]\, b4_nUAi(184) => \b4_nUAi[184]\, 
        b4_nUAi(183) => \b4_nUAi[183]\, b4_nUAi(182) => 
        \b4_nUAi[182]\, b4_nUAi(181) => \b4_nUAi[181]\, 
        b4_nUAi(180) => \b4_nUAi[180]\, b4_nUAi(179) => 
        \b4_nUAi[179]\, b4_nUAi(178) => \b4_nUAi[178]\, 
        b4_nUAi(177) => \b4_nUAi[177]\, b4_nUAi(176) => 
        \b4_nUAi[176]\, b4_nUAi(175) => \b4_nUAi[175]\, 
        b4_nUAi(174) => \b4_nUAi[174]\, b4_nUAi(173) => 
        \b4_nUAi[173]\, b4_nUAi(172) => \b4_nUAi[172]\, 
        b4_nUAi(171) => \b4_nUAi[171]\, b4_nUAi(170) => 
        \b4_nUAi[170]\, b4_nUAi(169) => \b4_nUAi[169]\, 
        b4_nUAi(168) => \b4_nUAi[168]\, b4_nUAi(167) => 
        \b4_nUAi[167]\, b4_nUAi(166) => \b4_nUAi[166]\, 
        b4_nUAi(165) => \b4_nUAi[165]\, b4_nUAi(164) => 
        \b4_nUAi[164]\, b4_nUAi(163) => \b4_nUAi[163]\, 
        b4_nUAi(162) => \b4_nUAi[162]\, b4_nUAi(161) => 
        \b4_nUAi[161]\, b4_nUAi(160) => \b4_nUAi[160]\, 
        b4_nUAi(159) => \b4_nUAi[159]\, b4_nUAi(158) => 
        \b4_nUAi[158]\, b4_nUAi(157) => \b4_nUAi[157]\, 
        b4_nUAi(156) => \b4_nUAi[156]\, b4_nUAi(155) => 
        \b4_nUAi[155]\, b4_nUAi(154) => \b4_nUAi[154]\, 
        b4_nUAi(153) => \b4_nUAi[153]\, b4_nUAi(152) => 
        \b4_nUAi[152]\, b4_nUAi(151) => \b4_nUAi[151]\, 
        b4_nUAi(150) => \b4_nUAi[150]\, b4_nUAi(149) => 
        \b4_nUAi[149]\, b4_nUAi(148) => \b4_nUAi[148]\, 
        b4_nUAi(147) => \b4_nUAi[147]\, b4_nUAi(146) => 
        \b4_nUAi[146]\, b4_nUAi(145) => \b4_nUAi[145]\, 
        b4_nUAi(144) => \b4_nUAi[144]\, b4_nUAi(143) => 
        \b4_nUAi[143]\, b4_nUAi(142) => \b4_nUAi[142]\, 
        b4_nUAi(141) => \b4_nUAi[141]\, b4_nUAi(140) => 
        \b4_nUAi[140]\, b4_nUAi(139) => \b4_nUAi[139]\, 
        b4_nUAi(138) => \b4_nUAi[138]\, b4_nUAi(137) => 
        \b4_nUAi[137]\, b4_nUAi(136) => \b4_nUAi[136]\, 
        b4_nUAi(135) => \b4_nUAi[135]\, b4_nUAi(134) => 
        \b4_nUAi[134]\, b4_nUAi(133) => \b4_nUAi[133]\, 
        b4_nUAi(132) => \b4_nUAi[132]\, b4_nUAi(131) => 
        \b4_nUAi[131]\, b4_nUAi(130) => \b4_nUAi[130]\, 
        b4_nUAi(129) => \b4_nUAi[129]\, b4_nUAi(128) => 
        \b4_nUAi[128]\, b4_nUAi(127) => \b4_nUAi[127]\, 
        b4_nUAi(126) => \b4_nUAi[126]\, b4_nUAi(125) => 
        \b4_nUAi[125]\, b4_nUAi(124) => \b4_nUAi[124]\, 
        b4_nUAi(123) => \b4_nUAi[123]\, b4_nUAi(122) => 
        \b4_nUAi[122]\, b4_nUAi(121) => \b4_nUAi[121]\, 
        b4_nUAi(120) => \b4_nUAi[120]\, b4_nUAi(119) => 
        \b4_nUAi[119]\, b4_nUAi(118) => \b4_nUAi[118]\, 
        b4_nUAi(117) => \b4_nUAi[117]\, b4_nUAi(116) => 
        \b4_nUAi[116]\, b4_nUAi(115) => \b4_nUAi[115]\, 
        b4_nUAi(114) => \b4_nUAi[114]\, b4_nUAi(113) => 
        \b4_nUAi[113]\, b4_nUAi(112) => \b4_nUAi[112]\, 
        b4_nUAi(111) => \b4_nUAi[111]\, b4_nUAi(110) => 
        \b4_nUAi[110]\, b4_nUAi(109) => \b4_nUAi[109]\, 
        b4_nUAi(108) => \b4_nUAi[108]\, b4_nUAi(107) => 
        \b4_nUAi[107]\, b4_nUAi(106) => \b4_nUAi[106]\, 
        b4_nUAi(105) => \b4_nUAi[105]\, b4_nUAi(104) => 
        \b4_nUAi[104]\, b4_nUAi(103) => \b4_nUAi[103]\, 
        b4_nUAi(102) => \b4_nUAi[102]\, b4_nUAi(101) => 
        \b4_nUAi[101]\, b4_nUAi(100) => \b4_nUAi[100]\, 
        b4_nUAi(99) => \b4_nUAi[99]\, b4_nUAi(98) => 
        \b4_nUAi[98]\, b4_nUAi(97) => \b4_nUAi[97]\, b4_nUAi(96)
         => \b4_nUAi[96]\, b4_nUAi(95) => \b4_nUAi[95]\, 
        b4_nUAi(94) => \b4_nUAi[94]\, b4_nUAi(93) => 
        \b4_nUAi[93]\, b4_nUAi(92) => \b4_nUAi[92]\, b4_nUAi(91)
         => \b4_nUAi[91]\, b4_nUAi(90) => \b4_nUAi[90]\, 
        b4_nUAi(89) => \b4_nUAi[89]\, b4_nUAi(88) => 
        \b4_nUAi[88]\, b4_nUAi(87) => \b4_nUAi[87]\, b4_nUAi(86)
         => \b4_nUAi[86]\, b4_nUAi(85) => \b4_nUAi[85]\, 
        b4_nUAi(84) => \b4_nUAi[84]\, b4_nUAi(83) => 
        \b4_nUAi[83]\, b4_nUAi(82) => \b4_nUAi[82]\, b4_nUAi(81)
         => \b4_nUAi[81]\, b4_nUAi(80) => \b4_nUAi[80]\, 
        b4_nUAi(79) => \b4_nUAi[79]\, b4_nUAi(78) => 
        \b4_nUAi[78]\, b4_nUAi(77) => \b4_nUAi[77]\, b4_nUAi(76)
         => \b4_nUAi[76]\, b4_nUAi(75) => \b4_nUAi[75]\, 
        b4_nUAi(74) => \b4_nUAi[74]\, b4_nUAi(73) => 
        \b4_nUAi[73]\, b4_nUAi(72) => \b4_nUAi[72]\, b4_nUAi(71)
         => \b4_nUAi[71]\, b4_nUAi(70) => \b4_nUAi[70]\, 
        b4_nUAi(69) => \b4_nUAi[69]\, b4_nUAi(68) => 
        \b4_nUAi[68]\, b4_nUAi(67) => \b4_nUAi[67]\, b4_nUAi(66)
         => \b4_nUAi[66]\, b4_nUAi(65) => \b4_nUAi[65]\, 
        b4_nUAi(64) => \b4_nUAi[64]\, b4_nUAi(63) => 
        \b4_nUAi[63]\, b4_nUAi(62) => \b4_nUAi[62]\, b4_nUAi(61)
         => \b4_nUAi[61]\, b4_nUAi(60) => \b4_nUAi[60]\, 
        b4_nUAi(59) => \b4_nUAi[59]\, b4_nUAi(58) => 
        \b4_nUAi[58]\, b4_nUAi(57) => \b4_nUAi[57]\, b4_nUAi(56)
         => \b4_nUAi[56]\, b4_nUAi(55) => \b4_nUAi[55]\, 
        b4_nUAi(54) => \b4_nUAi[54]\, b4_nUAi(53) => 
        \b4_nUAi[53]\, b4_nUAi(52) => \b4_nUAi[52]\, b4_nUAi(51)
         => \b4_nUAi[51]\, b4_nUAi(50) => \b4_nUAi[50]\, 
        b4_nUAi(49) => \b4_nUAi[49]\, b4_nUAi(48) => 
        \b4_nUAi[48]\, b4_nUAi(47) => \b4_nUAi[47]\, b4_nUAi(46)
         => \b4_nUAi[46]\, b4_nUAi(45) => \b4_nUAi[45]\, 
        b4_nUAi(44) => \b4_nUAi[44]\, b4_nUAi(43) => 
        \b4_nUAi[43]\, b4_nUAi(42) => \b4_nUAi[42]\, b4_nUAi(41)
         => \b4_nUAi[41]\, b4_nUAi(40) => \b4_nUAi[40]\, 
        b4_nUAi(39) => \b4_nUAi[39]\, b4_nUAi(38) => 
        \b4_nUAi[38]\, b4_nUAi(37) => \b4_nUAi[37]\, b4_nUAi(36)
         => \b4_nUAi[36]\, b4_nUAi(35) => \b4_nUAi[35]\, 
        b4_nUAi(34) => \b4_nUAi[34]\, b4_nUAi(33) => 
        \b4_nUAi[33]\, b4_nUAi(32) => \b4_nUAi[32]\, b4_nUAi(31)
         => \b4_nUAi[31]\, b4_nUAi(30) => \b4_nUAi[30]\, 
        b4_nUAi(29) => \b4_nUAi[29]\, b4_nUAi(28) => 
        \b4_nUAi[28]\, b4_nUAi(27) => \b4_nUAi[27]\, b4_nUAi(26)
         => \b4_nUAi[26]\, b4_nUAi(25) => \b4_nUAi[25]\, 
        b4_nUAi(24) => \b4_nUAi[24]\, b4_nUAi(23) => 
        \b4_nUAi[23]\, b4_nUAi(22) => \b4_nUAi[22]\, b4_nUAi(21)
         => \b4_nUAi[21]\, b4_nUAi(20) => \b4_nUAi[20]\, 
        b4_nUAi(19) => \b4_nUAi[19]\, b4_nUAi(18) => 
        \b4_nUAi[18]\, b4_nUAi(17) => \b4_nUAi[17]\, b4_nUAi(16)
         => \b4_nUAi[16]\, b4_nUAi(15) => \b4_nUAi[15]\, 
        b4_nUAi(14) => \b4_nUAi[14]\, b4_nUAi(13) => 
        \b4_nUAi[13]\, b4_nUAi(12) => \b4_nUAi[12]\, b4_nUAi(11)
         => \b4_nUAi[11]\, b4_nUAi(10) => \b4_nUAi[10]\, 
        b4_nUAi(9) => \b4_nUAi[9]\, b4_nUAi(8) => \b4_nUAi[8]\, 
        b4_nUAi(7) => \b4_nUAi[7]\, b4_nUAi(6) => \b4_nUAi[6]\, 
        b4_nUAi(5) => \b4_nUAi[5]\, b4_nUAi(4) => \b4_nUAi[4]\, 
        b4_nUAi(3) => \b4_nUAi[3]\, b4_nUAi(2) => \b4_nUAi[2]\, 
        b4_nUAi(1) => \b4_nUAi[1]\, b4_nUAi(0) => \b4_nUAi[0]\, 
        b10_nYBzIXrKbK_0 => b10_nYBzIXrKbK_0, CommsFPGA_CCC_0_GL0
         => CommsFPGA_CCC_0_GL0, b12_PSyi_XlK_qHv => 
        \b12_PSyi_XlK_qHv\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b8_nR_ymqrG_12s_5s_0_0s_0s_1_2046_x_0 is

    port( IICE_comm2iice  : in    std_logic_vector(11 downto 7);
          b6_nUT_IF       : out   std_logic_vector(11 downto 0);
          b6_nfs_IF       : out   std_logic_vector(4 downto 0);
          b6_nfs_IF_i_0   : out   std_logic;
          b9_vbTtJX_ab    : in    std_logic;
          b11_vABZ3qsY_qH : out   std_logic;
          b10_vbTtJX_Y2x  : out   std_logic;
          b10_PKFoLX_Y2x  : out   std_logic;
          b7_nUTQ_9u      : in    std_logic;
          b8_nUTQ_XlK     : out   std_logic;
          b9_PKFoLX_ab    : in    std_logic
        );

end b8_nR_ymqrG_12s_5s_0_0s_0s_1_2046_x_0;

architecture DEF_ARCH of b8_nR_ymqrG_12s_5s_0_0s_0s_1_2046_x_0 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \b6_nfs_IF[1]\, \b3_nfs[1]\, \b6_nfs_IF_i_0\, 
        \b10_nUT_M9kYfr[2]_net_1\, VCC_net_1, 
        \b10_nUT_M9kYfr[3]_net_1\, \b10_nUT_M9kYfr4\, GND_net_1, 
        \b10_nUT_M9kYfr[4]_net_1\, \b10_nUT_M9kYfr[5]_net_1\, 
        \b10_nUT_M9kYfr[6]_net_1\, \b10_nUT_M9kYfr[7]_net_1\, 
        \b10_nUT_M9kYfr[8]_net_1\, \b10_nUT_M9kYfr[9]_net_1\, 
        \b10_nUT_M9kYfr[10]_net_1\, \b10_nUT_M9kYfr[11]_net_1\, 
        \b8_nUTQ_XlK\, \b10_nfs_M9kYfr[1]_net_1\, 
        \b10_nfs_M9kYfr[2]_net_1\, \b10_nfs_M9kYfr[3]_net_1\, 
        \b10_nfs_M9kYfr[4]_net_1\, \b10_nfs_M9kYfr4\, 
        \b10_PKFoLX_Y2x\, \b10_nUT_M9kYfr[1]_net_1\, 
        \b10_vbTtJX_Y2x\, \b15_vABZ3qsY_ub3Rme3\ : std_logic;

begin 

    b6_nfs_IF(1) <= \b6_nfs_IF[1]\;
    b6_nfs_IF_i_0 <= \b6_nfs_IF_i_0\;
    b10_vbTtJX_Y2x <= \b10_vbTtJX_Y2x\;
    b10_PKFoLX_Y2x <= \b10_PKFoLX_Y2x\;
    b8_nUTQ_XlK <= \b8_nUTQ_XlK\;

    \genblk2.b3_nUT[10]\ : SLE
      port map(D => \b10_nUT_M9kYfr[10]_net_1\, CLK => 
        IICE_comm2iice(8), EN => b9_PKFoLX_ab, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => b6_nUT_IF(10));
    
    \genblk1.b3_nfs[4]\ : SLE
      port map(D => \b10_nfs_M9kYfr[4]_net_1\, CLK => 
        IICE_comm2iice(8), EN => b7_nUTQ_9u, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => b6_nfs_IF(4));
    
    \b10_nUT_M9kYfr[6]\ : SLE
      port map(D => \b10_nUT_M9kYfr[7]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \b10_nUT_M9kYfr4\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b10_nUT_M9kYfr[6]_net_1\);
    
    \genblk2.b3_nUT[9]\ : SLE
      port map(D => \b10_nUT_M9kYfr[9]_net_1\, CLK => 
        IICE_comm2iice(8), EN => b9_PKFoLX_ab, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => b6_nUT_IF(9));
    
    \genblk2.b3_nUT[6]\ : SLE
      port map(D => \b10_nUT_M9kYfr[6]_net_1\, CLK => 
        IICE_comm2iice(8), EN => b9_PKFoLX_ab, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => b6_nUT_IF(6));
    
    \b10_nUT_M9kYfr[9]\ : SLE
      port map(D => \b10_nUT_M9kYfr[10]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \b10_nUT_M9kYfr4\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b10_nUT_M9kYfr[9]_net_1\);
    
    b10_nfs_M9kYfr4 : CFG2
      generic map(INIT => x"8")

      port map(A => b7_nUTQ_9u, B => IICE_comm2iice(10), Y => 
        \b10_nfs_M9kYfr4\);
    
    \genblk2.b3_nUT[3]\ : SLE
      port map(D => \b10_nUT_M9kYfr[3]_net_1\, CLK => 
        IICE_comm2iice(8), EN => b9_PKFoLX_ab, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => b6_nUT_IF(3));
    
    \b10_nfs_M9kYfr[2]\ : SLE
      port map(D => \b10_nfs_M9kYfr[3]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \b10_nfs_M9kYfr4\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b10_nfs_M9kYfr[2]_net_1\);
    
    \genblk2.b3_nUT[2]\ : SLE
      port map(D => \b10_nUT_M9kYfr[2]_net_1\, CLK => 
        IICE_comm2iice(8), EN => b9_PKFoLX_ab, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => b6_nUT_IF(2));
    
    \b10_nUT_M9kYfr[3]\ : SLE
      port map(D => \b10_nUT_M9kYfr[4]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \b10_nUT_M9kYfr4\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b10_nUT_M9kYfr[3]_net_1\);
    
    b15_vABZ3qsY_ub3Rme : SLE
      port map(D => IICE_comm2iice(7), CLK => IICE_comm2iice(11), 
        EN => \b15_vABZ3qsY_ub3Rme3\, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b10_vbTtJX_Y2x\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \b10_nfs_M9kYfr[3]\ : SLE
      port map(D => \b10_nfs_M9kYfr[4]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \b10_nfs_M9kYfr4\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b10_nfs_M9kYfr[3]_net_1\);
    
    \genblk1.b3_nfs[3]\ : SLE
      port map(D => \b10_nfs_M9kYfr[3]_net_1\, CLK => 
        IICE_comm2iice(8), EN => b7_nUTQ_9u, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => b6_nfs_IF(3));
    
    \genblk1.b3_nfs_RNIU185[1]\ : CLKINT
      port map(A => \b3_nfs[1]\, Y => \b6_nfs_IF[1]\);
    
    \genblk2.b3_nUT[7]\ : SLE
      port map(D => \b10_nUT_M9kYfr[7]_net_1\, CLK => 
        IICE_comm2iice(8), EN => b9_PKFoLX_ab, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => b6_nUT_IF(7));
    
    \genblk1.b3_nfs[1]\ : SLE
      port map(D => \b10_nfs_M9kYfr[1]_net_1\, CLK => 
        IICE_comm2iice(8), EN => b7_nUTQ_9u, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b3_nfs[1]\);
    
    \b10_nfs_M9kYfr[1]\ : SLE
      port map(D => \b10_nfs_M9kYfr[2]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \b10_nfs_M9kYfr4\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b10_nfs_M9kYfr[1]_net_1\);
    
    \b10_nUT_M9kYfr[4]\ : SLE
      port map(D => \b10_nUT_M9kYfr[5]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \b10_nUT_M9kYfr4\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b10_nUT_M9kYfr[4]_net_1\);
    
    \genblk2.b3_nUT[0]\ : SLE
      port map(D => \b10_PKFoLX_Y2x\, CLK => IICE_comm2iice(8), 
        EN => b9_PKFoLX_ab, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => b6_nUT_IF(0));
    
    \b10_nUT_M9kYfr[1]\ : SLE
      port map(D => \b10_nUT_M9kYfr[2]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \b10_nUT_M9kYfr4\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b10_nUT_M9kYfr[1]_net_1\);
    
    \b10_nUT_M9kYfr[0]\ : SLE
      port map(D => \b10_nUT_M9kYfr[1]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \b10_nUT_M9kYfr4\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \b10_PKFoLX_Y2x\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \genblk2.b3_nUT[8]\ : SLE
      port map(D => \b10_nUT_M9kYfr[8]_net_1\, CLK => 
        IICE_comm2iice(8), EN => b9_PKFoLX_ab, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => b6_nUT_IF(8));
    
    \b10_nfs_M9kYfr[4]\ : SLE
      port map(D => IICE_comm2iice(7), CLK => IICE_comm2iice(11), 
        EN => \b10_nfs_M9kYfr4\, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b10_nfs_M9kYfr[4]_net_1\);
    
    \genblk2.b3_nUT[4]\ : SLE
      port map(D => \b10_nUT_M9kYfr[4]_net_1\, CLK => 
        IICE_comm2iice(8), EN => b9_PKFoLX_ab, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => b6_nUT_IF(4));
    
    \b10_nUT_M9kYfr[11]\ : SLE
      port map(D => IICE_comm2iice(7), CLK => IICE_comm2iice(11), 
        EN => \b10_nUT_M9kYfr4\, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b10_nUT_M9kYfr[11]_net_1\);
    
    \b10_nfs_M9kYfr[0]\ : SLE
      port map(D => \b10_nfs_M9kYfr[1]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \b10_nfs_M9kYfr4\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \b8_nUTQ_XlK\);
    
    \b10_nUT_M9kYfr[7]\ : SLE
      port map(D => \b10_nUT_M9kYfr[8]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \b10_nUT_M9kYfr4\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b10_nUT_M9kYfr[7]_net_1\);
    
    b10_nUT_M9kYfr4 : CFG2
      generic map(INIT => x"8")

      port map(A => b9_PKFoLX_ab, B => IICE_comm2iice(10), Y => 
        \b10_nUT_M9kYfr4\);
    
    \b10_nUT_M9kYfr[8]\ : SLE
      port map(D => \b10_nUT_M9kYfr[9]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \b10_nUT_M9kYfr4\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b10_nUT_M9kYfr[8]_net_1\);
    
    \genblk1.b3_nfs[2]\ : SLE
      port map(D => \b10_nfs_M9kYfr[2]_net_1\, CLK => 
        IICE_comm2iice(8), EN => b7_nUTQ_9u, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => b6_nfs_IF(2));
    
    \genblk1.b3_nfs[0]\ : SLE
      port map(D => \b8_nUTQ_XlK\, CLK => IICE_comm2iice(8), EN
         => b7_nUTQ_9u, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b6_nfs_IF(0));
    
    \genblk3.b8_vABZ3qsY\ : SLE
      port map(D => \b10_vbTtJX_Y2x\, CLK => IICE_comm2iice(8), 
        EN => b9_vbTtJX_ab, ALn => \b6_nfs_IF_i_0\, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => b11_vABZ3qsY_qH);
    
    \b10_nUT_M9kYfr[5]\ : SLE
      port map(D => \b10_nUT_M9kYfr[6]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \b10_nUT_M9kYfr4\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b10_nUT_M9kYfr[5]_net_1\);
    
    \b10_nUT_M9kYfr[10]\ : SLE
      port map(D => \b10_nUT_M9kYfr[11]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \b10_nUT_M9kYfr4\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b10_nUT_M9kYfr[10]_net_1\);
    
    \genblk1.b3_nfs_RNIU185_0[1]\ : CFG1
      generic map(INIT => "01")

      port map(A => \b6_nfs_IF[1]\, Y => \b6_nfs_IF_i_0\);
    
    \genblk2.b3_nUT[5]\ : SLE
      port map(D => \b10_nUT_M9kYfr[5]_net_1\, CLK => 
        IICE_comm2iice(8), EN => b9_PKFoLX_ab, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => b6_nUT_IF(5));
    
    b15_vABZ3qsY_ub3Rme3 : CFG2
      generic map(INIT => x"8")

      port map(A => b9_vbTtJX_ab, B => IICE_comm2iice(10), Y => 
        \b15_vABZ3qsY_ub3Rme3\);
    
    \b10_nUT_M9kYfr[2]\ : SLE
      port map(D => \b10_nUT_M9kYfr[3]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \b10_nUT_M9kYfr4\, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b10_nUT_M9kYfr[2]_net_1\);
    
    \genblk2.b3_nUT[1]\ : SLE
      port map(D => \b10_nUT_M9kYfr[1]_net_1\, CLK => 
        IICE_comm2iice(8), EN => b9_PKFoLX_ab, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => b6_nUT_IF(1));
    
    \genblk2.b3_nUT[11]\ : SLE
      port map(D => \b10_nUT_M9kYfr[11]_net_1\, CLK => 
        IICE_comm2iice(8), EN => b9_PKFoLX_ab, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => b6_nUT_IF(11));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity clock2_en_reg_en_5s_x_0 is

    port( status_b2sclk       : out   std_logic_vector(3 downto 0);
          b6_Ocm0rW           : in    std_logic_vector(2 downto 0);
          b13_nAzGfFM_sLsv3_0 : in    std_logic;
          IICE_comm2iice_0    : in    std_logic;
          b6_nfs_IF_i_0       : in    std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic
        );

end clock2_en_reg_en_5s_x_0;

architecture DEF_ARCH of clock2_en_reg_en_5s_x_0 is 

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \src_ack\, src_ack_i, VCC_net_1, \int_data[1]_net_1\, 
        \dout4\, GND_net_1, \int_data[2]_net_1\, 
        \int_data[3]_net_1\, \int_data[0]_net_1\, \in_en\, 
        \src_req\, \un1_in_en_1\, \dst_req\, \dst_req_d\, 
        \dst_ack\, \in_en4\ : std_logic;

begin 


    un1_in_en_1 : CFG2
      generic map(INIT => x"E")

      port map(A => \in_en\, B => \src_ack\, Y => \un1_in_en_1\);
    
    \dout[1]\ : SLE
      port map(D => \int_data[1]_net_1\, CLK => IICE_comm2iice_0, 
        EN => \dout4\, ALn => b6_nfs_IF_i_0, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => status_b2sclk(1));
    
    dst_ack : CFG2
      generic map(INIT => x"E")

      port map(A => \dst_req\, B => \dst_req_d\, Y => \dst_ack\);
    
    \dout[3]\ : SLE
      port map(D => \int_data[3]_net_1\, CLK => IICE_comm2iice_0, 
        EN => \dout4\, ALn => b6_nfs_IF_i_0, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => status_b2sclk(3));
    
    \int_data[1]\ : SLE
      port map(D => b6_Ocm0rW(1), CLK => CommsFPGA_CCC_0_GL0, EN
         => \in_en\, ALn => b6_nfs_IF_i_0, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \int_data[1]_net_1\);
    
    \dout[2]\ : SLE
      port map(D => \int_data[2]_net_1\, CLK => IICE_comm2iice_0, 
        EN => \dout4\, ALn => b6_nfs_IF_i_0, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => status_b2sclk(2));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    in_en : SLE
      port map(D => \in_en4\, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => b6_nfs_IF_i_0, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \in_en\);
    
    src_ack : SLE
      port map(D => \dst_ack\, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => b6_nfs_IF_i_0, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \src_ack\);
    
    \int_data[0]\ : SLE
      port map(D => b6_Ocm0rW(0), CLK => CommsFPGA_CCC_0_GL0, EN
         => \in_en\, ALn => b6_nfs_IF_i_0, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \int_data[0]_net_1\);
    
    \int_data[2]\ : SLE
      port map(D => b6_Ocm0rW(2), CLK => CommsFPGA_CCC_0_GL0, EN
         => \in_en\, ALn => b6_nfs_IF_i_0, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \int_data[2]_net_1\);
    
    \dout[0]\ : SLE
      port map(D => \int_data[0]_net_1\, CLK => IICE_comm2iice_0, 
        EN => \dout4\, ALn => b6_nfs_IF_i_0, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => status_b2sclk(0));
    
    dst_req : SLE
      port map(D => \src_req\, CLK => IICE_comm2iice_0, EN => 
        VCC_net_1, ALn => b6_nfs_IF_i_0, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \dst_req\);
    
    src_req_RNO : CFG1
      generic map(INIT => "01")

      port map(A => \src_ack\, Y => src_ack_i);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \int_data[3]\ : SLE
      port map(D => b13_nAzGfFM_sLsv3_0, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \in_en\, ALn => b6_nfs_IF_i_0, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \int_data[3]_net_1\);
    
    dout4 : CFG2
      generic map(INIT => x"2")

      port map(A => \dst_req\, B => \dst_req_d\, Y => \dout4\);
    
    src_req : SLE
      port map(D => src_ack_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_in_en_1\, ALn => b6_nfs_IF_i_0, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \src_req\);
    
    in_en4 : CFG3
      generic map(INIT => x"01")

      port map(A => \src_req\, B => \in_en\, C => \src_ack\, Y
         => \in_en4\);
    
    dst_req_d : SLE
      port map(D => \dst_req\, CLK => IICE_comm2iice_0, EN => 
        VCC_net_1, ALn => b6_nfs_IF_i_0, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \dst_req_d\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b7_OCByLXC_Z1_x_0 is

    port( IICE_comm2iice      : in    std_logic_vector(11 downto 7);
          b9_PKFoLX_ab        : in    std_logic;
          b8_nUTQ_XlK         : out   std_logic;
          b7_nUTQ_9u          : in    std_logic;
          b10_PKFoLX_Y2x      : out   std_logic;
          b10_vbTtJX_Y2x      : out   std_logic;
          b9_vbTtJX_ab        : in    std_logic;
          b8_ubTt3_YG         : in    std_logic;
          N_145_i             : out   std_logic;
          b13_wRBtT_ME83hHx   : in    std_logic;
          b9_ubTt3_Mxf        : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          b5_voSc3_i          : out   std_logic;
          b5_voSc3            : out   std_logic
        );

end b7_OCByLXC_Z1_x_0;

architecture DEF_ARCH of b7_OCByLXC_Z1_x_0 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component b8_nR_ymqrG_12s_5s_0_0s_0s_1_2046_x_0
    port( IICE_comm2iice  : in    std_logic_vector(11 downto 7) := (others => 'U');
          b6_nUT_IF       : out   std_logic_vector(11 downto 0);
          b6_nfs_IF       : out   std_logic_vector(4 downto 0);
          b6_nfs_IF_i_0   : out   std_logic;
          b9_vbTtJX_ab    : in    std_logic := 'U';
          b11_vABZ3qsY_qH : out   std_logic;
          b10_vbTtJX_Y2x  : out   std_logic;
          b10_PKFoLX_Y2x  : out   std_logic;
          b7_nUTQ_9u      : in    std_logic := 'U';
          b8_nUTQ_XlK     : out   std_logic;
          b9_PKFoLX_ab    : in    std_logic := 'U'
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component clock2_en_reg_en_5s_x_0
    port( status_b2sclk       : out   std_logic_vector(3 downto 0);
          b6_Ocm0rW           : in    std_logic_vector(2 downto 0) := (others => 'U');
          b13_nAzGfFM_sLsv3_0 : in    std_logic := 'U';
          IICE_comm2iice_0    : in    std_logic := 'U';
          b6_nfs_IF_i_0       : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U'
        );
  end component;

    signal \b5_voSc3\, \b12_voSc3_gmasbb\, 
        \b15_uRrc2XfY_rbN_gs[24]_net_1\, VCC_net_1, 
        \b15_uRrc2XfY_rbN_gr[24]_net_1\, GND_net_1, 
        \b15_uRrc2XfY_rbN_gs[25]_net_1\, 
        \b15_uRrc2XfY_rbN_gr[25]_net_1\, 
        \b15_uRrc2XfY_rbN_gs[26]_net_1\, 
        \b15_uRrc2XfY_rbN_gr[26]_net_1\, 
        \b15_uRrc2XfY_rbN_gs[27]_net_1\, 
        \b15_uRrc2XfY_rbN_gr[27]_net_1\, \b3_nfs[0]_net_1\, 
        \b6_nfs_IF[0]\, \b3_nfs[1]_net_1\, \b6_nfs_IF[1]\, 
        \b3_nfs[2]_net_1\, \b6_nfs_IF[2]\, \b3_nfs[3]_net_1\, 
        \b6_nfs_IF[3]\, \b3_nfs[4]_net_1\, \b6_nfs_IF[4]\, 
        \b15_uRrc2XfY_rbN_gs[9]_net_1\, 
        \b15_uRrc2XfY_rbN_gr[9]_net_1\, 
        \b15_uRrc2XfY_rbN_gs[10]_net_1\, 
        \b15_uRrc2XfY_rbN_gr[10]_net_1\, 
        \b15_uRrc2XfY_rbN_gs[11]_net_1\, 
        \b15_uRrc2XfY_rbN_gr[11]_net_1\, 
        \b15_uRrc2XfY_rbN_gs[12]_net_1\, 
        \b15_uRrc2XfY_rbN_gr[12]_net_1\, 
        \b15_uRrc2XfY_rbN_gs[13]_net_1\, 
        \b15_uRrc2XfY_rbN_gr[13]_net_1\, 
        \b15_uRrc2XfY_rbN_gs[14]_net_1\, 
        \b15_uRrc2XfY_rbN_gr[14]_net_1\, 
        \b15_uRrc2XfY_rbN_gs[15]_net_1\, 
        \b15_uRrc2XfY_rbN_gr[15]_net_1\, 
        \b15_uRrc2XfY_rbN_gs[16]_net_1\, 
        \b15_uRrc2XfY_rbN_gr[16]_net_1\, 
        \b15_uRrc2XfY_rbN_gs[17]_net_1\, 
        \b15_uRrc2XfY_rbN_gr[17]_net_1\, 
        \b15_uRrc2XfY_rbN_gs[18]_net_1\, 
        \b15_uRrc2XfY_rbN_gr[18]_net_1\, 
        \b15_uRrc2XfY_rbN_gs[19]_net_1\, 
        \b15_uRrc2XfY_rbN_gr[19]_net_1\, 
        \b15_uRrc2XfY_rbN_gs[20]_net_1\, 
        \b15_uRrc2XfY_rbN_gr[20]_net_1\, 
        \b15_uRrc2XfY_rbN_gs[21]_net_1\, 
        \b15_uRrc2XfY_rbN_gr[21]_net_1\, 
        \b15_uRrc2XfY_rbN_gs[22]_net_1\, 
        \b15_uRrc2XfY_rbN_gr[22]_net_1\, 
        \b15_uRrc2XfY_rbN_gs[23]_net_1\, 
        \b15_uRrc2XfY_rbN_gr[23]_net_1\, \b7_nYhI39s[5]_net_1\, 
        \b7_nYhI39s[6]_net_1\, \b7_nYhI39s[7]_net_1\, 
        \b7_nYhI39s[8]_net_1\, \b7_nYhI39s[9]_net_1\, 
        \b7_nYhI39s[10]_net_1\, \b7_nYhI39s[11]_net_1\, 
        \b15_uRrc2XfY_rbN_gs[0]_net_1\, 
        \b15_uRrc2XfY_rbN_gr[0]_net_1\, 
        \b15_uRrc2XfY_rbN_gs[1]_net_1\, 
        \b15_uRrc2XfY_rbN_gr[1]_net_1\, 
        \b15_uRrc2XfY_rbN_gs[2]_net_1\, 
        \b15_uRrc2XfY_rbN_gr[2]_net_1\, 
        \b15_uRrc2XfY_rbN_gs[3]_net_1\, 
        \b15_uRrc2XfY_rbN_gr[3]_net_1\, 
        \b15_uRrc2XfY_rbN_gs[5]_net_1\, 
        \b15_uRrc2XfY_rbN_gr[5]_net_1\, 
        \b15_uRrc2XfY_rbN_gs[6]_net_1\, 
        \b15_uRrc2XfY_rbN_gr[6]_net_1\, 
        \b15_uRrc2XfY_rbN_gs[7]_net_1\, 
        \b15_uRrc2XfY_rbN_gr[7]_net_1\, 
        \b15_uRrc2XfY_rbN_gs[8]_net_1\, 
        \b15_uRrc2XfY_rbN_gr[8]_net_1\, N_144_i, N_151_i, 
        \un13[2]_net_1\, \b13_nAzGfFM_sLsv3[5]_net_1\, 
        b11_vABZ3qsY_qH, \b7_nYhI39s[0]_net_1\, 
        \b7_nYhI39s[1]_net_1\, \b7_nYhI39s[2]_net_1\, 
        \b7_nYhI39s[3]_net_1\, \b7_nYhI39s[4]_net_1\, 
        \status_b2sclk[0]\, \status_b2sclk[1]\, 
        \status_b2sclk[2]\, \status_b2sclk[3]\, 
        \b13_nAzGfFM_sLsv3[2]_net_1\, 
        \b12_uRrc2XfY_rbN[27]_net_1\, 
        \b12_uRrc2XfY_rbN_5[27]_net_1\, 
        \un1_b12_uRrc2XfY_rbN10_i\, \b3_nUT[0]_net_1\, 
        \b6_nfs_IF_i[1]\, \b6_nUT_IF[0]\, \b3_nUT[1]_net_1\, 
        \b6_nUT_IF[1]\, \b3_nUT[2]_net_1\, \b6_nUT_IF[2]\, 
        \b3_nUT[3]_net_1\, \b6_nUT_IF[3]\, \b3_nUT[4]_net_1\, 
        \b6_nUT_IF[4]\, \b3_nUT[5]_net_1\, \b6_nUT_IF[5]\, 
        \b3_nUT[6]_net_1\, \b6_nUT_IF[6]\, \b3_nUT[7]_net_1\, 
        \b6_nUT_IF[7]\, \b3_nUT[8]_net_1\, \b6_nUT_IF[8]\, 
        \b3_nUT[9]_net_1\, \b6_nUT_IF[9]\, \b3_nUT[10]_net_1\, 
        \b6_nUT_IF[10]\, \b3_nUT[11]_net_1\, \b6_nUT_IF[11]\, 
        \b12_uRrc2XfY_rbN[12]_net_1\, 
        \b12_uRrc2XfY_rbN_5[12]_net_1\, 
        \b12_uRrc2XfY_rbN[13]_net_1\, 
        \b12_uRrc2XfY_rbN_5[13]_net_1\, 
        \b12_uRrc2XfY_rbN[14]_net_1\, 
        \b12_uRrc2XfY_rbN_5[14]_net_1\, 
        \b12_uRrc2XfY_rbN[15]_net_1\, 
        \b12_uRrc2XfY_rbN_5[15]_net_1\, 
        \b12_uRrc2XfY_rbN[16]_net_1\, 
        \b12_uRrc2XfY_rbN_5[16]_net_1\, 
        \b12_uRrc2XfY_rbN[17]_net_1\, 
        \b12_uRrc2XfY_rbN_5[17]_net_1\, 
        \b12_uRrc2XfY_rbN[18]_net_1\, 
        \b12_uRrc2XfY_rbN_5[18]_net_1\, 
        \b12_uRrc2XfY_rbN[19]_net_1\, 
        \b12_uRrc2XfY_rbN_5[19]_net_1\, 
        \b12_uRrc2XfY_rbN[20]_net_1\, 
        \b12_uRrc2XfY_rbN_5[20]_net_1\, 
        \b12_uRrc2XfY_rbN[21]_net_1\, 
        \b12_uRrc2XfY_rbN_5[21]_net_1\, 
        \b12_uRrc2XfY_rbN[22]_net_1\, 
        \b12_uRrc2XfY_rbN_5[22]_net_1\, 
        \b12_uRrc2XfY_rbN[23]_net_1\, 
        \b12_uRrc2XfY_rbN_5[23]_net_1\, 
        \b12_uRrc2XfY_rbN[24]_net_1\, 
        \b12_uRrc2XfY_rbN_5[24]_net_1\, 
        \b12_uRrc2XfY_rbN[25]_net_1\, 
        \b12_uRrc2XfY_rbN_5[25]_net_1\, 
        \b12_uRrc2XfY_rbN[26]_net_1\, 
        \b12_uRrc2XfY_rbN_5[26]_net_1\, 
        \b12_uRrc2XfY_rbN_5[0]_net_1\, 
        \b12_uRrc2XfY_rbN[1]_net_1\, 
        \b12_uRrc2XfY_rbN_5[1]_net_1\, 
        \b12_uRrc2XfY_rbN[2]_net_1\, 
        \b12_uRrc2XfY_rbN_5[2]_net_1\, 
        \b12_uRrc2XfY_rbN[3]_net_1\, 
        \b12_uRrc2XfY_rbN_5[3]_net_1\, 
        \b12_uRrc2XfY_rbN[4]_net_1\, 
        \b12_uRrc2XfY_rbN_5[4]_net_1\, 
        \b12_uRrc2XfY_rbN[5]_net_1\, 
        \b12_uRrc2XfY_rbN_5[5]_net_1\, 
        \b12_uRrc2XfY_rbN[6]_net_1\, 
        \b12_uRrc2XfY_rbN_5[6]_net_1\, 
        \b12_uRrc2XfY_rbN[7]_net_1\, 
        \b12_uRrc2XfY_rbN_5[7]_net_1\, 
        \b12_uRrc2XfY_rbN[8]_net_1\, 
        \b12_uRrc2XfY_rbN_5[8]_net_1\, 
        \b12_uRrc2XfY_rbN[9]_net_1\, 
        \b12_uRrc2XfY_rbN_5[9]_net_1\, 
        \b12_uRrc2XfY_rbN[10]_net_1\, 
        \b12_uRrc2XfY_rbN_5[10]_net_1\, 
        \b12_uRrc2XfY_rbN[11]_net_1\, 
        \b12_uRrc2XfY_rbN_5[11]_net_1\, b10_nYhI3_umjB, 
        \b10_nYhI3_umjB_1\, \b13_nAzGfFM_sLsv3[0]_net_1\, 
        \b13_nAzGfFM_sLsv3[1]_net_1\, 
        \b13_nAzGfFM_sLsv3_ns[1]_net_1\, 
        \b13_nAzGfFM_sLsv3_ns[2]_net_1\, 
        \b13_nAzGfFM_sLsv3[3]_net_1\, \b13_nAzGfFM_sLsv3_ns[3]\, 
        \b13_nAzGfFM_sLsv3[4]_net_1\, 
        \b13_nAzGfFM_sLsv3_ns[4]_net_1\, 
        \b13_nAzGfFM_sLsv3_ns[5]_net_1\, \b8_vABZ3qsY\, 
        \b7_nYhI39s_lm[0]\, b7_nYhI39se, \b7_nYhI39s_lm[1]\, 
        \b7_nYhI39s_lm[2]\, \b7_nYhI39s_lm[3]\, 
        \b7_nYhI39s_lm[4]\, \b7_nYhI39s_lm[5]\, 
        \b7_nYhI39s_lm[6]\, \b7_nYhI39s_lm[7]\, 
        \b7_nYhI39s_lm[8]\, \b7_nYhI39s_lm[9]\, 
        \b7_nYhI39s_lm[10]\, \b7_nYhI39s_lm[11]\, 
        \b7_nYhI39s_cry[0]_net_1\, \b7_nYhI39s_cry_Y[0]\, 
        \b7_nYhI39s_cry[1]_net_1\, \b7_nYhI39s_s[1]\, 
        \b7_nYhI39s_cry[2]_net_1\, \b7_nYhI39s_s[2]\, 
        \b7_nYhI39s_cry[3]_net_1\, \b7_nYhI39s_s[3]\, 
        \b7_nYhI39s_cry[4]_net_1\, \b7_nYhI39s_s[4]\, 
        \b7_nYhI39s_cry[5]_net_1\, \b7_nYhI39s_s[5]\, 
        \b7_nYhI39s_cry[6]_net_1\, \b7_nYhI39s_s[6]\, 
        \b7_nYhI39s_cry[7]_net_1\, \b7_nYhI39s_s[7]\, 
        \b7_nYhI39s_cry[8]_net_1\, \b7_nYhI39s_s[8]\, 
        \b7_nYhI39s_cry[9]_net_1\, \b7_nYhI39s_s[9]\, 
        \b7_nYhI39s_s[11]_net_1\, \b7_nYhI39s_cry[10]_net_1\, 
        \b7_nYhI39s_s[10]\, N_74, \b6_Ocm0rW[2]\, 
        b7_nYhI39slde_1_0, N_61, N_63_2, N_324, 
        \b10_nYhI3_umjB_0_sqmuxa_8\, \b10_nYhI3_umjB_0_sqmuxa_7\, 
        \b10_nYhI3_umjB_0_sqmuxa_6\, N_62, N_71, \b6_Ocm0rW[0]\, 
        N_140, \b6_Ocm0rW[1]\, b10_xoU0_WMrtX_0_sqmuxa_1, 
        b6_nUT_fF, N_86, \b10_nYhI3_umjB_0_sqmuxa\ : std_logic;
    signal nc1 : std_logic;

    for all : b8_nR_ymqrG_12s_5s_0_0s_0s_1_2046_x_0
	Use entity work.b8_nR_ymqrG_12s_5s_0_0s_0s_1_2046_x_0(DEF_ARCH);
    for all : clock2_en_reg_en_5s_x_0
	Use entity work.clock2_en_reg_en_5s_x_0(DEF_ARCH);
begin 

    b5_voSc3 <= \b5_voSc3\;

    \b3_nUT[0]\ : SLE
      port map(D => \b6_nUT_IF[0]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => \b6_nfs_IF_i[1]\, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b3_nUT[0]_net_1\);
    
    \b12_uRrc2XfY_rbN_5[6]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \b12_uRrc2XfY_rbN[7]_net_1\, B => 
        IICE_comm2iice(9), C => \b15_uRrc2XfY_rbN_gs[6]_net_1\, Y
         => \b12_uRrc2XfY_rbN_5[6]_net_1\);
    
    b10_nYhI3_umjB_0_sqmuxa_6 : CFG4
      generic map(INIT => x"0001")

      port map(A => \b7_nYhI39s[11]_net_1\, B => 
        \b7_nYhI39s[8]_net_1\, C => \b7_nYhI39s[6]_net_1\, D => 
        \b7_nYhI39s[2]_net_1\, Y => \b10_nYhI3_umjB_0_sqmuxa_6\);
    
    \b15_uRrc2XfY_rbN_gs[12]\ : SLE
      port map(D => \b15_uRrc2XfY_rbN_gr[12]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gs[12]_net_1\);
    
    \b12_uRrc2XfY_rbN[11]\ : SLE
      port map(D => \b12_uRrc2XfY_rbN_5[11]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \un1_b12_uRrc2XfY_rbN10_i\, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b12_uRrc2XfY_rbN[11]_net_1\);
    
    \b15_uRrc2XfY_rbN_gr[0]\ : SLE
      port map(D => \status_b2sclk[0]\, CLK => IICE_comm2iice(11), 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b15_uRrc2XfY_rbN_gr[0]_net_1\);
    
    b11_nUTGT_khWqH : b8_nR_ymqrG_12s_5s_0_0s_0s_1_2046_x_0
      port map(IICE_comm2iice(11) => IICE_comm2iice(11), 
        IICE_comm2iice(10) => IICE_comm2iice(10), 
        IICE_comm2iice(9) => nc1, IICE_comm2iice(8) => 
        IICE_comm2iice(8), IICE_comm2iice(7) => IICE_comm2iice(7), 
        b6_nUT_IF(11) => \b6_nUT_IF[11]\, b6_nUT_IF(10) => 
        \b6_nUT_IF[10]\, b6_nUT_IF(9) => \b6_nUT_IF[9]\, 
        b6_nUT_IF(8) => \b6_nUT_IF[8]\, b6_nUT_IF(7) => 
        \b6_nUT_IF[7]\, b6_nUT_IF(6) => \b6_nUT_IF[6]\, 
        b6_nUT_IF(5) => \b6_nUT_IF[5]\, b6_nUT_IF(4) => 
        \b6_nUT_IF[4]\, b6_nUT_IF(3) => \b6_nUT_IF[3]\, 
        b6_nUT_IF(2) => \b6_nUT_IF[2]\, b6_nUT_IF(1) => 
        \b6_nUT_IF[1]\, b6_nUT_IF(0) => \b6_nUT_IF[0]\, 
        b6_nfs_IF(4) => \b6_nfs_IF[4]\, b6_nfs_IF(3) => 
        \b6_nfs_IF[3]\, b6_nfs_IF(2) => \b6_nfs_IF[2]\, 
        b6_nfs_IF(1) => \b6_nfs_IF[1]\, b6_nfs_IF(0) => 
        \b6_nfs_IF[0]\, b6_nfs_IF_i_0 => \b6_nfs_IF_i[1]\, 
        b9_vbTtJX_ab => b9_vbTtJX_ab, b11_vABZ3qsY_qH => 
        b11_vABZ3qsY_qH, b10_vbTtJX_Y2x => b10_vbTtJX_Y2x, 
        b10_PKFoLX_Y2x => b10_PKFoLX_Y2x, b7_nUTQ_9u => 
        b7_nUTQ_9u, b8_nUTQ_XlK => b8_nUTQ_XlK, b9_PKFoLX_ab => 
        b9_PKFoLX_ab);
    
    \b3_nUT[6]\ : SLE
      port map(D => \b6_nUT_IF[6]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => \b6_nfs_IF_i[1]\, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b3_nUT[6]_net_1\);
    
    \b7_nYhI39s_lm_0[6]\ : CFG4
      generic map(INIT => x"AAC0")

      port map(A => \b7_nYhI39s_s[6]\, B => \b3_nUT[6]_net_1\, C
         => N_71, D => b6_nUT_fF, Y => \b7_nYhI39s_lm[6]\);
    
    b12_voSc3_gmasbb_RNI0GM6 : CLKINT
      port map(A => \b12_voSc3_gmasbb\, Y => \b5_voSc3\);
    
    b10_xoU0_WMrtX_0_sqmuxa : CFG3
      generic map(INIT => x"80")

      port map(A => b10_nYhI3_umjB, B => N_62, C => N_61, Y => 
        N_74);
    
    \b12_uRrc2XfY_rbN_5[17]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \b12_uRrc2XfY_rbN[18]_net_1\, B => 
        IICE_comm2iice(9), C => \b15_uRrc2XfY_rbN_gs[17]_net_1\, 
        Y => \b12_uRrc2XfY_rbN_5[17]_net_1\);
    
    \b12_uRrc2XfY_rbN[4]\ : SLE
      port map(D => \b12_uRrc2XfY_rbN_5[4]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \un1_b12_uRrc2XfY_rbN10_i\, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b12_uRrc2XfY_rbN[4]_net_1\);
    
    \b3_nUT[11]\ : SLE
      port map(D => \b6_nUT_IF[11]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => \b6_nfs_IF_i[1]\, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b3_nUT[11]_net_1\);
    
    \b12_uRrc2XfY_rbN[0]\ : SLE
      port map(D => \b12_uRrc2XfY_rbN_5[0]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \un1_b12_uRrc2XfY_rbN10_i\, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => b9_ubTt3_Mxf);
    
    \b15_uRrc2XfY_rbN_gs[1]\ : SLE
      port map(D => \b15_uRrc2XfY_rbN_gr[1]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gs[1]_net_1\);
    
    \b15_uRrc2XfY_rbN_gs[10]\ : SLE
      port map(D => \b15_uRrc2XfY_rbN_gr[10]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gs[10]_net_1\);
    
    \b3_nfs[1]\ : SLE
      port map(D => \b6_nfs_IF[1]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b3_nfs[1]_net_1\);
    
    b10_nYhI3_umjB_0_sqmuxa_8 : CFG4
      generic map(INIT => x"0001")

      port map(A => \b7_nYhI39s[7]_net_1\, B => 
        \b7_nYhI39s[5]_net_1\, C => \b7_nYhI39s[4]_net_1\, D => 
        \b7_nYhI39s[3]_net_1\, Y => \b10_nYhI3_umjB_0_sqmuxa_8\);
    
    \b7_nYhI39s_cry[2]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \b7_nYhI39s[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \b7_nYhI39s_cry[1]_net_1\, S => \b7_nYhI39s_s[2]\, Y => 
        OPEN, FCO => \b7_nYhI39s_cry[2]_net_1\);
    
    \b15_uRrc2XfY_rbN_gs[5]\ : SLE
      port map(D => \b15_uRrc2XfY_rbN_gr[5]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gs[5]_net_1\);
    
    \b15_uRrc2XfY_rbN_gs[27]\ : SLE
      port map(D => \b15_uRrc2XfY_rbN_gr[27]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gs[27]_net_1\);
    
    \b7_nYhI39s_cry[8]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \b7_nYhI39s[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \b7_nYhI39s_cry[7]_net_1\, S => \b7_nYhI39s_s[8]\, Y => 
        OPEN, FCO => \b7_nYhI39s_cry[8]_net_1\);
    
    \b15_uRrc2XfY_rbN_gr[18]\ : SLE
      port map(D => \b7_nYhI39s[2]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gr[18]_net_1\);
    
    \b12_uRrc2XfY_rbN[14]\ : SLE
      port map(D => \b12_uRrc2XfY_rbN_5[14]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \un1_b12_uRrc2XfY_rbN10_i\, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b12_uRrc2XfY_rbN[14]_net_1\);
    
    \b7_nYhI39s[3]\ : SLE
      port map(D => \b7_nYhI39s_lm[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b7_nYhI39se, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b7_nYhI39s[3]_net_1\);
    
    \b15_uRrc2XfY_rbN_gr[23]\ : SLE
      port map(D => \b7_nYhI39s[7]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gr[23]_net_1\);
    
    \b12_uRrc2XfY_rbN_5[26]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \b12_uRrc2XfY_rbN[27]_net_1\, B => 
        IICE_comm2iice(9), C => \b15_uRrc2XfY_rbN_gs[26]_net_1\, 
        Y => \b12_uRrc2XfY_rbN_5[26]_net_1\);
    
    \b15_uRrc2XfY_rbN_gs[24]\ : SLE
      port map(D => \b15_uRrc2XfY_rbN_gr[24]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gs[24]_net_1\);
    
    \b13_nAzGfFM_sLsv3[0]\ : SLE
      port map(D => GND_net_1, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => \b6_nfs_IF_i[1]\, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b13_nAzGfFM_sLsv3[0]_net_1\);
    
    \b12_uRrc2XfY_rbN[13]\ : SLE
      port map(D => \b12_uRrc2XfY_rbN_5[13]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \un1_b12_uRrc2XfY_rbN10_i\, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b12_uRrc2XfY_rbN[13]_net_1\);
    
    \b13_nAzGfFM_sLsv3[1]\ : SLE
      port map(D => \b13_nAzGfFM_sLsv3_ns[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        \b6_nfs_IF_i[1]\, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \b13_nAzGfFM_sLsv3[1]_net_1\);
    
    \b12_uRrc2XfY_rbN[25]\ : SLE
      port map(D => \b12_uRrc2XfY_rbN_5[25]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \un1_b12_uRrc2XfY_rbN10_i\, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b12_uRrc2XfY_rbN[25]_net_1\);
    
    \b15_uRrc2XfY_rbN_gr[13]\ : SLE
      port map(D => \un13[2]_net_1\, CLK => IICE_comm2iice(11), 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b15_uRrc2XfY_rbN_gr[13]_net_1\);
    
    \b13_nAzGfFM_sLsv3_ns_a3[3]\ : CFG2
      generic map(INIT => x"2")

      port map(A => N_140, B => b10_nYhI3_umjB, Y => 
        \b13_nAzGfFM_sLsv3_ns[3]\);
    
    b10_nYhI3_umjB_0_sqmuxa : CFG4
      generic map(INIT => x"8000")

      port map(A => \b10_nYhI3_umjB_0_sqmuxa_8\, B => 
        \b10_nYhI3_umjB_0_sqmuxa_7\, C => b6_nUT_fF, D => 
        \b10_nYhI3_umjB_0_sqmuxa_6\, Y => 
        \b10_nYhI3_umjB_0_sqmuxa\);
    
    \b15_uRrc2XfY_rbN_gr_RNO[12]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \b13_nAzGfFM_sLsv3[2]_net_1\, B => 
        \b13_nAzGfFM_sLsv3[3]_net_1\, Y => N_151_i);
    
    \b15_uRrc2XfY_rbN_gs[19]\ : SLE
      port map(D => \b15_uRrc2XfY_rbN_gr[19]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gs[19]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \b12_uRrc2XfY_rbN_5[23]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \b12_uRrc2XfY_rbN[24]_net_1\, B => 
        IICE_comm2iice(9), C => \b15_uRrc2XfY_rbN_gs[23]_net_1\, 
        Y => \b12_uRrc2XfY_rbN_5[23]_net_1\);
    
    \b12_uRrc2XfY_rbN[19]\ : SLE
      port map(D => \b12_uRrc2XfY_rbN_5[19]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \un1_b12_uRrc2XfY_rbN10_i\, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b12_uRrc2XfY_rbN[19]_net_1\);
    
    \b12_uRrc2XfY_rbN_5[24]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \b12_uRrc2XfY_rbN[25]_net_1\, B => 
        IICE_comm2iice(9), C => \b15_uRrc2XfY_rbN_gs[24]_net_1\, 
        Y => \b12_uRrc2XfY_rbN_5[24]_net_1\);
    
    \b7_nYhI39s_cry[5]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \b7_nYhI39s[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \b7_nYhI39s_cry[4]_net_1\, S => \b7_nYhI39s_s[5]\, Y => 
        OPEN, FCO => \b7_nYhI39s_cry[5]_net_1\);
    
    \b15_uRrc2XfY_rbN_gs[25]\ : SLE
      port map(D => \b15_uRrc2XfY_rbN_gr[25]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gs[25]_net_1\);
    
    \b12_uRrc2XfY_rbN[6]\ : SLE
      port map(D => \b12_uRrc2XfY_rbN_5[6]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \un1_b12_uRrc2XfY_rbN10_i\, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b12_uRrc2XfY_rbN[6]_net_1\);
    
    \b3_nUT[1]\ : SLE
      port map(D => \b6_nUT_IF[1]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => \b6_nfs_IF_i[1]\, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b3_nUT[1]_net_1\);
    
    \b15_uRrc2XfY_rbN_gs[17]\ : SLE
      port map(D => \b15_uRrc2XfY_rbN_gr[17]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gs[17]_net_1\);
    
    \b7_nYhI39s[6]\ : SLE
      port map(D => \b7_nYhI39s_lm[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b7_nYhI39se, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b7_nYhI39s[6]_net_1\);
    
    \b15_uRrc2XfY_rbN_gs[6]\ : SLE
      port map(D => \b15_uRrc2XfY_rbN_gr[6]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gs[6]_net_1\);
    
    \b15_uRrc2XfY_rbN_gs[14]\ : SLE
      port map(D => \b15_uRrc2XfY_rbN_gr[14]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gs[14]_net_1\);
    
    \b7_nYhI39s_lm_0[0]\ : CFG4
      generic map(INIT => x"AAC0")

      port map(A => \b7_nYhI39s_cry_Y[0]\, B => \b3_nUT[0]_net_1\, 
        C => N_71, D => b6_nUT_fF, Y => \b7_nYhI39s_lm[0]\);
    
    b6_nUT_fF_0_sqmuxa : CFG3
      generic map(INIT => x"80")

      port map(A => \b13_nAzGfFM_sLsv3[1]_net_1\, B => N_61, C
         => b10_nYhI3_umjB, Y => N_71);
    
    \b12_uRrc2XfY_rbN[8]\ : SLE
      port map(D => \b12_uRrc2XfY_rbN_5[8]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \un1_b12_uRrc2XfY_rbN10_i\, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b12_uRrc2XfY_rbN[8]_net_1\);
    
    un1_b12_uRrc2XfY_rbN10_i : CFG3
      generic map(INIT => x"E0")

      port map(A => IICE_comm2iice(10), B => IICE_comm2iice(9), C
         => b8_ubTt3_YG, Y => \un1_b12_uRrc2XfY_rbN10_i\);
    
    \b7_nYhI39s[5]\ : SLE
      port map(D => \b7_nYhI39s_lm[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b7_nYhI39se, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b7_nYhI39s[5]_net_1\);
    
    \b12_uRrc2XfY_rbN[1]\ : SLE
      port map(D => \b12_uRrc2XfY_rbN_5[1]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \un1_b12_uRrc2XfY_rbN10_i\, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b12_uRrc2XfY_rbN[1]_net_1\);
    
    \b15_uRrc2XfY_rbN_gr[3]\ : SLE
      port map(D => \status_b2sclk[3]\, CLK => IICE_comm2iice(11), 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b15_uRrc2XfY_rbN_gr[3]_net_1\);
    
    \b13_nAzGfFM_sLsv3_RNIVBP6[2]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \b13_nAzGfFM_sLsv3[2]_net_1\, B => 
        \b13_nAzGfFM_sLsv3[3]_net_1\, C => 
        \b13_nAzGfFM_sLsv3[1]_net_1\, Y => N_145_i);
    
    \b7_nYhI39s_cry[10]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \b7_nYhI39s[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \b7_nYhI39s_cry[9]_net_1\, S => \b7_nYhI39s_s[10]\, Y => 
        OPEN, FCO => \b7_nYhI39s_cry[10]_net_1\);
    
    \b3_nUT[3]\ : SLE
      port map(D => \b6_nUT_IF[3]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => \b6_nfs_IF_i[1]\, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b3_nUT[3]_net_1\);
    
    \b15_uRrc2XfY_rbN_gs[15]\ : SLE
      port map(D => \b15_uRrc2XfY_rbN_gr[15]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gs[15]_net_1\);
    
    \b15_uRrc2XfY_rbN_gr[22]\ : SLE
      port map(D => \b7_nYhI39s[6]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gr[22]_net_1\);
    
    \b3_nfs[0]\ : SLE
      port map(D => \b6_nfs_IF[0]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b3_nfs[0]_net_1\);
    
    \b12_uRrc2XfY_rbN_5[22]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \b12_uRrc2XfY_rbN[23]_net_1\, B => 
        IICE_comm2iice(9), C => \b15_uRrc2XfY_rbN_gs[22]_net_1\, 
        Y => \b12_uRrc2XfY_rbN_5[22]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \b7_nYhI39s_lm_0[2]\ : CFG4
      generic map(INIT => x"AAC0")

      port map(A => \b7_nYhI39s_s[2]\, B => \b3_nUT[2]_net_1\, C
         => N_71, D => b6_nUT_fF, Y => \b7_nYhI39s_lm[2]\);
    
    \b12_uRrc2XfY_rbN_5[1]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \b12_uRrc2XfY_rbN[2]_net_1\, B => 
        IICE_comm2iice(9), C => \b15_uRrc2XfY_rbN_gs[1]_net_1\, Y
         => \b12_uRrc2XfY_rbN_5[1]_net_1\);
    
    \b15_uRrc2XfY_rbN_gr_RNO[11]\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \b13_nAzGfFM_sLsv3[5]_net_1\, B => 
        \b13_nAzGfFM_sLsv3[3]_net_1\, C => 
        \b13_nAzGfFM_sLsv3[1]_net_1\, Y => N_144_i);
    
    \b7_nYhI39s_s[11]\ : ARI1
      generic map(INIT => x"45500")

      port map(A => VCC_net_1, B => \b7_nYhI39s[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \b7_nYhI39s_cry[10]_net_1\, S => \b7_nYhI39s_s[11]_net_1\, 
        Y => OPEN, FCO => OPEN);
    
    \b15_uRrc2XfY_rbN_gr[12]\ : SLE
      port map(D => N_151_i, CLK => IICE_comm2iice(11), EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b15_uRrc2XfY_rbN_gr[12]_net_1\);
    
    \b12_uRrc2XfY_rbN_5[2]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \b12_uRrc2XfY_rbN[3]_net_1\, B => 
        IICE_comm2iice(9), C => \b15_uRrc2XfY_rbN_gs[2]_net_1\, Y
         => \b12_uRrc2XfY_rbN_5[2]_net_1\);
    
    \b15_uRrc2XfY_rbN_gs[9]\ : SLE
      port map(D => \b15_uRrc2XfY_rbN_gr[9]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gs[9]_net_1\);
    
    \b7_nYhI39s[4]\ : SLE
      port map(D => \b7_nYhI39s_lm[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b7_nYhI39se, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b7_nYhI39s[4]_net_1\);
    
    b10_nYhI3_umjB_1_RNO : CFG3
      generic map(INIT => x"01")

      port map(A => \b13_nAzGfFM_sLsv3[0]_net_1\, B => b6_nUT_fF, 
        C => N_71, Y => N_86);
    
    \b12_uRrc2XfY_rbN_5[8]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \b12_uRrc2XfY_rbN[9]_net_1\, B => 
        IICE_comm2iice(9), C => \b15_uRrc2XfY_rbN_gs[8]_net_1\, Y
         => \b12_uRrc2XfY_rbN_5[8]_net_1\);
    
    \b15_uRrc2XfY_rbN_gr[20]\ : SLE
      port map(D => \b7_nYhI39s[4]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gr[20]_net_1\);
    
    \b7_nYhI39s[9]\ : SLE
      port map(D => \b7_nYhI39s_lm[9]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b7_nYhI39se, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b7_nYhI39s[9]_net_1\);
    
    \b13_nAzGfFM_sLsv3_ns[1]\ : CFG3
      generic map(INIT => x"F2")

      port map(A => \b13_nAzGfFM_sLsv3[1]_net_1\, B => N_74, C
         => \b13_nAzGfFM_sLsv3[0]_net_1\, Y => 
        \b13_nAzGfFM_sLsv3_ns[1]_net_1\);
    
    \b12_uRrc2XfY_rbN[15]\ : SLE
      port map(D => \b12_uRrc2XfY_rbN_5[15]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \un1_b12_uRrc2XfY_rbN10_i\, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b12_uRrc2XfY_rbN[15]_net_1\);
    
    \b12_uRrc2XfY_rbN_5[11]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \b12_uRrc2XfY_rbN[12]_net_1\, B => 
        IICE_comm2iice(9), C => \b15_uRrc2XfY_rbN_gs[11]_net_1\, 
        Y => \b12_uRrc2XfY_rbN_5[11]_net_1\);
    
    b6_nUT_fF9 : CFG4
      generic map(INIT => x"AAA8")

      port map(A => \b8_vABZ3qsY\, B => \b3_nfs[0]_net_1\, C => 
        \b3_nfs[2]_net_1\, D => N_63_2, Y => N_61);
    
    \b15_uRrc2XfY_rbN_gr[10]\ : SLE
      port map(D => \b6_nfs_IF[4]\, CLK => IICE_comm2iice(11), EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b15_uRrc2XfY_rbN_gr[10]_net_1\);
    
    \b7_nYhI39s_cry[6]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \b7_nYhI39s[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \b7_nYhI39s_cry[5]_net_1\, S => \b7_nYhI39s_s[6]\, Y => 
        OPEN, FCO => \b7_nYhI39s_cry[6]_net_1\);
    
    b10_nYhI3_umjB_2 : SLE
      port map(D => \b10_nYhI3_umjB_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => b10_nYhI3_umjB);
    
    b6_Ocm0rW7 : CFG3
      generic map(INIT => x"01")

      port map(A => \b3_nfs[2]_net_1\, B => N_63_2, C => 
        \b3_nfs[1]_net_1\, Y => N_62);
    
    \b7_nYhI39s_cry[9]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \b7_nYhI39s[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \b7_nYhI39s_cry[8]_net_1\, S => \b7_nYhI39s_s[9]\, Y => 
        OPEN, FCO => \b7_nYhI39s_cry[9]_net_1\);
    
    \b13_nAzGfFM_sLsv3_ns_o3[3]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => b13_wRBtT_ME83hHx, B => 
        \b13_nAzGfFM_sLsv3[2]_net_1\, C => 
        \b13_nAzGfFM_sLsv3[3]_net_1\, Y => N_140);
    
    \b13_nAzGfFM_sLsv3_ns[4]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \b13_nAzGfFM_sLsv3[4]_net_1\, B => 
        b10_nYhI3_umjB, C => N_140, Y => 
        \b13_nAzGfFM_sLsv3_ns[4]_net_1\);
    
    \b15_uRrc2XfY_rbN_gs[26]\ : SLE
      port map(D => \b15_uRrc2XfY_rbN_gr[26]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gs[26]_net_1\);
    
    \b12_uRrc2XfY_rbN_5[15]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \b12_uRrc2XfY_rbN[16]_net_1\, B => 
        IICE_comm2iice(9), C => \b15_uRrc2XfY_rbN_gs[15]_net_1\, 
        Y => \b12_uRrc2XfY_rbN_5[15]_net_1\);
    
    \b12_uRrc2XfY_rbN_5[27]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \b15_uRrc2XfY_rbN_gs[27]_net_1\, B => 
        IICE_comm2iice(7), C => IICE_comm2iice(9), Y => 
        \b12_uRrc2XfY_rbN_5[27]_net_1\);
    
    \b12_uRrc2XfY_rbN_5[10]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \b12_uRrc2XfY_rbN[11]_net_1\, B => 
        IICE_comm2iice(9), C => \b15_uRrc2XfY_rbN_gs[10]_net_1\, 
        Y => \b12_uRrc2XfY_rbN_5[10]_net_1\);
    
    b12_voSc3_gmasbb_RNI0GM6_0 : CFG1
      generic map(INIT => "01")

      port map(A => \b5_voSc3\, Y => b5_voSc3_i);
    
    \b12_uRrc2XfY_rbN_5[0]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \b12_uRrc2XfY_rbN[1]_net_1\, B => 
        IICE_comm2iice(9), C => \b15_uRrc2XfY_rbN_gs[0]_net_1\, Y
         => \b12_uRrc2XfY_rbN_5[0]_net_1\);
    
    \b13_nAzGfFM_sLsv3[5]\ : SLE
      port map(D => \b13_nAzGfFM_sLsv3_ns[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        \b6_nfs_IF_i[1]\, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \b13_nAzGfFM_sLsv3[5]_net_1\);
    
    \b15_uRrc2XfY_rbN_gs[21]\ : SLE
      port map(D => \b15_uRrc2XfY_rbN_gr[21]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gs[21]_net_1\);
    
    \b15_uRrc2XfY_rbN_gs[0]\ : SLE
      port map(D => \b15_uRrc2XfY_rbN_gr[0]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gs[0]_net_1\);
    
    \b12_uRrc2XfY_rbN_5[18]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \b12_uRrc2XfY_rbN[19]_net_1\, B => 
        IICE_comm2iice(9), C => \b15_uRrc2XfY_rbN_gs[18]_net_1\, 
        Y => \b12_uRrc2XfY_rbN_5[18]_net_1\);
    
    \b15_uRrc2XfY_rbN_gr[7]\ : SLE
      port map(D => \b6_nfs_IF[1]\, CLK => IICE_comm2iice(11), EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b15_uRrc2XfY_rbN_gr[7]_net_1\);
    
    \b6_Ocm0rW_0[2]\ : CFG4
      generic map(INIT => x"FEFA")

      port map(A => \b13_nAzGfFM_sLsv3[3]_net_1\, B => 
        \b13_nAzGfFM_sLsv3[1]_net_1\, C => 
        \b13_nAzGfFM_sLsv3[2]_net_1\, D => N_74, Y => 
        \b6_Ocm0rW[2]\);
    
    \b15_uRrc2XfY_rbN_gs[8]\ : SLE
      port map(D => \b15_uRrc2XfY_rbN_gr[8]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gs[8]_net_1\);
    
    iclksync : clock2_en_reg_en_5s_x_0
      port map(status_b2sclk(3) => \status_b2sclk[3]\, 
        status_b2sclk(2) => \status_b2sclk[2]\, status_b2sclk(1)
         => \status_b2sclk[1]\, status_b2sclk(0) => 
        \status_b2sclk[0]\, b6_Ocm0rW(2) => \b6_Ocm0rW[2]\, 
        b6_Ocm0rW(1) => \b6_Ocm0rW[1]\, b6_Ocm0rW(0) => 
        \b6_Ocm0rW[0]\, b13_nAzGfFM_sLsv3_0 => 
        \b13_nAzGfFM_sLsv3[5]_net_1\, IICE_comm2iice_0 => 
        IICE_comm2iice(11), b6_nfs_IF_i_0 => \b6_nfs_IF_i[1]\, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0);
    
    \b3_nUT[10]\ : SLE
      port map(D => \b6_nUT_IF[10]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => \b6_nfs_IF_i[1]\, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b3_nUT[10]_net_1\);
    
    b12_voSc3_gmasbb : SLE
      port map(D => \b13_nAzGfFM_sLsv3[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b12_voSc3_gmasbb\);
    
    \b15_uRrc2XfY_rbN_gr[6]\ : SLE
      port map(D => \b6_nfs_IF[0]\, CLK => IICE_comm2iice(11), EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b15_uRrc2XfY_rbN_gr[6]_net_1\);
    
    \b15_uRrc2XfY_rbN_gr[27]\ : SLE
      port map(D => \b7_nYhI39s[11]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gr[27]_net_1\);
    
    \b12_uRrc2XfY_rbN[26]\ : SLE
      port map(D => \b12_uRrc2XfY_rbN_5[26]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \un1_b12_uRrc2XfY_rbN10_i\, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b12_uRrc2XfY_rbN[26]_net_1\);
    
    \b3_nUT[9]\ : SLE
      port map(D => \b6_nUT_IF[9]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => \b6_nfs_IF_i[1]\, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b3_nUT[9]_net_1\);
    
    \b15_uRrc2XfY_rbN_gr[19]\ : SLE
      port map(D => \b7_nYhI39s[3]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gr[19]_net_1\);
    
    \un13[2]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \b13_nAzGfFM_sLsv3[4]_net_1\, B => 
        \b13_nAzGfFM_sLsv3[5]_net_1\, Y => \un13[2]_net_1\);
    
    \b15_uRrc2XfY_rbN_gr[24]\ : SLE
      port map(D => \b7_nYhI39s[8]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gr[24]_net_1\);
    
    \b7_nYhI39s_lm_0[4]\ : CFG4
      generic map(INIT => x"AAC0")

      port map(A => \b7_nYhI39s_s[4]\, B => \b3_nUT[4]_net_1\, C
         => N_71, D => b6_nUT_fF, Y => \b7_nYhI39s_lm[4]\);
    
    \b7_nYhI39s[0]\ : SLE
      port map(D => \b7_nYhI39s_lm[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b7_nYhI39se, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b7_nYhI39s[0]_net_1\);
    
    \b12_uRrc2XfY_rbN[5]\ : SLE
      port map(D => \b12_uRrc2XfY_rbN_5[5]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \un1_b12_uRrc2XfY_rbN10_i\, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b12_uRrc2XfY_rbN[5]_net_1\);
    
    \b12_uRrc2XfY_rbN[18]\ : SLE
      port map(D => \b12_uRrc2XfY_rbN_5[18]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \un1_b12_uRrc2XfY_rbN10_i\, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b12_uRrc2XfY_rbN[18]_net_1\);
    
    \b7_nYhI39s[11]\ : SLE
      port map(D => \b7_nYhI39s_lm[11]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b7_nYhI39se, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b7_nYhI39s[11]_net_1\);
    
    \b15_uRrc2XfY_rbN_gs[16]\ : SLE
      port map(D => \b15_uRrc2XfY_rbN_gr[16]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gs[16]_net_1\);
    
    \b6_Ocm0rW_0[1]\ : CFG4
      generic map(INIT => x"DCFC")

      port map(A => b10_nYhI3_umjB, B => 
        \b13_nAzGfFM_sLsv3[4]_net_1\, C => N_324, D => N_62, Y
         => \b6_Ocm0rW[1]\);
    
    \b12_uRrc2XfY_rbN_5[7]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \b12_uRrc2XfY_rbN[8]_net_1\, B => 
        IICE_comm2iice(9), C => \b15_uRrc2XfY_rbN_gs[7]_net_1\, Y
         => \b12_uRrc2XfY_rbN_5[7]_net_1\);
    
    \b12_uRrc2XfY_rbN[3]\ : SLE
      port map(D => \b12_uRrc2XfY_rbN_5[3]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \un1_b12_uRrc2XfY_rbN10_i\, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b12_uRrc2XfY_rbN[3]_net_1\);
    
    \b12_uRrc2XfY_rbN[27]\ : SLE
      port map(D => \b12_uRrc2XfY_rbN_5[27]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \un1_b12_uRrc2XfY_rbN10_i\, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b12_uRrc2XfY_rbN[27]_net_1\);
    
    \b15_uRrc2XfY_rbN_gr[17]\ : SLE
      port map(D => \b7_nYhI39s[1]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gr[17]_net_1\);
    
    \b7_nYhI39s[2]\ : SLE
      port map(D => \b7_nYhI39s_lm[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b7_nYhI39se, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b7_nYhI39s[2]_net_1\);
    
    \b15_uRrc2XfY_rbN_gs[2]\ : SLE
      port map(D => \b15_uRrc2XfY_rbN_gr[2]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gs[2]_net_1\);
    
    \b7_nYhI39s[8]\ : SLE
      port map(D => \b7_nYhI39s_lm[8]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b7_nYhI39se, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b7_nYhI39s[8]_net_1\);
    
    \b7_nYhI39s_cry[1]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \b7_nYhI39s[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \b7_nYhI39s_cry[0]_net_1\, S => \b7_nYhI39s_s[1]\, Y => 
        OPEN, FCO => \b7_nYhI39s_cry[1]_net_1\);
    
    \b15_uRrc2XfY_rbN_gs[11]\ : SLE
      port map(D => \b15_uRrc2XfY_rbN_gr[11]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gs[11]_net_1\);
    
    \b15_uRrc2XfY_rbN_gr[14]\ : SLE
      port map(D => \b13_nAzGfFM_sLsv3[5]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gr[14]_net_1\);
    
    \b15_uRrc2XfY_rbN_gs[3]\ : SLE
      port map(D => \b15_uRrc2XfY_rbN_gr[3]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gs[3]_net_1\);
    
    \b3_nUT[5]\ : SLE
      port map(D => \b6_nUT_IF[5]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => \b6_nfs_IF_i[1]\, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b3_nUT[5]_net_1\);
    
    \b12_uRrc2XfY_rbN[22]\ : SLE
      port map(D => \b12_uRrc2XfY_rbN_5[22]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \un1_b12_uRrc2XfY_rbN10_i\, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b12_uRrc2XfY_rbN[22]_net_1\);
    
    \b3_nfs[4]\ : SLE
      port map(D => \b6_nfs_IF[4]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b3_nfs[4]_net_1\);
    
    \b15_uRrc2XfY_rbN_gr[8]\ : SLE
      port map(D => \b6_nfs_IF[2]\, CLK => IICE_comm2iice(11), EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b15_uRrc2XfY_rbN_gr[8]_net_1\);
    
    \b12_uRrc2XfY_rbN_5[3]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \b12_uRrc2XfY_rbN[4]_net_1\, B => 
        IICE_comm2iice(9), C => \b15_uRrc2XfY_rbN_gs[3]_net_1\, Y
         => \b12_uRrc2XfY_rbN_5[3]_net_1\);
    
    \b13_nAzGfFM_sLsv3_RNIO4SI[3]\ : CFG3
      generic map(INIT => x"1D")

      port map(A => \b13_nAzGfFM_sLsv3[1]_net_1\, B => 
        \b13_nAzGfFM_sLsv3[3]_net_1\, C => b10_nYhI3_umjB, Y => 
        b7_nYhI39slde_1_0);
    
    \b3_nfs[2]\ : SLE
      port map(D => \b6_nfs_IF[2]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b3_nfs[2]_net_1\);
    
    \b15_uRrc2XfY_rbN_gr[25]\ : SLE
      port map(D => \b7_nYhI39s[9]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gr[25]_net_1\);
    
    \b3_nUT[8]\ : SLE
      port map(D => \b6_nUT_IF[8]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => \b6_nfs_IF_i[1]\, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b3_nUT[8]_net_1\);
    
    \b12_uRrc2XfY_rbN[20]\ : SLE
      port map(D => \b12_uRrc2XfY_rbN_5[20]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \un1_b12_uRrc2XfY_rbN10_i\, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b12_uRrc2XfY_rbN[20]_net_1\);
    
    \b12_uRrc2XfY_rbN[9]\ : SLE
      port map(D => \b12_uRrc2XfY_rbN_5[9]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \un1_b12_uRrc2XfY_rbN10_i\, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b12_uRrc2XfY_rbN[9]_net_1\);
    
    \b7_nYhI39s_lm_0[8]\ : CFG4
      generic map(INIT => x"AAC0")

      port map(A => \b7_nYhI39s_s[8]\, B => \b3_nUT[8]_net_1\, C
         => N_71, D => b6_nUT_fF, Y => \b7_nYhI39s_lm[8]\);
    
    \b15_uRrc2XfY_rbN_gs[23]\ : SLE
      port map(D => \b15_uRrc2XfY_rbN_gr[23]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gs[23]_net_1\);
    
    \b6_Ocm0rW_0[0]\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_324, B => \b13_nAzGfFM_sLsv3[2]_net_1\, Y
         => \b6_Ocm0rW[0]\);
    
    b6_nUT_fF_0 : CFG4
      generic map(INIT => x"BAAA")

      port map(A => \b13_nAzGfFM_sLsv3[3]_net_1\, B => 
        b10_nYhI3_umjB, C => \b13_nAzGfFM_sLsv3[1]_net_1\, D => 
        N_61, Y => b6_nUT_fF);
    
    \b12_uRrc2XfY_rbN_5[16]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \b12_uRrc2XfY_rbN[17]_net_1\, B => 
        IICE_comm2iice(9), C => \b15_uRrc2XfY_rbN_gs[16]_net_1\, 
        Y => \b12_uRrc2XfY_rbN_5[16]_net_1\);
    
    \b15_uRrc2XfY_rbN_gr[15]\ : SLE
      port map(D => b11_vABZ3qsY_qH, CLK => IICE_comm2iice(11), 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b15_uRrc2XfY_rbN_gr[15]_net_1\);
    
    \b13_nAzGfFM_sLsv3[4]\ : SLE
      port map(D => \b13_nAzGfFM_sLsv3_ns[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        \b6_nfs_IF_i[1]\, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \b13_nAzGfFM_sLsv3[4]_net_1\);
    
    \b12_uRrc2XfY_rbN[2]\ : SLE
      port map(D => \b12_uRrc2XfY_rbN_5[2]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \un1_b12_uRrc2XfY_rbN10_i\, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b12_uRrc2XfY_rbN[2]_net_1\);
    
    \b7_nYhI39s_cry[3]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \b7_nYhI39s[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \b7_nYhI39s_cry[2]_net_1\, S => \b7_nYhI39s_s[3]\, Y => 
        OPEN, FCO => \b7_nYhI39s_cry[3]_net_1\);
    
    \b6_Ocm0rW_0_a2[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_61, B => \b13_nAzGfFM_sLsv3[1]_net_1\, Y
         => N_324);
    
    \b3_nUT[7]\ : SLE
      port map(D => \b6_nUT_IF[7]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => \b6_nfs_IF_i[1]\, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b3_nUT[7]_net_1\);
    
    \b15_uRrc2XfY_rbN_gs[18]\ : SLE
      port map(D => \b15_uRrc2XfY_rbN_gr[18]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gs[18]_net_1\);
    
    \b12_uRrc2XfY_rbN_5[19]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \b12_uRrc2XfY_rbN[20]_net_1\, B => 
        IICE_comm2iice(9), C => \b15_uRrc2XfY_rbN_gs[19]_net_1\, 
        Y => \b12_uRrc2XfY_rbN_5[19]_net_1\);
    
    b10_nYhI3_umjB_0_sqmuxa_7 : CFG4
      generic map(INIT => x"0100")

      port map(A => \b7_nYhI39s[10]_net_1\, B => 
        \b7_nYhI39s[9]_net_1\, C => \b7_nYhI39s[1]_net_1\, D => 
        \b7_nYhI39s[0]_net_1\, Y => \b10_nYhI3_umjB_0_sqmuxa_7\);
    
    \b7_nYhI39s_cry[0]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \b7_nYhI39s[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => GND_net_1, S => OPEN, Y
         => \b7_nYhI39s_cry_Y[0]\, FCO => 
        \b7_nYhI39s_cry[0]_net_1\);
    
    \b12_uRrc2XfY_rbN[21]\ : SLE
      port map(D => \b12_uRrc2XfY_rbN_5[21]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \un1_b12_uRrc2XfY_rbN10_i\, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b12_uRrc2XfY_rbN[21]_net_1\);
    
    \b12_uRrc2XfY_rbN_5[13]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \b12_uRrc2XfY_rbN[14]_net_1\, B => 
        IICE_comm2iice(9), C => \b15_uRrc2XfY_rbN_gs[13]_net_1\, 
        Y => \b12_uRrc2XfY_rbN_5[13]_net_1\);
    
    \b7_nYhI39s_lm_0[3]\ : CFG4
      generic map(INIT => x"AAC0")

      port map(A => \b7_nYhI39s_s[3]\, B => \b3_nUT[3]_net_1\, C
         => N_71, D => b6_nUT_fF, Y => \b7_nYhI39s_lm[3]\);
    
    b10_xoU0_WMrtX_0_sqmuxa_1_0_a3 : CFG2
      generic map(INIT => x"8")

      port map(A => N_74, B => \b13_nAzGfFM_sLsv3[1]_net_1\, Y
         => b10_xoU0_WMrtX_0_sqmuxa_1);
    
    \b13_nAzGfFM_sLsv3_ns[5]\ : CFG4
      generic map(INIT => x"AAEA")

      port map(A => \b13_nAzGfFM_sLsv3[5]_net_1\, B => 
        \b13_nAzGfFM_sLsv3[2]_net_1\, C => \b3_nfs[4]_net_1\, D
         => b13_wRBtT_ME83hHx, Y => 
        \b13_nAzGfFM_sLsv3_ns[5]_net_1\);
    
    \b12_uRrc2XfY_rbN_5[14]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \b12_uRrc2XfY_rbN[15]_net_1\, B => 
        IICE_comm2iice(9), C => \b15_uRrc2XfY_rbN_gs[14]_net_1\, 
        Y => \b12_uRrc2XfY_rbN_5[14]_net_1\);
    
    b10_nYhI3_umjB_1 : CFG4
      generic map(INIT => x"00E2")

      port map(A => \b10_nYhI3_umjB_0_sqmuxa\, B => N_86, C => 
        b10_nYhI3_umjB, D => N_71, Y => \b10_nYhI3_umjB_1\);
    
    \b15_uRrc2XfY_rbN_gs[13]\ : SLE
      port map(D => \b15_uRrc2XfY_rbN_gr[13]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gs[13]_net_1\);
    
    \b7_nYhI39s_lm_0[1]\ : CFG4
      generic map(INIT => x"AACF")

      port map(A => \b7_nYhI39s_s[1]\, B => \b3_nUT[1]_net_1\, C
         => N_71, D => b6_nUT_fF, Y => \b7_nYhI39s_lm[1]\);
    
    \b7_nYhI39s_lm_0[10]\ : CFG4
      generic map(INIT => x"AAC0")

      port map(A => \b7_nYhI39s_s[10]\, B => \b3_nUT[10]_net_1\, 
        C => N_71, D => b6_nUT_fF, Y => \b7_nYhI39s_lm[10]\);
    
    \b12_uRrc2XfY_rbN[16]\ : SLE
      port map(D => \b12_uRrc2XfY_rbN_5[16]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \un1_b12_uRrc2XfY_rbN10_i\, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b12_uRrc2XfY_rbN[16]_net_1\);
    
    \b15_uRrc2XfY_rbN_gr[1]\ : SLE
      port map(D => \status_b2sclk[1]\, CLK => IICE_comm2iice(11), 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b15_uRrc2XfY_rbN_gr[1]_net_1\);
    
    \b7_nYhI39s_lm_0[7]\ : CFG4
      generic map(INIT => x"AAC0")

      port map(A => \b7_nYhI39s_s[7]\, B => \b3_nUT[7]_net_1\, C
         => N_71, D => b6_nUT_fF, Y => \b7_nYhI39s_lm[7]\);
    
    \b12_uRrc2XfY_rbN_5[5]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \b12_uRrc2XfY_rbN[6]_net_1\, B => 
        IICE_comm2iice(9), C => \b15_uRrc2XfY_rbN_gs[5]_net_1\, Y
         => \b12_uRrc2XfY_rbN_5[5]_net_1\);
    
    \b12_uRrc2XfY_rbN_5[21]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \b12_uRrc2XfY_rbN[22]_net_1\, B => 
        IICE_comm2iice(9), C => \b15_uRrc2XfY_rbN_gs[21]_net_1\, 
        Y => \b12_uRrc2XfY_rbN_5[21]_net_1\);
    
    \b12_uRrc2XfY_rbN[17]\ : SLE
      port map(D => \b12_uRrc2XfY_rbN_5[17]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \un1_b12_uRrc2XfY_rbN10_i\, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b12_uRrc2XfY_rbN[17]_net_1\);
    
    b8_vABZ3qsY : SLE
      port map(D => b11_vABZ3qsY_qH, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b8_vABZ3qsY\);
    
    \b12_uRrc2XfY_rbN[24]\ : SLE
      port map(D => \b12_uRrc2XfY_rbN_5[24]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \un1_b12_uRrc2XfY_rbN10_i\, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b12_uRrc2XfY_rbN[24]_net_1\);
    
    \b7_nYhI39s_cry[4]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \b7_nYhI39s[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \b7_nYhI39s_cry[3]_net_1\, S => \b7_nYhI39s_s[4]\, Y => 
        OPEN, FCO => \b7_nYhI39s_cry[4]_net_1\);
    
    \b12_uRrc2XfY_rbN_5[9]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \b12_uRrc2XfY_rbN[10]_net_1\, B => 
        IICE_comm2iice(9), C => \b15_uRrc2XfY_rbN_gs[9]_net_1\, Y
         => \b12_uRrc2XfY_rbN_5[9]_net_1\);
    
    \b12_uRrc2XfY_rbN[23]\ : SLE
      port map(D => \b12_uRrc2XfY_rbN_5[23]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \un1_b12_uRrc2XfY_rbN10_i\, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b12_uRrc2XfY_rbN[23]_net_1\);
    
    \b15_uRrc2XfY_rbN_gs[22]\ : SLE
      port map(D => \b15_uRrc2XfY_rbN_gr[22]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gs[22]_net_1\);
    
    \b12_uRrc2XfY_rbN[12]\ : SLE
      port map(D => \b12_uRrc2XfY_rbN_5[12]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \un1_b12_uRrc2XfY_rbN10_i\, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b12_uRrc2XfY_rbN[12]_net_1\);
    
    \b7_nYhI39s_lm_0[11]\ : CFG4
      generic map(INIT => x"AAC0")

      port map(A => \b7_nYhI39s_s[11]_net_1\, B => 
        \b3_nUT[11]_net_1\, C => N_71, D => b6_nUT_fF, Y => 
        \b7_nYhI39s_lm[11]\);
    
    \b13_nAzGfFM_sLsv3[2]\ : SLE
      port map(D => \b13_nAzGfFM_sLsv3_ns[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        \b6_nfs_IF_i[1]\, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \b13_nAzGfFM_sLsv3[2]_net_1\);
    
    \b12_uRrc2XfY_rbN_5[25]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \b12_uRrc2XfY_rbN[26]_net_1\, B => 
        IICE_comm2iice(9), C => \b15_uRrc2XfY_rbN_gs[25]_net_1\, 
        Y => \b12_uRrc2XfY_rbN_5[25]_net_1\);
    
    \b12_uRrc2XfY_rbN_5[20]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \b12_uRrc2XfY_rbN[21]_net_1\, B => 
        IICE_comm2iice(9), C => \b15_uRrc2XfY_rbN_gs[20]_net_1\, 
        Y => \b12_uRrc2XfY_rbN_5[20]_net_1\);
    
    \b7_nYhI39s[10]\ : SLE
      port map(D => \b7_nYhI39s_lm[10]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b7_nYhI39se, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b7_nYhI39s[10]_net_1\);
    
    \b12_uRrc2XfY_rbN_5[12]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \b12_uRrc2XfY_rbN[13]_net_1\, B => 
        IICE_comm2iice(9), C => \b15_uRrc2XfY_rbN_gs[12]_net_1\, 
        Y => \b12_uRrc2XfY_rbN_5[12]_net_1\);
    
    \b3_nUT[2]\ : SLE
      port map(D => \b6_nUT_IF[2]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => \b6_nfs_IF_i[1]\, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b3_nUT[2]_net_1\);
    
    \b15_uRrc2XfY_rbN_gr[26]\ : SLE
      port map(D => \b7_nYhI39s[10]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gr[26]_net_1\);
    
    \b3_nfs_RNIJV7V[3]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \b3_nfs[4]_net_1\, B => \b3_nfs[3]_net_1\, Y
         => N_63_2);
    
    \b12_uRrc2XfY_rbN[10]\ : SLE
      port map(D => \b12_uRrc2XfY_rbN_5[10]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \un1_b12_uRrc2XfY_rbN10_i\, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b12_uRrc2XfY_rbN[10]_net_1\);
    
    \b15_uRrc2XfY_rbN_gr[9]\ : SLE
      port map(D => \b6_nfs_IF[3]\, CLK => IICE_comm2iice(11), EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b15_uRrc2XfY_rbN_gr[9]_net_1\);
    
    \b13_nAzGfFM_sLsv3_RNIMCCQ[0]\ : CFG4
      generic map(INIT => x"E5E4")

      port map(A => \b13_nAzGfFM_sLsv3[3]_net_1\, B => 
        \b13_nAzGfFM_sLsv3[0]_net_1\, C => b7_nYhI39slde_1_0, D
         => N_61, Y => b7_nYhI39se);
    
    \b12_uRrc2XfY_rbN_5[4]\ : CFG2
      generic map(INIT => x"4")

      port map(A => IICE_comm2iice(9), B => 
        \b12_uRrc2XfY_rbN[5]_net_1\, Y => 
        \b12_uRrc2XfY_rbN_5[4]_net_1\);
    
    \b3_nfs[3]\ : SLE
      port map(D => \b6_nfs_IF[3]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b3_nfs[3]_net_1\);
    
    \b15_uRrc2XfY_rbN_gr[21]\ : SLE
      port map(D => \b7_nYhI39s[5]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gr[21]_net_1\);
    
    \b12_uRrc2XfY_rbN[7]\ : SLE
      port map(D => \b12_uRrc2XfY_rbN_5[7]_net_1\, CLK => 
        IICE_comm2iice(11), EN => \un1_b12_uRrc2XfY_rbN10_i\, ALn
         => VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \b12_uRrc2XfY_rbN[7]_net_1\);
    
    \b13_nAzGfFM_sLsv3[3]\ : SLE
      port map(D => \b13_nAzGfFM_sLsv3_ns[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        \b6_nfs_IF_i[1]\, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \b13_nAzGfFM_sLsv3[3]_net_1\);
    
    \b7_nYhI39s[1]\ : SLE
      port map(D => \b7_nYhI39s_lm[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b7_nYhI39se, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b7_nYhI39s[1]_net_1\);
    
    \b15_uRrc2XfY_rbN_gs[20]\ : SLE
      port map(D => \b15_uRrc2XfY_rbN_gr[20]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gs[20]_net_1\);
    
    \b15_uRrc2XfY_rbN_gr[16]\ : SLE
      port map(D => \b7_nYhI39s[0]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gr[16]_net_1\);
    
    \b7_nYhI39s[7]\ : SLE
      port map(D => \b7_nYhI39s_lm[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => b7_nYhI39se, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b7_nYhI39s[7]_net_1\);
    
    \b13_nAzGfFM_sLsv3_ns[2]\ : CFG4
      generic map(INIT => x"CCCE")

      port map(A => \b13_nAzGfFM_sLsv3[2]_net_1\, B => 
        b10_xoU0_WMrtX_0_sqmuxa_1, C => \b3_nfs[4]_net_1\, D => 
        b13_wRBtT_ME83hHx, Y => \b13_nAzGfFM_sLsv3_ns[2]_net_1\);
    
    \b15_uRrc2XfY_rbN_gs[7]\ : SLE
      port map(D => \b15_uRrc2XfY_rbN_gr[7]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gs[7]_net_1\);
    
    \b7_nYhI39s_lm_0[9]\ : CFG4
      generic map(INIT => x"AAC0")

      port map(A => \b7_nYhI39s_s[9]\, B => \b3_nUT[9]_net_1\, C
         => N_71, D => b6_nUT_fF, Y => \b7_nYhI39s_lm[9]\);
    
    \b3_nUT[4]\ : SLE
      port map(D => \b6_nUT_IF[4]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => \b6_nfs_IF_i[1]\, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b3_nUT[4]_net_1\);
    
    \b7_nYhI39s_cry[7]\ : ARI1
      generic map(INIT => x"65500")

      port map(A => VCC_net_1, B => \b7_nYhI39s[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \b7_nYhI39s_cry[6]_net_1\, S => \b7_nYhI39s_s[7]\, Y => 
        OPEN, FCO => \b7_nYhI39s_cry[7]_net_1\);
    
    \b15_uRrc2XfY_rbN_gr[5]\ : SLE
      port map(D => \b13_nAzGfFM_sLsv3[2]_net_1\, CLK => 
        IICE_comm2iice(11), EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b15_uRrc2XfY_rbN_gr[5]_net_1\);
    
    \b7_nYhI39s_lm_0[5]\ : CFG4
      generic map(INIT => x"AAC0")

      port map(A => \b7_nYhI39s_s[5]\, B => \b3_nUT[5]_net_1\, C
         => N_71, D => b6_nUT_fF, Y => \b7_nYhI39s_lm[5]\);
    
    \b15_uRrc2XfY_rbN_gr[2]\ : SLE
      port map(D => \status_b2sclk[2]\, CLK => IICE_comm2iice(11), 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b15_uRrc2XfY_rbN_gr[2]_net_1\);
    
    \b15_uRrc2XfY_rbN_gr[11]\ : SLE
      port map(D => N_144_i, CLK => IICE_comm2iice(11), EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b15_uRrc2XfY_rbN_gr[11]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity IICE_x is

    port( IICE_comm2iice                   : in    std_logic_vector(11 downto 0);
          up_EOP_del                       : in    std_logic_vector(5 downto 0);
          RX_FIFO_DIN                      : in    std_logic_vector(7 downto 0);
          RX_packet_depth                  : in    std_logic_vector(7 downto 0);
          RX_FIFO_DOUT                     : in    std_logic_vector(8 downto 0);
          un15                             : in    std_logic_vector(10 downto 0);
          ReadFIFO_Write_Ptr               : in    std_logic_vector(1 downto 0);
          RX_FIFO_DIN_pipe                 : in    std_logic_vector(8 downto 0);
          p2s_data                         : in    std_logic_vector(7 downto 0);
          packet_available_clear_reg       : in    std_logic_vector(2 downto 0);
          ReadFIFO_Read_Ptr                : in    std_logic_vector(1 downto 0);
          iRX_FIFO_UNDERRUN                : in    std_logic_vector(3 downto 0);
          int_reg                          : in    std_logic_vector(7 downto 1);
          iRX_FIFO_Empty                   : in    std_logic_vector(3 downto 0);
          iRX_FIFO_Full                    : in    std_logic_vector(3 downto 0);
          manches_in_dly                   : in    std_logic_vector(1 downto 0);
          CoreAPB3_0_APBmslave0_PWDATA     : in    std_logic_vector(7 downto 0);
          clkdiv                           : in    std_logic_vector(3 downto 0);
          CoreAPB3_0_APBmslave0_PADDR      : in    std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PRDATA     : in    std_logic_vector(7 downto 0);
          un6                              : in    std_logic_vector(5 downto 0);
          control_reg_0                    : in    std_logic;
          control_reg_2                    : in    std_logic;
          control_reg_3                    : in    std_logic;
          IICE_iice2comm                   : out   std_logic;
          iup_EOP                          : in    std_logic;
          m2s010_som_sb_0_GPIO_28_SW_RESET : in    std_logic;
          TX_FIFO_Full                     : in    std_logic;
          TX_FIFO_wr_en                    : in    std_logic;
          tx_packet_complt                 : in    std_logic;
          RX_packet_depth_status           : in    std_logic;
          RX_FIFO_Empty                    : in    std_logic;
          RX_FIFO_Full                     : in    std_logic;
          rx_FIFO_OVERFLOW_int             : in    std_logic;
          RX_FIFO_rd_en                    : in    std_logic;
          rx_FIFO_UNDERRUN_int             : in    std_logic;
          rx_packet_complt                 : in    std_logic;
          RESET                            : in    std_logic;
          rx_CRC_error_int                 : in    std_logic;
          rx_packet_avail_int              : in    std_logic;
          TX_FIFO_Empty                    : in    std_logic;
          CommsFPGA_CCC_0_LOCK             : in    std_logic;
          MANCH_OUT_P_c                    : in    std_logic;
          MANCHESTER_IN_c                  : in    std_logic;
          int_reg_clr                      : in    std_logic;
          irx_center_sample                : in    std_logic;
          TX_FIFO_RST                      : in    std_logic;
          rx_FIFO_rst_reg                  : in    std_logic;
          start_tx_FIFO                    : in    std_logic;
          internal_loopback                : in    std_logic;
          external_loopback                : in    std_logic;
          iNRZ_data                        : in    std_logic;
          CoreAPB3_0_APBmslave0_PWRITE     : in    std_logic;
          bd_reset                         : in    std_logic;
          m2s010_som_sb_0_POWER_ON_RESET_N : in    std_logic;
          block_int_until_rd               : in    std_logic;
          CoreAPB3_0_APBmslave0_PREADY     : in    std_logic;
          long_reset                       : in    std_logic;
          CommsFPGA_CCC_0_GL0              : in    std_logic
        );

end IICE_x;

architecture DEF_ARCH of IICE_x is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component b11_OFWNT9s_8tZ_Z3_x
    port( mdiclink_reg        : in    std_logic_vector(167 downto 0) := (others => 'U');
          b11_OFWNT9L_8tZ     : out   std_logic_vector(167 downto 0);
          IICE_comm2iice      : in    std_logic_vector(11 downto 0) := (others => 'U');
          N_145_i             : in    std_logic := 'U';
          N_1261_i            : out   std_logic;
          b5_voSc3            : in    std_logic := 'U';
          b9_OFWNT9_ab        : in    std_logic := 'U';
          b13_wRBtT_ME83hHx   : in    std_logic := 'U';
          b5_voSc3_i          : in    std_logic := 'U';
          b10_OFWNT9_Y2x      : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component b3_uKr_x
    port( b13_nvmFL_fx2rbuQ : in    std_logic_vector(6 downto 1) := (others => 'U');
          b11_uRrc_9urXBb   : in    std_logic := 'U';
          b3_PLy            : in    std_logic := 'U';
          b3_PLF            : out   std_logic;
          b7_PLy_PlM        : out   std_logic;
          b7_nUTQ_9u        : out   std_logic;
          b7_PSyi_9u        : out   std_logic;
          b9_OFWNT9_ab      : out   std_logic;
          b9_PbTt39_ab      : out   std_logic;
          b9_PKFoLX_ab      : out   std_logic;
          b9_vbTtJX_ab      : out   std_logic;
          b8_ubTt3_YG       : out   std_logic;
          b9_ibScJX_ab      : out   std_logic;
          b7_yYh0_9u        : out   std_logic;
          b8_nUTQ_XlK       : in    std_logic := 'U';
          b8_PSyi_XlK       : in    std_logic := 'U';
          b10_OFWNT9_Y2x    : in    std_logic := 'U';
          b10_PbTt39_Y2x    : in    std_logic := 'U';
          b10_PKFoLX_Y2x    : in    std_logic := 'U';
          b10_vbTtJX_Y2x    : in    std_logic := 'U';
          b9_ubTt3_Mxf      : in    std_logic := 'U';
          b10_ibScJX_Y2x    : in    std_logic := 'U';
          b8_yYh0_XlK       : in    std_logic := 'U'
        );
  end component;

  component b8_PfFzrNYI_x
    port( b11_OFWNT9L_8tZ     : in    std_logic_vector(167 downto 0) := (others => 'U');
          mdiclink_reg        : in    std_logic_vector(167 downto 0) := (others => 'U');
          IICE_comm2iice_4    : in    std_logic := 'U';
          IICE_comm2iice_0    : in    std_logic := 'U';
          IICE_comm2iice_3    : in    std_logic := 'U';
          b10_nYBzIXrKbK_0    : out   std_logic;
          b7_PSyi_9u          : in    std_logic := 'U';
          b12_PSyi_XlK_qHv    : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U'
        );
  end component;

  component b7_OCByLXC_Z1_x_0
    port( IICE_comm2iice      : in    std_logic_vector(11 downto 7) := (others => 'U');
          b9_PKFoLX_ab        : in    std_logic := 'U';
          b8_nUTQ_XlK         : out   std_logic;
          b7_nUTQ_9u          : in    std_logic := 'U';
          b10_PKFoLX_Y2x      : out   std_logic;
          b10_vbTtJX_Y2x      : out   std_logic;
          b9_vbTtJX_ab        : in    std_logic := 'U';
          b8_ubTt3_YG         : in    std_logic := 'U';
          N_145_i             : out   std_logic;
          b13_wRBtT_ME83hHx   : in    std_logic := 'U';
          b9_ubTt3_Mxf        : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          b5_voSc3_i          : out   std_logic;
          b5_voSc3            : out   std_logic
        );
  end component;

    signal \mdiclink_reg[10]_net_1\, VCC_net_1, GND_net_1, 
        \mdiclink_reg[9]_net_1\, \mdiclink_reg[8]_net_1\, 
        \mdiclink_reg[7]_net_1\, \mdiclink_reg[6]_net_1\, 
        \mdiclink_reg[5]_net_1\, \mdiclink_reg[4]_net_1\, 
        \mdiclink_reg[3]_net_1\, \mdiclink_reg[2]_net_1\, 
        \mdiclink_reg[1]_net_1\, \mdiclink_reg[0]_net_1\, 
        \mdiclink_reg[25]_net_1\, \mdiclink_reg[24]_net_1\, 
        \mdiclink_reg[23]_net_1\, \mdiclink_reg[22]_net_1\, 
        \mdiclink_reg[21]_net_1\, \mdiclink_reg[20]_net_1\, 
        \mdiclink_reg[19]_net_1\, \mdiclink_reg[18]_net_1\, 
        \mdiclink_reg[17]_net_1\, \mdiclink_reg[16]_net_1\, 
        \mdiclink_reg[15]_net_1\, \mdiclink_reg[14]_net_1\, 
        \mdiclink_reg[13]_net_1\, \mdiclink_reg[12]_net_1\, 
        \mdiclink_reg[11]_net_1\, \mdiclink_reg[40]_net_1\, 
        \mdiclink_reg[39]_net_1\, \mdiclink_reg[38]_net_1\, 
        \mdiclink_reg[37]_net_1\, \mdiclink_reg[36]_net_1\, 
        \mdiclink_reg[35]_net_1\, \mdiclink_reg[34]_net_1\, 
        \mdiclink_reg[33]_net_1\, \mdiclink_reg[32]_net_1\, 
        \mdiclink_reg[31]_net_1\, \mdiclink_reg[30]_net_1\, 
        \mdiclink_reg[29]_net_1\, \mdiclink_reg[28]_net_1\, 
        \mdiclink_reg[27]_net_1\, \mdiclink_reg[26]_net_1\, 
        \mdiclink_reg[55]_net_1\, \mdiclink_reg[54]_net_1\, 
        \mdiclink_reg[53]_net_1\, \mdiclink_reg[52]_net_1\, 
        \mdiclink_reg[51]_net_1\, \mdiclink_reg[50]_net_1\, 
        \mdiclink_reg[49]_net_1\, \mdiclink_reg[48]_net_1\, 
        \mdiclink_reg[47]_net_1\, \mdiclink_reg[46]_net_1\, 
        \mdiclink_reg[45]_net_1\, \mdiclink_reg[44]_net_1\, 
        \mdiclink_reg[43]_net_1\, \mdiclink_reg[42]_net_1\, 
        \mdiclink_reg[41]_net_1\, \mdiclink_reg[70]_net_1\, 
        \mdiclink_reg[69]_net_1\, \mdiclink_reg[68]_net_1\, 
        \mdiclink_reg[67]_net_1\, \mdiclink_reg[66]_net_1\, 
        \mdiclink_reg[65]_net_1\, \mdiclink_reg[64]_net_1\, 
        \mdiclink_reg[63]_net_1\, \mdiclink_reg[62]_net_1\, 
        \mdiclink_reg[61]_net_1\, \mdiclink_reg[60]_net_1\, 
        \mdiclink_reg[59]_net_1\, \mdiclink_reg[58]_net_1\, 
        \mdiclink_reg[57]_net_1\, \mdiclink_reg[56]_net_1\, 
        \mdiclink_reg[85]_net_1\, \mdiclink_reg[84]_net_1\, 
        \mdiclink_reg[83]_net_1\, \mdiclink_reg[82]_net_1\, 
        \mdiclink_reg[81]_net_1\, \mdiclink_reg[80]_net_1\, 
        \mdiclink_reg[79]_net_1\, \mdiclink_reg[78]_net_1\, 
        \mdiclink_reg[77]_net_1\, \mdiclink_reg[76]_net_1\, 
        \mdiclink_reg[75]_net_1\, \mdiclink_reg[74]_net_1\, 
        \mdiclink_reg[73]_net_1\, \mdiclink_reg[72]_net_1\, 
        \mdiclink_reg[71]_net_1\, \mdiclink_reg[100]_net_1\, 
        \mdiclink_reg[99]_net_1\, \mdiclink_reg[98]_net_1\, 
        \mdiclink_reg[97]_net_1\, \mdiclink_reg[96]_net_1\, 
        \mdiclink_reg[95]_net_1\, \mdiclink_reg[94]_net_1\, 
        \mdiclink_reg[93]_net_1\, \mdiclink_reg[92]_net_1\, 
        \mdiclink_reg[91]_net_1\, \mdiclink_reg[90]_net_1\, 
        \mdiclink_reg[89]_net_1\, \mdiclink_reg[88]_net_1\, 
        \mdiclink_reg[87]_net_1\, \mdiclink_reg[86]_net_1\, 
        \mdiclink_reg[115]_net_1\, \mdiclink_reg[114]_net_1\, 
        \mdiclink_reg[113]_net_1\, \mdiclink_reg[112]_net_1\, 
        \mdiclink_reg[111]_net_1\, \mdiclink_reg[110]_net_1\, 
        \mdiclink_reg[109]_net_1\, \mdiclink_reg[108]_net_1\, 
        \mdiclink_reg[107]_net_1\, \mdiclink_reg[106]_net_1\, 
        \mdiclink_reg[105]_net_1\, \mdiclink_reg[104]_net_1\, 
        \mdiclink_reg[103]_net_1\, \mdiclink_reg[102]_net_1\, 
        \mdiclink_reg[101]_net_1\, \mdiclink_reg[130]_net_1\, 
        \mdiclink_reg[129]_net_1\, \mdiclink_reg[128]_net_1\, 
        \mdiclink_reg[127]_net_1\, \mdiclink_reg[126]_net_1\, 
        \mdiclink_reg[125]_net_1\, \mdiclink_reg[124]_net_1\, 
        \mdiclink_reg[123]_net_1\, \mdiclink_reg[122]_net_1\, 
        \mdiclink_reg[121]_net_1\, \mdiclink_reg[120]_net_1\, 
        \mdiclink_reg[119]_net_1\, \mdiclink_reg[118]_net_1\, 
        \mdiclink_reg[117]_net_1\, \mdiclink_reg[116]_net_1\, 
        \mdiclink_reg[145]_net_1\, \mdiclink_reg[144]_net_1\, 
        \mdiclink_reg[143]_net_1\, \mdiclink_reg[142]_net_1\, 
        \mdiclink_reg[141]_net_1\, \mdiclink_reg[140]_net_1\, 
        \mdiclink_reg[139]_net_1\, \mdiclink_reg[138]_net_1\, 
        \mdiclink_reg[137]_net_1\, \mdiclink_reg[136]_net_1\, 
        \mdiclink_reg[135]_net_1\, \mdiclink_reg[134]_net_1\, 
        \mdiclink_reg[133]_net_1\, \mdiclink_reg[132]_net_1\, 
        \mdiclink_reg[131]_net_1\, \mdiclink_reg[160]_net_1\, 
        \mdiclink_reg[159]_net_1\, \mdiclink_reg[158]_net_1\, 
        \mdiclink_reg[157]_net_1\, \mdiclink_reg[156]_net_1\, 
        \mdiclink_reg[155]_net_1\, \mdiclink_reg[154]_net_1\, 
        \mdiclink_reg[153]_net_1\, \mdiclink_reg[152]_net_1\, 
        \mdiclink_reg[151]_net_1\, \mdiclink_reg[150]_net_1\, 
        \mdiclink_reg[149]_net_1\, \mdiclink_reg[148]_net_1\, 
        \mdiclink_reg[147]_net_1\, \mdiclink_reg[146]_net_1\, 
        \b13_wRBtT_ME83hHx\, \b10_nYBzIXrKbK[1]\, 
        \mdiclink_reg[167]_net_1\, \mdiclink_reg[166]_net_1\, 
        \mdiclink_reg[165]_net_1\, \mdiclink_reg[164]_net_1\, 
        \mdiclink_reg[163]_net_1\, \mdiclink_reg[162]_net_1\, 
        \mdiclink_reg[161]_net_1\, b4_PLyF, b7_nUTQ_9u, 
        b7_PSyi_9u, b9_OFWNT9_ab, b9_PbTt39_ab, b9_PKFoLX_ab, 
        b9_vbTtJX_ab, b8_ubTt3_YG, b9_ibScJX_ab, b7_yYh0_9u, 
        b8_nUTQ_XlK, b12_PSyi_XlK_qHv, b10_OFWNT9_Y2x, 
        b10_PKFoLX_Y2x, b10_vbTtJX_Y2x, b9_ubTt3_Mxf, N_1261_i, 
        N_145_i, b5_voSc3_i, b5_voSc3, \b11_OFWNT9L_8tZ[0]\, 
        \b11_OFWNT9L_8tZ[1]\, \b11_OFWNT9L_8tZ[2]\, 
        \b11_OFWNT9L_8tZ[3]\, \b11_OFWNT9L_8tZ[4]\, 
        \b11_OFWNT9L_8tZ[5]\, \b11_OFWNT9L_8tZ[6]\, 
        \b11_OFWNT9L_8tZ[7]\, \b11_OFWNT9L_8tZ[8]\, 
        \b11_OFWNT9L_8tZ[9]\, \b11_OFWNT9L_8tZ[10]\, 
        \b11_OFWNT9L_8tZ[11]\, \b11_OFWNT9L_8tZ[12]\, 
        \b11_OFWNT9L_8tZ[13]\, \b11_OFWNT9L_8tZ[14]\, 
        \b11_OFWNT9L_8tZ[15]\, \b11_OFWNT9L_8tZ[16]\, 
        \b11_OFWNT9L_8tZ[17]\, \b11_OFWNT9L_8tZ[18]\, 
        \b11_OFWNT9L_8tZ[19]\, \b11_OFWNT9L_8tZ[20]\, 
        \b11_OFWNT9L_8tZ[21]\, \b11_OFWNT9L_8tZ[22]\, 
        \b11_OFWNT9L_8tZ[23]\, \b11_OFWNT9L_8tZ[24]\, 
        \b11_OFWNT9L_8tZ[25]\, \b11_OFWNT9L_8tZ[26]\, 
        \b11_OFWNT9L_8tZ[27]\, \b11_OFWNT9L_8tZ[28]\, 
        \b11_OFWNT9L_8tZ[29]\, \b11_OFWNT9L_8tZ[30]\, 
        \b11_OFWNT9L_8tZ[31]\, \b11_OFWNT9L_8tZ[32]\, 
        \b11_OFWNT9L_8tZ[33]\, \b11_OFWNT9L_8tZ[34]\, 
        \b11_OFWNT9L_8tZ[35]\, \b11_OFWNT9L_8tZ[36]\, 
        \b11_OFWNT9L_8tZ[37]\, \b11_OFWNT9L_8tZ[38]\, 
        \b11_OFWNT9L_8tZ[39]\, \b11_OFWNT9L_8tZ[40]\, 
        \b11_OFWNT9L_8tZ[41]\, \b11_OFWNT9L_8tZ[42]\, 
        \b11_OFWNT9L_8tZ[43]\, \b11_OFWNT9L_8tZ[44]\, 
        \b11_OFWNT9L_8tZ[45]\, \b11_OFWNT9L_8tZ[46]\, 
        \b11_OFWNT9L_8tZ[47]\, \b11_OFWNT9L_8tZ[48]\, 
        \b11_OFWNT9L_8tZ[49]\, \b11_OFWNT9L_8tZ[50]\, 
        \b11_OFWNT9L_8tZ[51]\, \b11_OFWNT9L_8tZ[52]\, 
        \b11_OFWNT9L_8tZ[53]\, \b11_OFWNT9L_8tZ[54]\, 
        \b11_OFWNT9L_8tZ[55]\, \b11_OFWNT9L_8tZ[56]\, 
        \b11_OFWNT9L_8tZ[57]\, \b11_OFWNT9L_8tZ[58]\, 
        \b11_OFWNT9L_8tZ[59]\, \b11_OFWNT9L_8tZ[60]\, 
        \b11_OFWNT9L_8tZ[61]\, \b11_OFWNT9L_8tZ[62]\, 
        \b11_OFWNT9L_8tZ[63]\, \b11_OFWNT9L_8tZ[64]\, 
        \b11_OFWNT9L_8tZ[65]\, \b11_OFWNT9L_8tZ[66]\, 
        \b11_OFWNT9L_8tZ[67]\, \b11_OFWNT9L_8tZ[68]\, 
        \b11_OFWNT9L_8tZ[69]\, \b11_OFWNT9L_8tZ[70]\, 
        \b11_OFWNT9L_8tZ[71]\, \b11_OFWNT9L_8tZ[72]\, 
        \b11_OFWNT9L_8tZ[73]\, \b11_OFWNT9L_8tZ[74]\, 
        \b11_OFWNT9L_8tZ[75]\, \b11_OFWNT9L_8tZ[76]\, 
        \b11_OFWNT9L_8tZ[77]\, \b11_OFWNT9L_8tZ[78]\, 
        \b11_OFWNT9L_8tZ[79]\, \b11_OFWNT9L_8tZ[80]\, 
        \b11_OFWNT9L_8tZ[81]\, \b11_OFWNT9L_8tZ[82]\, 
        \b11_OFWNT9L_8tZ[83]\, \b11_OFWNT9L_8tZ[84]\, 
        \b11_OFWNT9L_8tZ[85]\, \b11_OFWNT9L_8tZ[86]\, 
        \b11_OFWNT9L_8tZ[87]\, \b11_OFWNT9L_8tZ[88]\, 
        \b11_OFWNT9L_8tZ[89]\, \b11_OFWNT9L_8tZ[90]\, 
        \b11_OFWNT9L_8tZ[91]\, \b11_OFWNT9L_8tZ[92]\, 
        \b11_OFWNT9L_8tZ[93]\, \b11_OFWNT9L_8tZ[94]\, 
        \b11_OFWNT9L_8tZ[95]\, \b11_OFWNT9L_8tZ[96]\, 
        \b11_OFWNT9L_8tZ[97]\, \b11_OFWNT9L_8tZ[98]\, 
        \b11_OFWNT9L_8tZ[99]\, \b11_OFWNT9L_8tZ[100]\, 
        \b11_OFWNT9L_8tZ[101]\, \b11_OFWNT9L_8tZ[102]\, 
        \b11_OFWNT9L_8tZ[103]\, \b11_OFWNT9L_8tZ[104]\, 
        \b11_OFWNT9L_8tZ[105]\, \b11_OFWNT9L_8tZ[106]\, 
        \b11_OFWNT9L_8tZ[107]\, \b11_OFWNT9L_8tZ[108]\, 
        \b11_OFWNT9L_8tZ[109]\, \b11_OFWNT9L_8tZ[110]\, 
        \b11_OFWNT9L_8tZ[111]\, \b11_OFWNT9L_8tZ[112]\, 
        \b11_OFWNT9L_8tZ[113]\, \b11_OFWNT9L_8tZ[114]\, 
        \b11_OFWNT9L_8tZ[115]\, \b11_OFWNT9L_8tZ[116]\, 
        \b11_OFWNT9L_8tZ[117]\, \b11_OFWNT9L_8tZ[118]\, 
        \b11_OFWNT9L_8tZ[119]\, \b11_OFWNT9L_8tZ[120]\, 
        \b11_OFWNT9L_8tZ[121]\, \b11_OFWNT9L_8tZ[122]\, 
        \b11_OFWNT9L_8tZ[123]\, \b11_OFWNT9L_8tZ[124]\, 
        \b11_OFWNT9L_8tZ[125]\, \b11_OFWNT9L_8tZ[126]\, 
        \b11_OFWNT9L_8tZ[127]\, \b11_OFWNT9L_8tZ[128]\, 
        \b11_OFWNT9L_8tZ[129]\, \b11_OFWNT9L_8tZ[130]\, 
        \b11_OFWNT9L_8tZ[131]\, \b11_OFWNT9L_8tZ[132]\, 
        \b11_OFWNT9L_8tZ[133]\, \b11_OFWNT9L_8tZ[134]\, 
        \b11_OFWNT9L_8tZ[135]\, \b11_OFWNT9L_8tZ[136]\, 
        \b11_OFWNT9L_8tZ[137]\, \b11_OFWNT9L_8tZ[138]\, 
        \b11_OFWNT9L_8tZ[139]\, \b11_OFWNT9L_8tZ[140]\, 
        \b11_OFWNT9L_8tZ[141]\, \b11_OFWNT9L_8tZ[142]\, 
        \b11_OFWNT9L_8tZ[143]\, \b11_OFWNT9L_8tZ[144]\, 
        \b11_OFWNT9L_8tZ[145]\, \b11_OFWNT9L_8tZ[146]\, 
        \b11_OFWNT9L_8tZ[147]\, \b11_OFWNT9L_8tZ[148]\, 
        \b11_OFWNT9L_8tZ[149]\, \b11_OFWNT9L_8tZ[150]\, 
        \b11_OFWNT9L_8tZ[151]\, \b11_OFWNT9L_8tZ[152]\, 
        \b11_OFWNT9L_8tZ[153]\, \b11_OFWNT9L_8tZ[154]\, 
        \b11_OFWNT9L_8tZ[155]\, \b11_OFWNT9L_8tZ[156]\, 
        \b11_OFWNT9L_8tZ[157]\, \b11_OFWNT9L_8tZ[158]\, 
        \b11_OFWNT9L_8tZ[159]\, \b11_OFWNT9L_8tZ[160]\, 
        \b11_OFWNT9L_8tZ[161]\, \b11_OFWNT9L_8tZ[162]\, 
        \b11_OFWNT9L_8tZ[163]\, \b11_OFWNT9L_8tZ[164]\, 
        \b11_OFWNT9L_8tZ[165]\, \b11_OFWNT9L_8tZ[166]\, 
        \b11_OFWNT9L_8tZ[167]\ : std_logic;
    signal nc2, nc1 : std_logic;

    for all : b11_OFWNT9s_8tZ_Z3_x
	Use entity work.b11_OFWNT9s_8tZ_Z3_x(DEF_ARCH);
    for all : b3_uKr_x
	Use entity work.b3_uKr_x(DEF_ARCH);
    for all : b8_PfFzrNYI_x
	Use entity work.b8_PfFzrNYI_x(DEF_ARCH);
    for all : b7_OCByLXC_Z1_x_0
	Use entity work.b7_OCByLXC_Z1_x_0(DEF_ARCH);
begin 


    \mdiclink_reg[162]\ : SLE
      port map(D => up_EOP_del(5), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[162]_net_1\);
    
    \mdiclink_reg[89]\ : SLE
      port map(D => packet_available_clear_reg(0), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[89]_net_1\);
    
    \mdiclink_reg[117]\ : SLE
      port map(D => RX_FIFO_DOUT(7), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[117]_net_1\);
    
    \mdiclink_reg[116]\ : SLE
      port map(D => RX_FIFO_DOUT(8), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[116]_net_1\);
    
    \mdiclink_reg[110]\ : SLE
      port map(D => RX_FIFO_DIN_pipe(5), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[110]_net_1\);
    
    \mdiclink_reg[90]\ : SLE
      port map(D => ReadFIFO_Read_Ptr(1), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[90]_net_1\);
    
    \mdiclink_reg[97]\ : SLE
      port map(D => un15(5), CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[97]_net_1\);
    
    \mdiclink_reg[108]\ : SLE
      port map(D => RX_FIFO_DIN_pipe(7), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[108]_net_1\);
    
    b3_SoW : b11_OFWNT9s_8tZ_Z3_x
      port map(mdiclink_reg(167) => \mdiclink_reg[167]_net_1\, 
        mdiclink_reg(166) => \mdiclink_reg[166]_net_1\, 
        mdiclink_reg(165) => \mdiclink_reg[165]_net_1\, 
        mdiclink_reg(164) => \mdiclink_reg[164]_net_1\, 
        mdiclink_reg(163) => \mdiclink_reg[163]_net_1\, 
        mdiclink_reg(162) => \mdiclink_reg[162]_net_1\, 
        mdiclink_reg(161) => \mdiclink_reg[161]_net_1\, 
        mdiclink_reg(160) => \mdiclink_reg[160]_net_1\, 
        mdiclink_reg(159) => \mdiclink_reg[159]_net_1\, 
        mdiclink_reg(158) => \mdiclink_reg[158]_net_1\, 
        mdiclink_reg(157) => \mdiclink_reg[157]_net_1\, 
        mdiclink_reg(156) => \mdiclink_reg[156]_net_1\, 
        mdiclink_reg(155) => \mdiclink_reg[155]_net_1\, 
        mdiclink_reg(154) => \mdiclink_reg[154]_net_1\, 
        mdiclink_reg(153) => \mdiclink_reg[153]_net_1\, 
        mdiclink_reg(152) => \mdiclink_reg[152]_net_1\, 
        mdiclink_reg(151) => \mdiclink_reg[151]_net_1\, 
        mdiclink_reg(150) => \mdiclink_reg[150]_net_1\, 
        mdiclink_reg(149) => \mdiclink_reg[149]_net_1\, 
        mdiclink_reg(148) => \mdiclink_reg[148]_net_1\, 
        mdiclink_reg(147) => \mdiclink_reg[147]_net_1\, 
        mdiclink_reg(146) => \mdiclink_reg[146]_net_1\, 
        mdiclink_reg(145) => \mdiclink_reg[145]_net_1\, 
        mdiclink_reg(144) => \mdiclink_reg[144]_net_1\, 
        mdiclink_reg(143) => \mdiclink_reg[143]_net_1\, 
        mdiclink_reg(142) => \mdiclink_reg[142]_net_1\, 
        mdiclink_reg(141) => \mdiclink_reg[141]_net_1\, 
        mdiclink_reg(140) => \mdiclink_reg[140]_net_1\, 
        mdiclink_reg(139) => \mdiclink_reg[139]_net_1\, 
        mdiclink_reg(138) => \mdiclink_reg[138]_net_1\, 
        mdiclink_reg(137) => \mdiclink_reg[137]_net_1\, 
        mdiclink_reg(136) => \mdiclink_reg[136]_net_1\, 
        mdiclink_reg(135) => \mdiclink_reg[135]_net_1\, 
        mdiclink_reg(134) => \mdiclink_reg[134]_net_1\, 
        mdiclink_reg(133) => \mdiclink_reg[133]_net_1\, 
        mdiclink_reg(132) => \mdiclink_reg[132]_net_1\, 
        mdiclink_reg(131) => \mdiclink_reg[131]_net_1\, 
        mdiclink_reg(130) => \mdiclink_reg[130]_net_1\, 
        mdiclink_reg(129) => \mdiclink_reg[129]_net_1\, 
        mdiclink_reg(128) => \mdiclink_reg[128]_net_1\, 
        mdiclink_reg(127) => \mdiclink_reg[127]_net_1\, 
        mdiclink_reg(126) => \mdiclink_reg[126]_net_1\, 
        mdiclink_reg(125) => \mdiclink_reg[125]_net_1\, 
        mdiclink_reg(124) => \mdiclink_reg[124]_net_1\, 
        mdiclink_reg(123) => \mdiclink_reg[123]_net_1\, 
        mdiclink_reg(122) => \mdiclink_reg[122]_net_1\, 
        mdiclink_reg(121) => \mdiclink_reg[121]_net_1\, 
        mdiclink_reg(120) => \mdiclink_reg[120]_net_1\, 
        mdiclink_reg(119) => \mdiclink_reg[119]_net_1\, 
        mdiclink_reg(118) => \mdiclink_reg[118]_net_1\, 
        mdiclink_reg(117) => \mdiclink_reg[117]_net_1\, 
        mdiclink_reg(116) => \mdiclink_reg[116]_net_1\, 
        mdiclink_reg(115) => \mdiclink_reg[115]_net_1\, 
        mdiclink_reg(114) => \mdiclink_reg[114]_net_1\, 
        mdiclink_reg(113) => \mdiclink_reg[113]_net_1\, 
        mdiclink_reg(112) => \mdiclink_reg[112]_net_1\, 
        mdiclink_reg(111) => \mdiclink_reg[111]_net_1\, 
        mdiclink_reg(110) => \mdiclink_reg[110]_net_1\, 
        mdiclink_reg(109) => \mdiclink_reg[109]_net_1\, 
        mdiclink_reg(108) => \mdiclink_reg[108]_net_1\, 
        mdiclink_reg(107) => \mdiclink_reg[107]_net_1\, 
        mdiclink_reg(106) => \mdiclink_reg[106]_net_1\, 
        mdiclink_reg(105) => \mdiclink_reg[105]_net_1\, 
        mdiclink_reg(104) => \mdiclink_reg[104]_net_1\, 
        mdiclink_reg(103) => \mdiclink_reg[103]_net_1\, 
        mdiclink_reg(102) => \mdiclink_reg[102]_net_1\, 
        mdiclink_reg(101) => \mdiclink_reg[101]_net_1\, 
        mdiclink_reg(100) => \mdiclink_reg[100]_net_1\, 
        mdiclink_reg(99) => \mdiclink_reg[99]_net_1\, 
        mdiclink_reg(98) => \mdiclink_reg[98]_net_1\, 
        mdiclink_reg(97) => \mdiclink_reg[97]_net_1\, 
        mdiclink_reg(96) => \mdiclink_reg[96]_net_1\, 
        mdiclink_reg(95) => \mdiclink_reg[95]_net_1\, 
        mdiclink_reg(94) => \mdiclink_reg[94]_net_1\, 
        mdiclink_reg(93) => \mdiclink_reg[93]_net_1\, 
        mdiclink_reg(92) => \mdiclink_reg[92]_net_1\, 
        mdiclink_reg(91) => \mdiclink_reg[91]_net_1\, 
        mdiclink_reg(90) => \mdiclink_reg[90]_net_1\, 
        mdiclink_reg(89) => \mdiclink_reg[89]_net_1\, 
        mdiclink_reg(88) => \mdiclink_reg[88]_net_1\, 
        mdiclink_reg(87) => \mdiclink_reg[87]_net_1\, 
        mdiclink_reg(86) => \mdiclink_reg[86]_net_1\, 
        mdiclink_reg(85) => \mdiclink_reg[85]_net_1\, 
        mdiclink_reg(84) => \mdiclink_reg[84]_net_1\, 
        mdiclink_reg(83) => \mdiclink_reg[83]_net_1\, 
        mdiclink_reg(82) => \mdiclink_reg[82]_net_1\, 
        mdiclink_reg(81) => \mdiclink_reg[81]_net_1\, 
        mdiclink_reg(80) => \mdiclink_reg[80]_net_1\, 
        mdiclink_reg(79) => \mdiclink_reg[79]_net_1\, 
        mdiclink_reg(78) => \mdiclink_reg[78]_net_1\, 
        mdiclink_reg(77) => \mdiclink_reg[77]_net_1\, 
        mdiclink_reg(76) => \mdiclink_reg[76]_net_1\, 
        mdiclink_reg(75) => \mdiclink_reg[75]_net_1\, 
        mdiclink_reg(74) => \mdiclink_reg[74]_net_1\, 
        mdiclink_reg(73) => \mdiclink_reg[73]_net_1\, 
        mdiclink_reg(72) => \mdiclink_reg[72]_net_1\, 
        mdiclink_reg(71) => \mdiclink_reg[71]_net_1\, 
        mdiclink_reg(70) => \mdiclink_reg[70]_net_1\, 
        mdiclink_reg(69) => \mdiclink_reg[69]_net_1\, 
        mdiclink_reg(68) => \mdiclink_reg[68]_net_1\, 
        mdiclink_reg(67) => \mdiclink_reg[67]_net_1\, 
        mdiclink_reg(66) => \mdiclink_reg[66]_net_1\, 
        mdiclink_reg(65) => \mdiclink_reg[65]_net_1\, 
        mdiclink_reg(64) => \mdiclink_reg[64]_net_1\, 
        mdiclink_reg(63) => \mdiclink_reg[63]_net_1\, 
        mdiclink_reg(62) => \mdiclink_reg[62]_net_1\, 
        mdiclink_reg(61) => \mdiclink_reg[61]_net_1\, 
        mdiclink_reg(60) => \mdiclink_reg[60]_net_1\, 
        mdiclink_reg(59) => \mdiclink_reg[59]_net_1\, 
        mdiclink_reg(58) => \mdiclink_reg[58]_net_1\, 
        mdiclink_reg(57) => \mdiclink_reg[57]_net_1\, 
        mdiclink_reg(56) => \mdiclink_reg[56]_net_1\, 
        mdiclink_reg(55) => \mdiclink_reg[55]_net_1\, 
        mdiclink_reg(54) => \mdiclink_reg[54]_net_1\, 
        mdiclink_reg(53) => \mdiclink_reg[53]_net_1\, 
        mdiclink_reg(52) => \mdiclink_reg[52]_net_1\, 
        mdiclink_reg(51) => \mdiclink_reg[51]_net_1\, 
        mdiclink_reg(50) => \mdiclink_reg[50]_net_1\, 
        mdiclink_reg(49) => \mdiclink_reg[49]_net_1\, 
        mdiclink_reg(48) => \mdiclink_reg[48]_net_1\, 
        mdiclink_reg(47) => \mdiclink_reg[47]_net_1\, 
        mdiclink_reg(46) => \mdiclink_reg[46]_net_1\, 
        mdiclink_reg(45) => \mdiclink_reg[45]_net_1\, 
        mdiclink_reg(44) => \mdiclink_reg[44]_net_1\, 
        mdiclink_reg(43) => \mdiclink_reg[43]_net_1\, 
        mdiclink_reg(42) => \mdiclink_reg[42]_net_1\, 
        mdiclink_reg(41) => \mdiclink_reg[41]_net_1\, 
        mdiclink_reg(40) => \mdiclink_reg[40]_net_1\, 
        mdiclink_reg(39) => \mdiclink_reg[39]_net_1\, 
        mdiclink_reg(38) => \mdiclink_reg[38]_net_1\, 
        mdiclink_reg(37) => \mdiclink_reg[37]_net_1\, 
        mdiclink_reg(36) => \mdiclink_reg[36]_net_1\, 
        mdiclink_reg(35) => \mdiclink_reg[35]_net_1\, 
        mdiclink_reg(34) => \mdiclink_reg[34]_net_1\, 
        mdiclink_reg(33) => \mdiclink_reg[33]_net_1\, 
        mdiclink_reg(32) => \mdiclink_reg[32]_net_1\, 
        mdiclink_reg(31) => \mdiclink_reg[31]_net_1\, 
        mdiclink_reg(30) => \mdiclink_reg[30]_net_1\, 
        mdiclink_reg(29) => \mdiclink_reg[29]_net_1\, 
        mdiclink_reg(28) => \mdiclink_reg[28]_net_1\, 
        mdiclink_reg(27) => \mdiclink_reg[27]_net_1\, 
        mdiclink_reg(26) => \mdiclink_reg[26]_net_1\, 
        mdiclink_reg(25) => \mdiclink_reg[25]_net_1\, 
        mdiclink_reg(24) => \mdiclink_reg[24]_net_1\, 
        mdiclink_reg(23) => \mdiclink_reg[23]_net_1\, 
        mdiclink_reg(22) => \mdiclink_reg[22]_net_1\, 
        mdiclink_reg(21) => \mdiclink_reg[21]_net_1\, 
        mdiclink_reg(20) => \mdiclink_reg[20]_net_1\, 
        mdiclink_reg(19) => \mdiclink_reg[19]_net_1\, 
        mdiclink_reg(18) => \mdiclink_reg[18]_net_1\, 
        mdiclink_reg(17) => \mdiclink_reg[17]_net_1\, 
        mdiclink_reg(16) => \mdiclink_reg[16]_net_1\, 
        mdiclink_reg(15) => \mdiclink_reg[15]_net_1\, 
        mdiclink_reg(14) => \mdiclink_reg[14]_net_1\, 
        mdiclink_reg(13) => \mdiclink_reg[13]_net_1\, 
        mdiclink_reg(12) => \mdiclink_reg[12]_net_1\, 
        mdiclink_reg(11) => \mdiclink_reg[11]_net_1\, 
        mdiclink_reg(10) => \mdiclink_reg[10]_net_1\, 
        mdiclink_reg(9) => \mdiclink_reg[9]_net_1\, 
        mdiclink_reg(8) => \mdiclink_reg[8]_net_1\, 
        mdiclink_reg(7) => \mdiclink_reg[7]_net_1\, 
        mdiclink_reg(6) => \mdiclink_reg[6]_net_1\, 
        mdiclink_reg(5) => \mdiclink_reg[5]_net_1\, 
        mdiclink_reg(4) => \mdiclink_reg[4]_net_1\, 
        mdiclink_reg(3) => \mdiclink_reg[3]_net_1\, 
        mdiclink_reg(2) => \mdiclink_reg[2]_net_1\, 
        mdiclink_reg(1) => \mdiclink_reg[1]_net_1\, 
        mdiclink_reg(0) => \mdiclink_reg[0]_net_1\, 
        b11_OFWNT9L_8tZ(167) => \b11_OFWNT9L_8tZ[167]\, 
        b11_OFWNT9L_8tZ(166) => \b11_OFWNT9L_8tZ[166]\, 
        b11_OFWNT9L_8tZ(165) => \b11_OFWNT9L_8tZ[165]\, 
        b11_OFWNT9L_8tZ(164) => \b11_OFWNT9L_8tZ[164]\, 
        b11_OFWNT9L_8tZ(163) => \b11_OFWNT9L_8tZ[163]\, 
        b11_OFWNT9L_8tZ(162) => \b11_OFWNT9L_8tZ[162]\, 
        b11_OFWNT9L_8tZ(161) => \b11_OFWNT9L_8tZ[161]\, 
        b11_OFWNT9L_8tZ(160) => \b11_OFWNT9L_8tZ[160]\, 
        b11_OFWNT9L_8tZ(159) => \b11_OFWNT9L_8tZ[159]\, 
        b11_OFWNT9L_8tZ(158) => \b11_OFWNT9L_8tZ[158]\, 
        b11_OFWNT9L_8tZ(157) => \b11_OFWNT9L_8tZ[157]\, 
        b11_OFWNT9L_8tZ(156) => \b11_OFWNT9L_8tZ[156]\, 
        b11_OFWNT9L_8tZ(155) => \b11_OFWNT9L_8tZ[155]\, 
        b11_OFWNT9L_8tZ(154) => \b11_OFWNT9L_8tZ[154]\, 
        b11_OFWNT9L_8tZ(153) => \b11_OFWNT9L_8tZ[153]\, 
        b11_OFWNT9L_8tZ(152) => \b11_OFWNT9L_8tZ[152]\, 
        b11_OFWNT9L_8tZ(151) => \b11_OFWNT9L_8tZ[151]\, 
        b11_OFWNT9L_8tZ(150) => \b11_OFWNT9L_8tZ[150]\, 
        b11_OFWNT9L_8tZ(149) => \b11_OFWNT9L_8tZ[149]\, 
        b11_OFWNT9L_8tZ(148) => \b11_OFWNT9L_8tZ[148]\, 
        b11_OFWNT9L_8tZ(147) => \b11_OFWNT9L_8tZ[147]\, 
        b11_OFWNT9L_8tZ(146) => \b11_OFWNT9L_8tZ[146]\, 
        b11_OFWNT9L_8tZ(145) => \b11_OFWNT9L_8tZ[145]\, 
        b11_OFWNT9L_8tZ(144) => \b11_OFWNT9L_8tZ[144]\, 
        b11_OFWNT9L_8tZ(143) => \b11_OFWNT9L_8tZ[143]\, 
        b11_OFWNT9L_8tZ(142) => \b11_OFWNT9L_8tZ[142]\, 
        b11_OFWNT9L_8tZ(141) => \b11_OFWNT9L_8tZ[141]\, 
        b11_OFWNT9L_8tZ(140) => \b11_OFWNT9L_8tZ[140]\, 
        b11_OFWNT9L_8tZ(139) => \b11_OFWNT9L_8tZ[139]\, 
        b11_OFWNT9L_8tZ(138) => \b11_OFWNT9L_8tZ[138]\, 
        b11_OFWNT9L_8tZ(137) => \b11_OFWNT9L_8tZ[137]\, 
        b11_OFWNT9L_8tZ(136) => \b11_OFWNT9L_8tZ[136]\, 
        b11_OFWNT9L_8tZ(135) => \b11_OFWNT9L_8tZ[135]\, 
        b11_OFWNT9L_8tZ(134) => \b11_OFWNT9L_8tZ[134]\, 
        b11_OFWNT9L_8tZ(133) => \b11_OFWNT9L_8tZ[133]\, 
        b11_OFWNT9L_8tZ(132) => \b11_OFWNT9L_8tZ[132]\, 
        b11_OFWNT9L_8tZ(131) => \b11_OFWNT9L_8tZ[131]\, 
        b11_OFWNT9L_8tZ(130) => \b11_OFWNT9L_8tZ[130]\, 
        b11_OFWNT9L_8tZ(129) => \b11_OFWNT9L_8tZ[129]\, 
        b11_OFWNT9L_8tZ(128) => \b11_OFWNT9L_8tZ[128]\, 
        b11_OFWNT9L_8tZ(127) => \b11_OFWNT9L_8tZ[127]\, 
        b11_OFWNT9L_8tZ(126) => \b11_OFWNT9L_8tZ[126]\, 
        b11_OFWNT9L_8tZ(125) => \b11_OFWNT9L_8tZ[125]\, 
        b11_OFWNT9L_8tZ(124) => \b11_OFWNT9L_8tZ[124]\, 
        b11_OFWNT9L_8tZ(123) => \b11_OFWNT9L_8tZ[123]\, 
        b11_OFWNT9L_8tZ(122) => \b11_OFWNT9L_8tZ[122]\, 
        b11_OFWNT9L_8tZ(121) => \b11_OFWNT9L_8tZ[121]\, 
        b11_OFWNT9L_8tZ(120) => \b11_OFWNT9L_8tZ[120]\, 
        b11_OFWNT9L_8tZ(119) => \b11_OFWNT9L_8tZ[119]\, 
        b11_OFWNT9L_8tZ(118) => \b11_OFWNT9L_8tZ[118]\, 
        b11_OFWNT9L_8tZ(117) => \b11_OFWNT9L_8tZ[117]\, 
        b11_OFWNT9L_8tZ(116) => \b11_OFWNT9L_8tZ[116]\, 
        b11_OFWNT9L_8tZ(115) => \b11_OFWNT9L_8tZ[115]\, 
        b11_OFWNT9L_8tZ(114) => \b11_OFWNT9L_8tZ[114]\, 
        b11_OFWNT9L_8tZ(113) => \b11_OFWNT9L_8tZ[113]\, 
        b11_OFWNT9L_8tZ(112) => \b11_OFWNT9L_8tZ[112]\, 
        b11_OFWNT9L_8tZ(111) => \b11_OFWNT9L_8tZ[111]\, 
        b11_OFWNT9L_8tZ(110) => \b11_OFWNT9L_8tZ[110]\, 
        b11_OFWNT9L_8tZ(109) => \b11_OFWNT9L_8tZ[109]\, 
        b11_OFWNT9L_8tZ(108) => \b11_OFWNT9L_8tZ[108]\, 
        b11_OFWNT9L_8tZ(107) => \b11_OFWNT9L_8tZ[107]\, 
        b11_OFWNT9L_8tZ(106) => \b11_OFWNT9L_8tZ[106]\, 
        b11_OFWNT9L_8tZ(105) => \b11_OFWNT9L_8tZ[105]\, 
        b11_OFWNT9L_8tZ(104) => \b11_OFWNT9L_8tZ[104]\, 
        b11_OFWNT9L_8tZ(103) => \b11_OFWNT9L_8tZ[103]\, 
        b11_OFWNT9L_8tZ(102) => \b11_OFWNT9L_8tZ[102]\, 
        b11_OFWNT9L_8tZ(101) => \b11_OFWNT9L_8tZ[101]\, 
        b11_OFWNT9L_8tZ(100) => \b11_OFWNT9L_8tZ[100]\, 
        b11_OFWNT9L_8tZ(99) => \b11_OFWNT9L_8tZ[99]\, 
        b11_OFWNT9L_8tZ(98) => \b11_OFWNT9L_8tZ[98]\, 
        b11_OFWNT9L_8tZ(97) => \b11_OFWNT9L_8tZ[97]\, 
        b11_OFWNT9L_8tZ(96) => \b11_OFWNT9L_8tZ[96]\, 
        b11_OFWNT9L_8tZ(95) => \b11_OFWNT9L_8tZ[95]\, 
        b11_OFWNT9L_8tZ(94) => \b11_OFWNT9L_8tZ[94]\, 
        b11_OFWNT9L_8tZ(93) => \b11_OFWNT9L_8tZ[93]\, 
        b11_OFWNT9L_8tZ(92) => \b11_OFWNT9L_8tZ[92]\, 
        b11_OFWNT9L_8tZ(91) => \b11_OFWNT9L_8tZ[91]\, 
        b11_OFWNT9L_8tZ(90) => \b11_OFWNT9L_8tZ[90]\, 
        b11_OFWNT9L_8tZ(89) => \b11_OFWNT9L_8tZ[89]\, 
        b11_OFWNT9L_8tZ(88) => \b11_OFWNT9L_8tZ[88]\, 
        b11_OFWNT9L_8tZ(87) => \b11_OFWNT9L_8tZ[87]\, 
        b11_OFWNT9L_8tZ(86) => \b11_OFWNT9L_8tZ[86]\, 
        b11_OFWNT9L_8tZ(85) => \b11_OFWNT9L_8tZ[85]\, 
        b11_OFWNT9L_8tZ(84) => \b11_OFWNT9L_8tZ[84]\, 
        b11_OFWNT9L_8tZ(83) => \b11_OFWNT9L_8tZ[83]\, 
        b11_OFWNT9L_8tZ(82) => \b11_OFWNT9L_8tZ[82]\, 
        b11_OFWNT9L_8tZ(81) => \b11_OFWNT9L_8tZ[81]\, 
        b11_OFWNT9L_8tZ(80) => \b11_OFWNT9L_8tZ[80]\, 
        b11_OFWNT9L_8tZ(79) => \b11_OFWNT9L_8tZ[79]\, 
        b11_OFWNT9L_8tZ(78) => \b11_OFWNT9L_8tZ[78]\, 
        b11_OFWNT9L_8tZ(77) => \b11_OFWNT9L_8tZ[77]\, 
        b11_OFWNT9L_8tZ(76) => \b11_OFWNT9L_8tZ[76]\, 
        b11_OFWNT9L_8tZ(75) => \b11_OFWNT9L_8tZ[75]\, 
        b11_OFWNT9L_8tZ(74) => \b11_OFWNT9L_8tZ[74]\, 
        b11_OFWNT9L_8tZ(73) => \b11_OFWNT9L_8tZ[73]\, 
        b11_OFWNT9L_8tZ(72) => \b11_OFWNT9L_8tZ[72]\, 
        b11_OFWNT9L_8tZ(71) => \b11_OFWNT9L_8tZ[71]\, 
        b11_OFWNT9L_8tZ(70) => \b11_OFWNT9L_8tZ[70]\, 
        b11_OFWNT9L_8tZ(69) => \b11_OFWNT9L_8tZ[69]\, 
        b11_OFWNT9L_8tZ(68) => \b11_OFWNT9L_8tZ[68]\, 
        b11_OFWNT9L_8tZ(67) => \b11_OFWNT9L_8tZ[67]\, 
        b11_OFWNT9L_8tZ(66) => \b11_OFWNT9L_8tZ[66]\, 
        b11_OFWNT9L_8tZ(65) => \b11_OFWNT9L_8tZ[65]\, 
        b11_OFWNT9L_8tZ(64) => \b11_OFWNT9L_8tZ[64]\, 
        b11_OFWNT9L_8tZ(63) => \b11_OFWNT9L_8tZ[63]\, 
        b11_OFWNT9L_8tZ(62) => \b11_OFWNT9L_8tZ[62]\, 
        b11_OFWNT9L_8tZ(61) => \b11_OFWNT9L_8tZ[61]\, 
        b11_OFWNT9L_8tZ(60) => \b11_OFWNT9L_8tZ[60]\, 
        b11_OFWNT9L_8tZ(59) => \b11_OFWNT9L_8tZ[59]\, 
        b11_OFWNT9L_8tZ(58) => \b11_OFWNT9L_8tZ[58]\, 
        b11_OFWNT9L_8tZ(57) => \b11_OFWNT9L_8tZ[57]\, 
        b11_OFWNT9L_8tZ(56) => \b11_OFWNT9L_8tZ[56]\, 
        b11_OFWNT9L_8tZ(55) => \b11_OFWNT9L_8tZ[55]\, 
        b11_OFWNT9L_8tZ(54) => \b11_OFWNT9L_8tZ[54]\, 
        b11_OFWNT9L_8tZ(53) => \b11_OFWNT9L_8tZ[53]\, 
        b11_OFWNT9L_8tZ(52) => \b11_OFWNT9L_8tZ[52]\, 
        b11_OFWNT9L_8tZ(51) => \b11_OFWNT9L_8tZ[51]\, 
        b11_OFWNT9L_8tZ(50) => \b11_OFWNT9L_8tZ[50]\, 
        b11_OFWNT9L_8tZ(49) => \b11_OFWNT9L_8tZ[49]\, 
        b11_OFWNT9L_8tZ(48) => \b11_OFWNT9L_8tZ[48]\, 
        b11_OFWNT9L_8tZ(47) => \b11_OFWNT9L_8tZ[47]\, 
        b11_OFWNT9L_8tZ(46) => \b11_OFWNT9L_8tZ[46]\, 
        b11_OFWNT9L_8tZ(45) => \b11_OFWNT9L_8tZ[45]\, 
        b11_OFWNT9L_8tZ(44) => \b11_OFWNT9L_8tZ[44]\, 
        b11_OFWNT9L_8tZ(43) => \b11_OFWNT9L_8tZ[43]\, 
        b11_OFWNT9L_8tZ(42) => \b11_OFWNT9L_8tZ[42]\, 
        b11_OFWNT9L_8tZ(41) => \b11_OFWNT9L_8tZ[41]\, 
        b11_OFWNT9L_8tZ(40) => \b11_OFWNT9L_8tZ[40]\, 
        b11_OFWNT9L_8tZ(39) => \b11_OFWNT9L_8tZ[39]\, 
        b11_OFWNT9L_8tZ(38) => \b11_OFWNT9L_8tZ[38]\, 
        b11_OFWNT9L_8tZ(37) => \b11_OFWNT9L_8tZ[37]\, 
        b11_OFWNT9L_8tZ(36) => \b11_OFWNT9L_8tZ[36]\, 
        b11_OFWNT9L_8tZ(35) => \b11_OFWNT9L_8tZ[35]\, 
        b11_OFWNT9L_8tZ(34) => \b11_OFWNT9L_8tZ[34]\, 
        b11_OFWNT9L_8tZ(33) => \b11_OFWNT9L_8tZ[33]\, 
        b11_OFWNT9L_8tZ(32) => \b11_OFWNT9L_8tZ[32]\, 
        b11_OFWNT9L_8tZ(31) => \b11_OFWNT9L_8tZ[31]\, 
        b11_OFWNT9L_8tZ(30) => \b11_OFWNT9L_8tZ[30]\, 
        b11_OFWNT9L_8tZ(29) => \b11_OFWNT9L_8tZ[29]\, 
        b11_OFWNT9L_8tZ(28) => \b11_OFWNT9L_8tZ[28]\, 
        b11_OFWNT9L_8tZ(27) => \b11_OFWNT9L_8tZ[27]\, 
        b11_OFWNT9L_8tZ(26) => \b11_OFWNT9L_8tZ[26]\, 
        b11_OFWNT9L_8tZ(25) => \b11_OFWNT9L_8tZ[25]\, 
        b11_OFWNT9L_8tZ(24) => \b11_OFWNT9L_8tZ[24]\, 
        b11_OFWNT9L_8tZ(23) => \b11_OFWNT9L_8tZ[23]\, 
        b11_OFWNT9L_8tZ(22) => \b11_OFWNT9L_8tZ[22]\, 
        b11_OFWNT9L_8tZ(21) => \b11_OFWNT9L_8tZ[21]\, 
        b11_OFWNT9L_8tZ(20) => \b11_OFWNT9L_8tZ[20]\, 
        b11_OFWNT9L_8tZ(19) => \b11_OFWNT9L_8tZ[19]\, 
        b11_OFWNT9L_8tZ(18) => \b11_OFWNT9L_8tZ[18]\, 
        b11_OFWNT9L_8tZ(17) => \b11_OFWNT9L_8tZ[17]\, 
        b11_OFWNT9L_8tZ(16) => \b11_OFWNT9L_8tZ[16]\, 
        b11_OFWNT9L_8tZ(15) => \b11_OFWNT9L_8tZ[15]\, 
        b11_OFWNT9L_8tZ(14) => \b11_OFWNT9L_8tZ[14]\, 
        b11_OFWNT9L_8tZ(13) => \b11_OFWNT9L_8tZ[13]\, 
        b11_OFWNT9L_8tZ(12) => \b11_OFWNT9L_8tZ[12]\, 
        b11_OFWNT9L_8tZ(11) => \b11_OFWNT9L_8tZ[11]\, 
        b11_OFWNT9L_8tZ(10) => \b11_OFWNT9L_8tZ[10]\, 
        b11_OFWNT9L_8tZ(9) => \b11_OFWNT9L_8tZ[9]\, 
        b11_OFWNT9L_8tZ(8) => \b11_OFWNT9L_8tZ[8]\, 
        b11_OFWNT9L_8tZ(7) => \b11_OFWNT9L_8tZ[7]\, 
        b11_OFWNT9L_8tZ(6) => \b11_OFWNT9L_8tZ[6]\, 
        b11_OFWNT9L_8tZ(5) => \b11_OFWNT9L_8tZ[5]\, 
        b11_OFWNT9L_8tZ(4) => \b11_OFWNT9L_8tZ[4]\, 
        b11_OFWNT9L_8tZ(3) => \b11_OFWNT9L_8tZ[3]\, 
        b11_OFWNT9L_8tZ(2) => \b11_OFWNT9L_8tZ[2]\, 
        b11_OFWNT9L_8tZ(1) => \b11_OFWNT9L_8tZ[1]\, 
        b11_OFWNT9L_8tZ(0) => \b11_OFWNT9L_8tZ[0]\, 
        IICE_comm2iice(11) => IICE_comm2iice(11), 
        IICE_comm2iice(10) => IICE_comm2iice(10), 
        IICE_comm2iice(9) => IICE_comm2iice(9), IICE_comm2iice(8)
         => nc2, IICE_comm2iice(7) => nc1, IICE_comm2iice(6) => 
        IICE_comm2iice(6), IICE_comm2iice(5) => IICE_comm2iice(5), 
        IICE_comm2iice(4) => IICE_comm2iice(4), IICE_comm2iice(3)
         => IICE_comm2iice(3), IICE_comm2iice(2) => 
        IICE_comm2iice(2), IICE_comm2iice(1) => IICE_comm2iice(1), 
        IICE_comm2iice(0) => IICE_comm2iice(0), N_145_i => 
        N_145_i, N_1261_i => N_1261_i, b5_voSc3 => b5_voSc3, 
        b9_OFWNT9_ab => b9_OFWNT9_ab, b13_wRBtT_ME83hHx => 
        \b13_wRBtT_ME83hHx\, b5_voSc3_i => b5_voSc3_i, 
        b10_OFWNT9_Y2x => b10_OFWNT9_Y2x, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0);
    
    \mdiclink_reg[155]\ : SLE
      port map(D => RX_FIFO_Empty, CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[155]_net_1\);
    
    \mdiclink_reg[134]\ : SLE
      port map(D => RX_packet_depth(4), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[134]_net_1\);
    
    \mdiclink_reg[61]\ : SLE
      port map(D => irx_center_sample, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[61]_net_1\);
    
    \mdiclink_reg[129]\ : SLE
      port map(D => rx_FIFO_UNDERRUN_int, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[129]_net_1\);
    
    \mdiclink_reg[2]\ : SLE
      port map(D => un6(2), CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[2]_net_1\);
    
    \mdiclink_reg[85]\ : SLE
      port map(D => p2s_data(1), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[85]_net_1\);
    
    \mdiclink_reg[49]\ : SLE
      port map(D => manches_in_dly(1), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[49]_net_1\);
    
    \mdiclink_reg[127]\ : SLE
      port map(D => rx_FIFO_OVERFLOW_int, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[127]_net_1\);
    
    \mdiclink_reg[63]\ : SLE
      port map(D => iRX_FIFO_Empty(2), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[63]_net_1\);
    
    \mdiclink_reg[126]\ : SLE
      port map(D => RX_FIFO_Full, CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[126]_net_1\);
    
    \mdiclink_reg[120]\ : SLE
      port map(D => RX_FIFO_DOUT(4), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[120]_net_1\);
    
    \mdiclink_reg[80]\ : SLE
      port map(D => p2s_data(6), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[80]_net_1\);
    
    \mdiclink_reg[159]\ : SLE
      port map(D => TX_FIFO_wr_en, CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[159]_net_1\);
    
    \mdiclink_reg[52]\ : SLE
      port map(D => int_reg(7), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[52]_net_1\);
    
    \mdiclink_reg[87]\ : SLE
      port map(D => packet_available_clear_reg(2), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[87]_net_1\);
    
    \mdiclink_reg[68]\ : SLE
      port map(D => iRX_FIFO_Full(1), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[68]_net_1\);
    
    \mdiclink_reg[31]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[31]_net_1\);
    
    \mdiclink_reg[103]\ : SLE
      port map(D => ReadFIFO_Write_Ptr(1), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[103]_net_1\);
    
    \mdiclink_reg[66]\ : SLE
      port map(D => iRX_FIFO_Full(3), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[66]_net_1\);
    
    \mdiclink_reg[45]\ : SLE
      port map(D => control_reg_3, CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[45]_net_1\);
    
    \mdiclink_reg[157]\ : SLE
      port map(D => TX_FIFO_Empty, CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[157]_net_1\);
    
    \mdiclink_reg[54]\ : SLE
      port map(D => int_reg(5), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[54]_net_1\);
    
    \mdiclink_reg[156]\ : SLE
      port map(D => m2s010_som_sb_0_GPIO_28_SW_RESET, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[156]_net_1\);
    
    \mdiclink_reg[150]\ : SLE
      port map(D => GND_net_1, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[150]_net_1\);
    
    \mdiclink_reg[33]\ : SLE
      port map(D => bd_reset, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[33]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \mdiclink_reg[40]\ : SLE
      port map(D => GND_net_1, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[40]_net_1\);
    
    \mdiclink_reg[105]\ : SLE
      port map(D => RESET, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[105]_net_1\);
    
    \mdiclink_reg[47]\ : SLE
      port map(D => external_loopback, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[47]_net_1\);
    
    \mdiclink_reg[148]\ : SLE
      port map(D => GND_net_1, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[148]_net_1\);
    
    \mdiclink_reg[114]\ : SLE
      port map(D => RX_FIFO_DIN_pipe(1), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[114]_net_1\);
    
    \mdiclink_reg[38]\ : SLE
      port map(D => clkdiv(1), CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[38]_net_1\);
    
    \mdiclink_reg[36]\ : SLE
      port map(D => clkdiv(3), CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[36]_net_1\);
    
    \mdiclink_reg[21]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PRDATA(0), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[21]_net_1\);
    
    \mdiclink_reg[109]\ : SLE
      port map(D => RX_FIFO_DIN_pipe(6), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[109]_net_1\);
    
    \mdiclink_reg[59]\ : SLE
      port map(D => GND_net_1, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[59]_net_1\);
    
    \mdiclink_reg[23]\ : SLE
      port map(D => long_reset, CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[23]_net_1\);
    
    \mdiclink_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PADDR(7), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[6]_net_1\);
    
    \mdiclink_reg[124]\ : SLE
      port map(D => RX_FIFO_DOUT(0), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[124]_net_1\);
    
    \mdiclink_reg[11]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PADDR(2), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[11]_net_1\);
    
    \mdiclink_reg[143]\ : SLE
      port map(D => RX_FIFO_DIN(4), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[143]_net_1\);
    
    \mdiclink_reg[131]\ : SLE
      port map(D => RX_packet_depth(7), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[131]_net_1\);
    
    \mdiclink_reg[9]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PADDR(4), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[9]_net_1\);
    
    \mdiclink_reg[28]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[28]_net_1\);
    
    \mdiclink_reg[163]\ : SLE
      port map(D => up_EOP_del(4), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[163]_net_1\);
    
    \mdiclink_reg[107]\ : SLE
      port map(D => RX_FIFO_DIN_pipe(8), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[107]_net_1\);
    
    \mdiclink_reg[106]\ : SLE
      port map(D => rx_CRC_error_int, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[106]_net_1\);
    
    \mdiclink_reg[100]\ : SLE
      port map(D => un15(8), CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[100]_net_1\);
    
    \mdiclink_reg[26]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[26]_net_1\);
    
    \mdiclink_reg[71]\ : SLE
      port map(D => iRX_FIFO_UNDERRUN(2), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[71]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \mdiclink_reg[55]\ : SLE
      port map(D => int_reg(4), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[55]_net_1\);
    
    \mdiclink_reg[13]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PADDR(0), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[13]_net_1\);
    
    \mdiclink_reg[132]\ : SLE
      port map(D => RX_packet_depth(6), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[132]_net_1\);
    
    \mdiclink_reg[62]\ : SLE
      port map(D => iRX_FIFO_Empty(3), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[62]_net_1\);
    
    \mdiclink_reg[145]\ : SLE
      port map(D => RX_FIFO_DIN(2), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[145]_net_1\);
    
    \mdiclink_reg[154]\ : SLE
      port map(D => RX_FIFO_Full, CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[154]_net_1\);
    
    \mdiclink_reg[165]\ : SLE
      port map(D => up_EOP_del(2), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[165]_net_1\);
    
    \mdiclink_reg[18]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PRDATA(3), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[18]_net_1\);
    
    \mdiclink_reg[8]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PADDR(5), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[8]_net_1\);
    
    \mdiclink_reg[50]\ : SLE
      port map(D => manches_in_dly(0), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[50]_net_1\);
    
    \mdiclink_reg[73]\ : SLE
      port map(D => iRX_FIFO_UNDERRUN(0), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[73]_net_1\);
    
    \mdiclink_reg[16]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PRDATA(5), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[16]_net_1\);
    
    \mdiclink_reg[64]\ : SLE
      port map(D => iRX_FIFO_Empty(1), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[64]_net_1\);
    
    \mdiclink_reg[57]\ : SLE
      port map(D => int_reg(2), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[57]_net_1\);
    
    \mdiclink_reg[78]\ : SLE
      port map(D => MANCHESTER_IN_c, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[78]_net_1\);
    
    \mdiclink_reg[32]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWRITE, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[32]_net_1\);
    
    \mdiclink_reg[149]\ : SLE
      port map(D => GND_net_1, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[149]_net_1\);
    
    \mdiclink_reg[76]\ : SLE
      port map(D => CommsFPGA_CCC_0_LOCK, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[76]_net_1\);
    
    \mdiclink_reg[91]\ : SLE
      port map(D => ReadFIFO_Read_Ptr(0), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[91]_net_1\);
    
    \mdiclink_reg[111]\ : SLE
      port map(D => RX_FIFO_DIN_pipe(4), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[111]_net_1\);
    
    \mdiclink_reg[147]\ : SLE
      port map(D => RX_FIFO_DIN(0), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[147]_net_1\);
    
    \mdiclink_reg[34]\ : SLE
      port map(D => m2s010_som_sb_0_POWER_ON_RESET_N, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[34]_net_1\);
    
    \mdiclink_reg[146]\ : SLE
      port map(D => RX_FIFO_DIN(1), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[146]_net_1\);
    
    \mdiclink_reg[140]\ : SLE
      port map(D => RX_FIFO_DIN(7), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[140]_net_1\);
    
    b8_uKr_IFLY : b3_uKr_x
      port map(b13_nvmFL_fx2rbuQ(6) => IICE_comm2iice(0), 
        b13_nvmFL_fx2rbuQ(5) => IICE_comm2iice(1), 
        b13_nvmFL_fx2rbuQ(4) => IICE_comm2iice(2), 
        b13_nvmFL_fx2rbuQ(3) => IICE_comm2iice(3), 
        b13_nvmFL_fx2rbuQ(2) => IICE_comm2iice(4), 
        b13_nvmFL_fx2rbuQ(1) => IICE_comm2iice(5), 
        b11_uRrc_9urXBb => IICE_comm2iice(6), b3_PLy => 
        IICE_comm2iice(7), b3_PLF => IICE_iice2comm, b7_PLy_PlM
         => b4_PLyF, b7_nUTQ_9u => b7_nUTQ_9u, b7_PSyi_9u => 
        b7_PSyi_9u, b9_OFWNT9_ab => b9_OFWNT9_ab, b9_PbTt39_ab
         => b9_PbTt39_ab, b9_PKFoLX_ab => b9_PKFoLX_ab, 
        b9_vbTtJX_ab => b9_vbTtJX_ab, b8_ubTt3_YG => b8_ubTt3_YG, 
        b9_ibScJX_ab => b9_ibScJX_ab, b7_yYh0_9u => b7_yYh0_9u, 
        b8_nUTQ_XlK => b8_nUTQ_XlK, b8_PSyi_XlK => 
        b12_PSyi_XlK_qHv, b10_OFWNT9_Y2x => b10_OFWNT9_Y2x, 
        b10_PbTt39_Y2x => GND_net_1, b10_PKFoLX_Y2x => 
        b10_PKFoLX_Y2x, b10_vbTtJX_Y2x => b10_vbTtJX_Y2x, 
        b9_ubTt3_Mxf => b9_ubTt3_Mxf, b10_ibScJX_Y2x => GND_net_1, 
        b8_yYh0_XlK => N_1261_i);
    
    \mdiclink_reg[167]\ : SLE
      port map(D => up_EOP_del(0), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[167]_net_1\);
    
    \mdiclink_reg[166]\ : SLE
      port map(D => up_EOP_del(1), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[166]_net_1\);
    
    \mdiclink_reg[1]\ : SLE
      port map(D => GND_net_1, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[1]_net_1\);
    
    \mdiclink_reg[160]\ : SLE
      port map(D => tx_packet_complt, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[160]_net_1\);
    
    \mdiclink_reg[93]\ : SLE
      port map(D => un15(1), CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[93]_net_1\);
    
    \mdiclink_reg[69]\ : SLE
      port map(D => iRX_FIFO_Full(0), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[69]_net_1\);
    
    \mdiclink_reg[104]\ : SLE
      port map(D => ReadFIFO_Write_Ptr(0), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[104]_net_1\);
    
    \mdiclink_reg[112]\ : SLE
      port map(D => RX_FIFO_DIN_pipe(3), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[112]_net_1\);
    
    b4_PfFz : b8_PfFzrNYI_x
      port map(b11_OFWNT9L_8tZ(167) => \b11_OFWNT9L_8tZ[167]\, 
        b11_OFWNT9L_8tZ(166) => \b11_OFWNT9L_8tZ[166]\, 
        b11_OFWNT9L_8tZ(165) => \b11_OFWNT9L_8tZ[165]\, 
        b11_OFWNT9L_8tZ(164) => \b11_OFWNT9L_8tZ[164]\, 
        b11_OFWNT9L_8tZ(163) => \b11_OFWNT9L_8tZ[163]\, 
        b11_OFWNT9L_8tZ(162) => \b11_OFWNT9L_8tZ[162]\, 
        b11_OFWNT9L_8tZ(161) => \b11_OFWNT9L_8tZ[161]\, 
        b11_OFWNT9L_8tZ(160) => \b11_OFWNT9L_8tZ[160]\, 
        b11_OFWNT9L_8tZ(159) => \b11_OFWNT9L_8tZ[159]\, 
        b11_OFWNT9L_8tZ(158) => \b11_OFWNT9L_8tZ[158]\, 
        b11_OFWNT9L_8tZ(157) => \b11_OFWNT9L_8tZ[157]\, 
        b11_OFWNT9L_8tZ(156) => \b11_OFWNT9L_8tZ[156]\, 
        b11_OFWNT9L_8tZ(155) => \b11_OFWNT9L_8tZ[155]\, 
        b11_OFWNT9L_8tZ(154) => \b11_OFWNT9L_8tZ[154]\, 
        b11_OFWNT9L_8tZ(153) => \b11_OFWNT9L_8tZ[153]\, 
        b11_OFWNT9L_8tZ(152) => \b11_OFWNT9L_8tZ[152]\, 
        b11_OFWNT9L_8tZ(151) => \b11_OFWNT9L_8tZ[151]\, 
        b11_OFWNT9L_8tZ(150) => \b11_OFWNT9L_8tZ[150]\, 
        b11_OFWNT9L_8tZ(149) => \b11_OFWNT9L_8tZ[149]\, 
        b11_OFWNT9L_8tZ(148) => \b11_OFWNT9L_8tZ[148]\, 
        b11_OFWNT9L_8tZ(147) => \b11_OFWNT9L_8tZ[147]\, 
        b11_OFWNT9L_8tZ(146) => \b11_OFWNT9L_8tZ[146]\, 
        b11_OFWNT9L_8tZ(145) => \b11_OFWNT9L_8tZ[145]\, 
        b11_OFWNT9L_8tZ(144) => \b11_OFWNT9L_8tZ[144]\, 
        b11_OFWNT9L_8tZ(143) => \b11_OFWNT9L_8tZ[143]\, 
        b11_OFWNT9L_8tZ(142) => \b11_OFWNT9L_8tZ[142]\, 
        b11_OFWNT9L_8tZ(141) => \b11_OFWNT9L_8tZ[141]\, 
        b11_OFWNT9L_8tZ(140) => \b11_OFWNT9L_8tZ[140]\, 
        b11_OFWNT9L_8tZ(139) => \b11_OFWNT9L_8tZ[139]\, 
        b11_OFWNT9L_8tZ(138) => \b11_OFWNT9L_8tZ[138]\, 
        b11_OFWNT9L_8tZ(137) => \b11_OFWNT9L_8tZ[137]\, 
        b11_OFWNT9L_8tZ(136) => \b11_OFWNT9L_8tZ[136]\, 
        b11_OFWNT9L_8tZ(135) => \b11_OFWNT9L_8tZ[135]\, 
        b11_OFWNT9L_8tZ(134) => \b11_OFWNT9L_8tZ[134]\, 
        b11_OFWNT9L_8tZ(133) => \b11_OFWNT9L_8tZ[133]\, 
        b11_OFWNT9L_8tZ(132) => \b11_OFWNT9L_8tZ[132]\, 
        b11_OFWNT9L_8tZ(131) => \b11_OFWNT9L_8tZ[131]\, 
        b11_OFWNT9L_8tZ(130) => \b11_OFWNT9L_8tZ[130]\, 
        b11_OFWNT9L_8tZ(129) => \b11_OFWNT9L_8tZ[129]\, 
        b11_OFWNT9L_8tZ(128) => \b11_OFWNT9L_8tZ[128]\, 
        b11_OFWNT9L_8tZ(127) => \b11_OFWNT9L_8tZ[127]\, 
        b11_OFWNT9L_8tZ(126) => \b11_OFWNT9L_8tZ[126]\, 
        b11_OFWNT9L_8tZ(125) => \b11_OFWNT9L_8tZ[125]\, 
        b11_OFWNT9L_8tZ(124) => \b11_OFWNT9L_8tZ[124]\, 
        b11_OFWNT9L_8tZ(123) => \b11_OFWNT9L_8tZ[123]\, 
        b11_OFWNT9L_8tZ(122) => \b11_OFWNT9L_8tZ[122]\, 
        b11_OFWNT9L_8tZ(121) => \b11_OFWNT9L_8tZ[121]\, 
        b11_OFWNT9L_8tZ(120) => \b11_OFWNT9L_8tZ[120]\, 
        b11_OFWNT9L_8tZ(119) => \b11_OFWNT9L_8tZ[119]\, 
        b11_OFWNT9L_8tZ(118) => \b11_OFWNT9L_8tZ[118]\, 
        b11_OFWNT9L_8tZ(117) => \b11_OFWNT9L_8tZ[117]\, 
        b11_OFWNT9L_8tZ(116) => \b11_OFWNT9L_8tZ[116]\, 
        b11_OFWNT9L_8tZ(115) => \b11_OFWNT9L_8tZ[115]\, 
        b11_OFWNT9L_8tZ(114) => \b11_OFWNT9L_8tZ[114]\, 
        b11_OFWNT9L_8tZ(113) => \b11_OFWNT9L_8tZ[113]\, 
        b11_OFWNT9L_8tZ(112) => \b11_OFWNT9L_8tZ[112]\, 
        b11_OFWNT9L_8tZ(111) => \b11_OFWNT9L_8tZ[111]\, 
        b11_OFWNT9L_8tZ(110) => \b11_OFWNT9L_8tZ[110]\, 
        b11_OFWNT9L_8tZ(109) => \b11_OFWNT9L_8tZ[109]\, 
        b11_OFWNT9L_8tZ(108) => \b11_OFWNT9L_8tZ[108]\, 
        b11_OFWNT9L_8tZ(107) => \b11_OFWNT9L_8tZ[107]\, 
        b11_OFWNT9L_8tZ(106) => \b11_OFWNT9L_8tZ[106]\, 
        b11_OFWNT9L_8tZ(105) => \b11_OFWNT9L_8tZ[105]\, 
        b11_OFWNT9L_8tZ(104) => \b11_OFWNT9L_8tZ[104]\, 
        b11_OFWNT9L_8tZ(103) => \b11_OFWNT9L_8tZ[103]\, 
        b11_OFWNT9L_8tZ(102) => \b11_OFWNT9L_8tZ[102]\, 
        b11_OFWNT9L_8tZ(101) => \b11_OFWNT9L_8tZ[101]\, 
        b11_OFWNT9L_8tZ(100) => \b11_OFWNT9L_8tZ[100]\, 
        b11_OFWNT9L_8tZ(99) => \b11_OFWNT9L_8tZ[99]\, 
        b11_OFWNT9L_8tZ(98) => \b11_OFWNT9L_8tZ[98]\, 
        b11_OFWNT9L_8tZ(97) => \b11_OFWNT9L_8tZ[97]\, 
        b11_OFWNT9L_8tZ(96) => \b11_OFWNT9L_8tZ[96]\, 
        b11_OFWNT9L_8tZ(95) => \b11_OFWNT9L_8tZ[95]\, 
        b11_OFWNT9L_8tZ(94) => \b11_OFWNT9L_8tZ[94]\, 
        b11_OFWNT9L_8tZ(93) => \b11_OFWNT9L_8tZ[93]\, 
        b11_OFWNT9L_8tZ(92) => \b11_OFWNT9L_8tZ[92]\, 
        b11_OFWNT9L_8tZ(91) => \b11_OFWNT9L_8tZ[91]\, 
        b11_OFWNT9L_8tZ(90) => \b11_OFWNT9L_8tZ[90]\, 
        b11_OFWNT9L_8tZ(89) => \b11_OFWNT9L_8tZ[89]\, 
        b11_OFWNT9L_8tZ(88) => \b11_OFWNT9L_8tZ[88]\, 
        b11_OFWNT9L_8tZ(87) => \b11_OFWNT9L_8tZ[87]\, 
        b11_OFWNT9L_8tZ(86) => \b11_OFWNT9L_8tZ[86]\, 
        b11_OFWNT9L_8tZ(85) => \b11_OFWNT9L_8tZ[85]\, 
        b11_OFWNT9L_8tZ(84) => \b11_OFWNT9L_8tZ[84]\, 
        b11_OFWNT9L_8tZ(83) => \b11_OFWNT9L_8tZ[83]\, 
        b11_OFWNT9L_8tZ(82) => \b11_OFWNT9L_8tZ[82]\, 
        b11_OFWNT9L_8tZ(81) => \b11_OFWNT9L_8tZ[81]\, 
        b11_OFWNT9L_8tZ(80) => \b11_OFWNT9L_8tZ[80]\, 
        b11_OFWNT9L_8tZ(79) => \b11_OFWNT9L_8tZ[79]\, 
        b11_OFWNT9L_8tZ(78) => \b11_OFWNT9L_8tZ[78]\, 
        b11_OFWNT9L_8tZ(77) => \b11_OFWNT9L_8tZ[77]\, 
        b11_OFWNT9L_8tZ(76) => \b11_OFWNT9L_8tZ[76]\, 
        b11_OFWNT9L_8tZ(75) => \b11_OFWNT9L_8tZ[75]\, 
        b11_OFWNT9L_8tZ(74) => \b11_OFWNT9L_8tZ[74]\, 
        b11_OFWNT9L_8tZ(73) => \b11_OFWNT9L_8tZ[73]\, 
        b11_OFWNT9L_8tZ(72) => \b11_OFWNT9L_8tZ[72]\, 
        b11_OFWNT9L_8tZ(71) => \b11_OFWNT9L_8tZ[71]\, 
        b11_OFWNT9L_8tZ(70) => \b11_OFWNT9L_8tZ[70]\, 
        b11_OFWNT9L_8tZ(69) => \b11_OFWNT9L_8tZ[69]\, 
        b11_OFWNT9L_8tZ(68) => \b11_OFWNT9L_8tZ[68]\, 
        b11_OFWNT9L_8tZ(67) => \b11_OFWNT9L_8tZ[67]\, 
        b11_OFWNT9L_8tZ(66) => \b11_OFWNT9L_8tZ[66]\, 
        b11_OFWNT9L_8tZ(65) => \b11_OFWNT9L_8tZ[65]\, 
        b11_OFWNT9L_8tZ(64) => \b11_OFWNT9L_8tZ[64]\, 
        b11_OFWNT9L_8tZ(63) => \b11_OFWNT9L_8tZ[63]\, 
        b11_OFWNT9L_8tZ(62) => \b11_OFWNT9L_8tZ[62]\, 
        b11_OFWNT9L_8tZ(61) => \b11_OFWNT9L_8tZ[61]\, 
        b11_OFWNT9L_8tZ(60) => \b11_OFWNT9L_8tZ[60]\, 
        b11_OFWNT9L_8tZ(59) => \b11_OFWNT9L_8tZ[59]\, 
        b11_OFWNT9L_8tZ(58) => \b11_OFWNT9L_8tZ[58]\, 
        b11_OFWNT9L_8tZ(57) => \b11_OFWNT9L_8tZ[57]\, 
        b11_OFWNT9L_8tZ(56) => \b11_OFWNT9L_8tZ[56]\, 
        b11_OFWNT9L_8tZ(55) => \b11_OFWNT9L_8tZ[55]\, 
        b11_OFWNT9L_8tZ(54) => \b11_OFWNT9L_8tZ[54]\, 
        b11_OFWNT9L_8tZ(53) => \b11_OFWNT9L_8tZ[53]\, 
        b11_OFWNT9L_8tZ(52) => \b11_OFWNT9L_8tZ[52]\, 
        b11_OFWNT9L_8tZ(51) => \b11_OFWNT9L_8tZ[51]\, 
        b11_OFWNT9L_8tZ(50) => \b11_OFWNT9L_8tZ[50]\, 
        b11_OFWNT9L_8tZ(49) => \b11_OFWNT9L_8tZ[49]\, 
        b11_OFWNT9L_8tZ(48) => \b11_OFWNT9L_8tZ[48]\, 
        b11_OFWNT9L_8tZ(47) => \b11_OFWNT9L_8tZ[47]\, 
        b11_OFWNT9L_8tZ(46) => \b11_OFWNT9L_8tZ[46]\, 
        b11_OFWNT9L_8tZ(45) => \b11_OFWNT9L_8tZ[45]\, 
        b11_OFWNT9L_8tZ(44) => \b11_OFWNT9L_8tZ[44]\, 
        b11_OFWNT9L_8tZ(43) => \b11_OFWNT9L_8tZ[43]\, 
        b11_OFWNT9L_8tZ(42) => \b11_OFWNT9L_8tZ[42]\, 
        b11_OFWNT9L_8tZ(41) => \b11_OFWNT9L_8tZ[41]\, 
        b11_OFWNT9L_8tZ(40) => \b11_OFWNT9L_8tZ[40]\, 
        b11_OFWNT9L_8tZ(39) => \b11_OFWNT9L_8tZ[39]\, 
        b11_OFWNT9L_8tZ(38) => \b11_OFWNT9L_8tZ[38]\, 
        b11_OFWNT9L_8tZ(37) => \b11_OFWNT9L_8tZ[37]\, 
        b11_OFWNT9L_8tZ(36) => \b11_OFWNT9L_8tZ[36]\, 
        b11_OFWNT9L_8tZ(35) => \b11_OFWNT9L_8tZ[35]\, 
        b11_OFWNT9L_8tZ(34) => \b11_OFWNT9L_8tZ[34]\, 
        b11_OFWNT9L_8tZ(33) => \b11_OFWNT9L_8tZ[33]\, 
        b11_OFWNT9L_8tZ(32) => \b11_OFWNT9L_8tZ[32]\, 
        b11_OFWNT9L_8tZ(31) => \b11_OFWNT9L_8tZ[31]\, 
        b11_OFWNT9L_8tZ(30) => \b11_OFWNT9L_8tZ[30]\, 
        b11_OFWNT9L_8tZ(29) => \b11_OFWNT9L_8tZ[29]\, 
        b11_OFWNT9L_8tZ(28) => \b11_OFWNT9L_8tZ[28]\, 
        b11_OFWNT9L_8tZ(27) => \b11_OFWNT9L_8tZ[27]\, 
        b11_OFWNT9L_8tZ(26) => \b11_OFWNT9L_8tZ[26]\, 
        b11_OFWNT9L_8tZ(25) => \b11_OFWNT9L_8tZ[25]\, 
        b11_OFWNT9L_8tZ(24) => \b11_OFWNT9L_8tZ[24]\, 
        b11_OFWNT9L_8tZ(23) => \b11_OFWNT9L_8tZ[23]\, 
        b11_OFWNT9L_8tZ(22) => \b11_OFWNT9L_8tZ[22]\, 
        b11_OFWNT9L_8tZ(21) => \b11_OFWNT9L_8tZ[21]\, 
        b11_OFWNT9L_8tZ(20) => \b11_OFWNT9L_8tZ[20]\, 
        b11_OFWNT9L_8tZ(19) => \b11_OFWNT9L_8tZ[19]\, 
        b11_OFWNT9L_8tZ(18) => \b11_OFWNT9L_8tZ[18]\, 
        b11_OFWNT9L_8tZ(17) => \b11_OFWNT9L_8tZ[17]\, 
        b11_OFWNT9L_8tZ(16) => \b11_OFWNT9L_8tZ[16]\, 
        b11_OFWNT9L_8tZ(15) => \b11_OFWNT9L_8tZ[15]\, 
        b11_OFWNT9L_8tZ(14) => \b11_OFWNT9L_8tZ[14]\, 
        b11_OFWNT9L_8tZ(13) => \b11_OFWNT9L_8tZ[13]\, 
        b11_OFWNT9L_8tZ(12) => \b11_OFWNT9L_8tZ[12]\, 
        b11_OFWNT9L_8tZ(11) => \b11_OFWNT9L_8tZ[11]\, 
        b11_OFWNT9L_8tZ(10) => \b11_OFWNT9L_8tZ[10]\, 
        b11_OFWNT9L_8tZ(9) => \b11_OFWNT9L_8tZ[9]\, 
        b11_OFWNT9L_8tZ(8) => \b11_OFWNT9L_8tZ[8]\, 
        b11_OFWNT9L_8tZ(7) => \b11_OFWNT9L_8tZ[7]\, 
        b11_OFWNT9L_8tZ(6) => \b11_OFWNT9L_8tZ[6]\, 
        b11_OFWNT9L_8tZ(5) => \b11_OFWNT9L_8tZ[5]\, 
        b11_OFWNT9L_8tZ(4) => \b11_OFWNT9L_8tZ[4]\, 
        b11_OFWNT9L_8tZ(3) => \b11_OFWNT9L_8tZ[3]\, 
        b11_OFWNT9L_8tZ(2) => \b11_OFWNT9L_8tZ[2]\, 
        b11_OFWNT9L_8tZ(1) => \b11_OFWNT9L_8tZ[1]\, 
        b11_OFWNT9L_8tZ(0) => \b11_OFWNT9L_8tZ[0]\, 
        mdiclink_reg(167) => \mdiclink_reg[167]_net_1\, 
        mdiclink_reg(166) => \mdiclink_reg[166]_net_1\, 
        mdiclink_reg(165) => \mdiclink_reg[165]_net_1\, 
        mdiclink_reg(164) => \mdiclink_reg[164]_net_1\, 
        mdiclink_reg(163) => \mdiclink_reg[163]_net_1\, 
        mdiclink_reg(162) => \mdiclink_reg[162]_net_1\, 
        mdiclink_reg(161) => \mdiclink_reg[161]_net_1\, 
        mdiclink_reg(160) => \mdiclink_reg[160]_net_1\, 
        mdiclink_reg(159) => \mdiclink_reg[159]_net_1\, 
        mdiclink_reg(158) => \mdiclink_reg[158]_net_1\, 
        mdiclink_reg(157) => \mdiclink_reg[157]_net_1\, 
        mdiclink_reg(156) => \mdiclink_reg[156]_net_1\, 
        mdiclink_reg(155) => \mdiclink_reg[155]_net_1\, 
        mdiclink_reg(154) => \mdiclink_reg[154]_net_1\, 
        mdiclink_reg(153) => \mdiclink_reg[153]_net_1\, 
        mdiclink_reg(152) => \mdiclink_reg[152]_net_1\, 
        mdiclink_reg(151) => \mdiclink_reg[151]_net_1\, 
        mdiclink_reg(150) => \mdiclink_reg[150]_net_1\, 
        mdiclink_reg(149) => \mdiclink_reg[149]_net_1\, 
        mdiclink_reg(148) => \mdiclink_reg[148]_net_1\, 
        mdiclink_reg(147) => \mdiclink_reg[147]_net_1\, 
        mdiclink_reg(146) => \mdiclink_reg[146]_net_1\, 
        mdiclink_reg(145) => \mdiclink_reg[145]_net_1\, 
        mdiclink_reg(144) => \mdiclink_reg[144]_net_1\, 
        mdiclink_reg(143) => \mdiclink_reg[143]_net_1\, 
        mdiclink_reg(142) => \mdiclink_reg[142]_net_1\, 
        mdiclink_reg(141) => \mdiclink_reg[141]_net_1\, 
        mdiclink_reg(140) => \mdiclink_reg[140]_net_1\, 
        mdiclink_reg(139) => \mdiclink_reg[139]_net_1\, 
        mdiclink_reg(138) => \mdiclink_reg[138]_net_1\, 
        mdiclink_reg(137) => \mdiclink_reg[137]_net_1\, 
        mdiclink_reg(136) => \mdiclink_reg[136]_net_1\, 
        mdiclink_reg(135) => \mdiclink_reg[135]_net_1\, 
        mdiclink_reg(134) => \mdiclink_reg[134]_net_1\, 
        mdiclink_reg(133) => \mdiclink_reg[133]_net_1\, 
        mdiclink_reg(132) => \mdiclink_reg[132]_net_1\, 
        mdiclink_reg(131) => \mdiclink_reg[131]_net_1\, 
        mdiclink_reg(130) => \mdiclink_reg[130]_net_1\, 
        mdiclink_reg(129) => \mdiclink_reg[129]_net_1\, 
        mdiclink_reg(128) => \mdiclink_reg[128]_net_1\, 
        mdiclink_reg(127) => \mdiclink_reg[127]_net_1\, 
        mdiclink_reg(126) => \mdiclink_reg[126]_net_1\, 
        mdiclink_reg(125) => \mdiclink_reg[125]_net_1\, 
        mdiclink_reg(124) => \mdiclink_reg[124]_net_1\, 
        mdiclink_reg(123) => \mdiclink_reg[123]_net_1\, 
        mdiclink_reg(122) => \mdiclink_reg[122]_net_1\, 
        mdiclink_reg(121) => \mdiclink_reg[121]_net_1\, 
        mdiclink_reg(120) => \mdiclink_reg[120]_net_1\, 
        mdiclink_reg(119) => \mdiclink_reg[119]_net_1\, 
        mdiclink_reg(118) => \mdiclink_reg[118]_net_1\, 
        mdiclink_reg(117) => \mdiclink_reg[117]_net_1\, 
        mdiclink_reg(116) => \mdiclink_reg[116]_net_1\, 
        mdiclink_reg(115) => \mdiclink_reg[115]_net_1\, 
        mdiclink_reg(114) => \mdiclink_reg[114]_net_1\, 
        mdiclink_reg(113) => \mdiclink_reg[113]_net_1\, 
        mdiclink_reg(112) => \mdiclink_reg[112]_net_1\, 
        mdiclink_reg(111) => \mdiclink_reg[111]_net_1\, 
        mdiclink_reg(110) => \mdiclink_reg[110]_net_1\, 
        mdiclink_reg(109) => \mdiclink_reg[109]_net_1\, 
        mdiclink_reg(108) => \mdiclink_reg[108]_net_1\, 
        mdiclink_reg(107) => \mdiclink_reg[107]_net_1\, 
        mdiclink_reg(106) => \mdiclink_reg[106]_net_1\, 
        mdiclink_reg(105) => \mdiclink_reg[105]_net_1\, 
        mdiclink_reg(104) => \mdiclink_reg[104]_net_1\, 
        mdiclink_reg(103) => \mdiclink_reg[103]_net_1\, 
        mdiclink_reg(102) => \mdiclink_reg[102]_net_1\, 
        mdiclink_reg(101) => \mdiclink_reg[101]_net_1\, 
        mdiclink_reg(100) => \mdiclink_reg[100]_net_1\, 
        mdiclink_reg(99) => \mdiclink_reg[99]_net_1\, 
        mdiclink_reg(98) => \mdiclink_reg[98]_net_1\, 
        mdiclink_reg(97) => \mdiclink_reg[97]_net_1\, 
        mdiclink_reg(96) => \mdiclink_reg[96]_net_1\, 
        mdiclink_reg(95) => \mdiclink_reg[95]_net_1\, 
        mdiclink_reg(94) => \mdiclink_reg[94]_net_1\, 
        mdiclink_reg(93) => \mdiclink_reg[93]_net_1\, 
        mdiclink_reg(92) => \mdiclink_reg[92]_net_1\, 
        mdiclink_reg(91) => \mdiclink_reg[91]_net_1\, 
        mdiclink_reg(90) => \mdiclink_reg[90]_net_1\, 
        mdiclink_reg(89) => \mdiclink_reg[89]_net_1\, 
        mdiclink_reg(88) => \mdiclink_reg[88]_net_1\, 
        mdiclink_reg(87) => \mdiclink_reg[87]_net_1\, 
        mdiclink_reg(86) => \mdiclink_reg[86]_net_1\, 
        mdiclink_reg(85) => \mdiclink_reg[85]_net_1\, 
        mdiclink_reg(84) => \mdiclink_reg[84]_net_1\, 
        mdiclink_reg(83) => \mdiclink_reg[83]_net_1\, 
        mdiclink_reg(82) => \mdiclink_reg[82]_net_1\, 
        mdiclink_reg(81) => \mdiclink_reg[81]_net_1\, 
        mdiclink_reg(80) => \mdiclink_reg[80]_net_1\, 
        mdiclink_reg(79) => \mdiclink_reg[79]_net_1\, 
        mdiclink_reg(78) => \mdiclink_reg[78]_net_1\, 
        mdiclink_reg(77) => \mdiclink_reg[77]_net_1\, 
        mdiclink_reg(76) => \mdiclink_reg[76]_net_1\, 
        mdiclink_reg(75) => \mdiclink_reg[75]_net_1\, 
        mdiclink_reg(74) => \mdiclink_reg[74]_net_1\, 
        mdiclink_reg(73) => \mdiclink_reg[73]_net_1\, 
        mdiclink_reg(72) => \mdiclink_reg[72]_net_1\, 
        mdiclink_reg(71) => \mdiclink_reg[71]_net_1\, 
        mdiclink_reg(70) => \mdiclink_reg[70]_net_1\, 
        mdiclink_reg(69) => \mdiclink_reg[69]_net_1\, 
        mdiclink_reg(68) => \mdiclink_reg[68]_net_1\, 
        mdiclink_reg(67) => \mdiclink_reg[67]_net_1\, 
        mdiclink_reg(66) => \mdiclink_reg[66]_net_1\, 
        mdiclink_reg(65) => \mdiclink_reg[65]_net_1\, 
        mdiclink_reg(64) => \mdiclink_reg[64]_net_1\, 
        mdiclink_reg(63) => \mdiclink_reg[63]_net_1\, 
        mdiclink_reg(62) => \mdiclink_reg[62]_net_1\, 
        mdiclink_reg(61) => \mdiclink_reg[61]_net_1\, 
        mdiclink_reg(60) => \mdiclink_reg[60]_net_1\, 
        mdiclink_reg(59) => \mdiclink_reg[59]_net_1\, 
        mdiclink_reg(58) => \mdiclink_reg[58]_net_1\, 
        mdiclink_reg(57) => \mdiclink_reg[57]_net_1\, 
        mdiclink_reg(56) => \mdiclink_reg[56]_net_1\, 
        mdiclink_reg(55) => \mdiclink_reg[55]_net_1\, 
        mdiclink_reg(54) => \mdiclink_reg[54]_net_1\, 
        mdiclink_reg(53) => \mdiclink_reg[53]_net_1\, 
        mdiclink_reg(52) => \mdiclink_reg[52]_net_1\, 
        mdiclink_reg(51) => \mdiclink_reg[51]_net_1\, 
        mdiclink_reg(50) => \mdiclink_reg[50]_net_1\, 
        mdiclink_reg(49) => \mdiclink_reg[49]_net_1\, 
        mdiclink_reg(48) => \mdiclink_reg[48]_net_1\, 
        mdiclink_reg(47) => \mdiclink_reg[47]_net_1\, 
        mdiclink_reg(46) => \mdiclink_reg[46]_net_1\, 
        mdiclink_reg(45) => \mdiclink_reg[45]_net_1\, 
        mdiclink_reg(44) => \mdiclink_reg[44]_net_1\, 
        mdiclink_reg(43) => \mdiclink_reg[43]_net_1\, 
        mdiclink_reg(42) => \mdiclink_reg[42]_net_1\, 
        mdiclink_reg(41) => \mdiclink_reg[41]_net_1\, 
        mdiclink_reg(40) => \mdiclink_reg[40]_net_1\, 
        mdiclink_reg(39) => \mdiclink_reg[39]_net_1\, 
        mdiclink_reg(38) => \mdiclink_reg[38]_net_1\, 
        mdiclink_reg(37) => \mdiclink_reg[37]_net_1\, 
        mdiclink_reg(36) => \mdiclink_reg[36]_net_1\, 
        mdiclink_reg(35) => \mdiclink_reg[35]_net_1\, 
        mdiclink_reg(34) => \mdiclink_reg[34]_net_1\, 
        mdiclink_reg(33) => \mdiclink_reg[33]_net_1\, 
        mdiclink_reg(32) => \mdiclink_reg[32]_net_1\, 
        mdiclink_reg(31) => \mdiclink_reg[31]_net_1\, 
        mdiclink_reg(30) => \mdiclink_reg[30]_net_1\, 
        mdiclink_reg(29) => \mdiclink_reg[29]_net_1\, 
        mdiclink_reg(28) => \mdiclink_reg[28]_net_1\, 
        mdiclink_reg(27) => \mdiclink_reg[27]_net_1\, 
        mdiclink_reg(26) => \mdiclink_reg[26]_net_1\, 
        mdiclink_reg(25) => \mdiclink_reg[25]_net_1\, 
        mdiclink_reg(24) => \mdiclink_reg[24]_net_1\, 
        mdiclink_reg(23) => \mdiclink_reg[23]_net_1\, 
        mdiclink_reg(22) => \mdiclink_reg[22]_net_1\, 
        mdiclink_reg(21) => \mdiclink_reg[21]_net_1\, 
        mdiclink_reg(20) => \mdiclink_reg[20]_net_1\, 
        mdiclink_reg(19) => \mdiclink_reg[19]_net_1\, 
        mdiclink_reg(18) => \mdiclink_reg[18]_net_1\, 
        mdiclink_reg(17) => \mdiclink_reg[17]_net_1\, 
        mdiclink_reg(16) => \mdiclink_reg[16]_net_1\, 
        mdiclink_reg(15) => \mdiclink_reg[15]_net_1\, 
        mdiclink_reg(14) => \mdiclink_reg[14]_net_1\, 
        mdiclink_reg(13) => \mdiclink_reg[13]_net_1\, 
        mdiclink_reg(12) => \mdiclink_reg[12]_net_1\, 
        mdiclink_reg(11) => \mdiclink_reg[11]_net_1\, 
        mdiclink_reg(10) => \mdiclink_reg[10]_net_1\, 
        mdiclink_reg(9) => \mdiclink_reg[9]_net_1\, 
        mdiclink_reg(8) => \mdiclink_reg[8]_net_1\, 
        mdiclink_reg(7) => \mdiclink_reg[7]_net_1\, 
        mdiclink_reg(6) => \mdiclink_reg[6]_net_1\, 
        mdiclink_reg(5) => \mdiclink_reg[5]_net_1\, 
        mdiclink_reg(4) => \mdiclink_reg[4]_net_1\, 
        mdiclink_reg(3) => \mdiclink_reg[3]_net_1\, 
        mdiclink_reg(2) => \mdiclink_reg[2]_net_1\, 
        mdiclink_reg(1) => \mdiclink_reg[1]_net_1\, 
        mdiclink_reg(0) => \mdiclink_reg[0]_net_1\, 
        IICE_comm2iice_4 => IICE_comm2iice(11), IICE_comm2iice_0
         => IICE_comm2iice(7), IICE_comm2iice_3 => 
        IICE_comm2iice(10), b10_nYBzIXrKbK_0 => 
        \b10_nYBzIXrKbK[1]\, b7_PSyi_9u => b7_PSyi_9u, 
        b12_PSyi_XlK_qHv => b12_PSyi_XlK_qHv, CommsFPGA_CCC_0_GL0
         => CommsFPGA_CCC_0_GL0);
    
    \mdiclink_reg[22]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PREADY, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[22]_net_1\);
    
    \mdiclink_reg[98]\ : SLE
      port map(D => GND_net_1, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[98]_net_1\);
    
    \mdiclink_reg[81]\ : SLE
      port map(D => p2s_data(5), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[81]_net_1\);
    
    \mdiclink_reg[121]\ : SLE
      port map(D => RX_FIFO_DOUT(3), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[121]_net_1\);
    
    \mdiclink_reg[96]\ : SLE
      port map(D => un15(4), CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[96]_net_1\);
    
    \mdiclink_reg[138]\ : SLE
      port map(D => RX_packet_depth(0), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[138]_net_1\);
    
    \mdiclink_reg[65]\ : SLE
      port map(D => iRX_FIFO_Empty(0), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[65]_net_1\);
    
    \mdiclink_reg[24]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[24]_net_1\);
    
    \mdiclink_reg[39]\ : SLE
      port map(D => clkdiv(0), CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[39]_net_1\);
    
    \mdiclink_reg[83]\ : SLE
      port map(D => p2s_data(3), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[83]_net_1\);
    
    \mdiclink_reg[12]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PADDR(1), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[12]_net_1\);
    
    \mdiclink_reg[122]\ : SLE
      port map(D => RX_FIFO_DOUT(2), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[122]_net_1\);
    
    \mdiclink_reg[60]\ : SLE
      port map(D => int_reg_clr, CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[60]_net_1\);
    
    \mdiclink_reg[41]\ : SLE
      port map(D => TX_FIFO_RST, CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[41]_net_1\);
    
    \mdiclink_reg[151]\ : SLE
      port map(D => RX_packet_depth_status, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[151]_net_1\);
    
    \mdiclink_reg[67]\ : SLE
      port map(D => iRX_FIFO_Full(2), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[67]_net_1\);
    
    \mdiclink_reg[88]\ : SLE
      port map(D => packet_available_clear_reg(1), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[88]_net_1\);
    
    \mdiclink_reg[4]\ : SLE
      port map(D => un6(4), CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[4]_net_1\);
    
    \mdiclink_reg[72]\ : SLE
      port map(D => iRX_FIFO_UNDERRUN(1), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[72]_net_1\);
    
    \mdiclink_reg[86]\ : SLE
      port map(D => p2s_data(0), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[86]_net_1\);
    
    \mdiclink_reg[14]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PRDATA(7), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[14]_net_1\);
    
    \mdiclink_reg[35]\ : SLE
      port map(D => block_int_until_rd, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[35]_net_1\);
    
    \mdiclink_reg[133]\ : SLE
      port map(D => RX_packet_depth(5), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[133]_net_1\);
    
    \mdiclink_reg[43]\ : SLE
      port map(D => start_tx_FIFO, CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[43]_net_1\);
    
    \mdiclink_reg[152]\ : SLE
      port map(D => TX_FIFO_Full, CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[152]_net_1\);
    
    \mdiclink_reg[144]\ : SLE
      port map(D => RX_FIFO_DIN(3), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[144]_net_1\);
    
    \mdiclink_reg[74]\ : SLE
      port map(D => rx_packet_avail_int, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[74]_net_1\);
    
    \mdiclink_reg[164]\ : SLE
      port map(D => up_EOP_del(3), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[164]_net_1\);
    
    b5_nUTGT : b7_OCByLXC_Z1_x_0
      port map(IICE_comm2iice(11) => IICE_comm2iice(11), 
        IICE_comm2iice(10) => IICE_comm2iice(10), 
        IICE_comm2iice(9) => IICE_comm2iice(9), IICE_comm2iice(8)
         => IICE_comm2iice(8), IICE_comm2iice(7) => 
        IICE_comm2iice(7), b9_PKFoLX_ab => b9_PKFoLX_ab, 
        b8_nUTQ_XlK => b8_nUTQ_XlK, b7_nUTQ_9u => b7_nUTQ_9u, 
        b10_PKFoLX_Y2x => b10_PKFoLX_Y2x, b10_vbTtJX_Y2x => 
        b10_vbTtJX_Y2x, b9_vbTtJX_ab => b9_vbTtJX_ab, b8_ubTt3_YG
         => b8_ubTt3_YG, N_145_i => N_145_i, b13_wRBtT_ME83hHx
         => \b13_wRBtT_ME83hHx\, b9_ubTt3_Mxf => b9_ubTt3_Mxf, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, b5_voSc3_i
         => b5_voSc3_i, b5_voSc3 => b5_voSc3);
    
    \mdiclink_reg[29]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[29]_net_1\);
    
    \mdiclink_reg[30]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[30]_net_1\);
    
    \mdiclink_reg[48]\ : SLE
      port map(D => control_reg_0, CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[48]_net_1\);
    
    \mdiclink_reg[37]\ : SLE
      port map(D => clkdiv(2), CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[37]_net_1\);
    
    \mdiclink_reg[46]\ : SLE
      port map(D => control_reg_2, CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[46]_net_1\);
    
    \mdiclink_reg[135]\ : SLE
      port map(D => RX_packet_depth(3), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[135]_net_1\);
    
    \mdiclink_reg[118]\ : SLE
      port map(D => RX_FIFO_DOUT(6), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[118]_net_1\);
    
    \mdiclink_reg[5]\ : SLE
      port map(D => un6(5), CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[5]_net_1\);
    
    \mdiclink_reg[19]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PRDATA(2), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[19]_net_1\);
    
    \mdiclink_reg[92]\ : SLE
      port map(D => un15(0), CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[92]_net_1\);
    
    \mdiclink_reg[25]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[25]_net_1\);
    
    \mdiclink_reg[3]\ : SLE
      port map(D => un6(3), CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[3]_net_1\);
    
    \mdiclink_reg[101]\ : SLE
      port map(D => un15(9), CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[101]_net_1\);
    
    \mdiclink_reg[139]\ : SLE
      port map(D => RX_packet_depth_status, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[139]_net_1\);
    
    \mdiclink_reg[79]\ : SLE
      port map(D => p2s_data(7), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[79]_net_1\);
    
    \mdiclink_reg[20]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PRDATA(1), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[20]_net_1\);
    
    \mdiclink_reg[94]\ : SLE
      port map(D => un15(2), CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[94]_net_1\);
    
    \mdiclink_reg[27]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[27]_net_1\);
    
    \mdiclink_reg[128]\ : SLE
      port map(D => RX_FIFO_rd_en, CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[128]_net_1\);
    
    \mdiclink_reg[51]\ : SLE
      port map(D => iNRZ_data, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[51]_net_1\);
    
    \mdiclink_reg[15]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PRDATA(6), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[15]_net_1\);
    
    \mdiclink_reg[102]\ : SLE
      port map(D => un15(10), CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[102]_net_1\);
    
    b13_wRBtT_ME83hHx : SLE
      port map(D => \b10_nYBzIXrKbK[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \b13_wRBtT_ME83hHx\);
    
    \mdiclink_reg[113]\ : SLE
      port map(D => RX_FIFO_DIN_pipe(2), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[113]_net_1\);
    
    \mdiclink_reg[137]\ : SLE
      port map(D => RX_packet_depth(1), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[137]_net_1\);
    
    \mdiclink_reg[136]\ : SLE
      port map(D => RX_packet_depth(2), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[136]_net_1\);
    
    \mdiclink_reg[82]\ : SLE
      port map(D => p2s_data(4), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[82]_net_1\);
    
    \mdiclink_reg[130]\ : SLE
      port map(D => rx_packet_complt, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[130]_net_1\);
    
    \mdiclink_reg[10]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PADDR(3), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[10]_net_1\);
    
    \mdiclink_reg[75]\ : SLE
      port map(D => TX_FIFO_Empty, CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[75]_net_1\);
    
    \mdiclink_reg[0]\ : SLE
      port map(D => un6(0), CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[0]_net_1\);
    
    \mdiclink_reg[53]\ : SLE
      port map(D => int_reg(6), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[53]_net_1\);
    
    \mdiclink_reg[17]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PRDATA(4), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[17]_net_1\);
    
    \mdiclink_reg[158]\ : SLE
      port map(D => TX_FIFO_Full, CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[158]_net_1\);
    
    \mdiclink_reg[115]\ : SLE
      port map(D => RX_FIFO_DIN_pipe(0), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[115]_net_1\);
    
    \mdiclink_reg[84]\ : SLE
      port map(D => p2s_data(2), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[84]_net_1\);
    
    \mdiclink_reg[58]\ : SLE
      port map(D => int_reg(1), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[58]_net_1\);
    
    \mdiclink_reg[70]\ : SLE
      port map(D => iRX_FIFO_UNDERRUN(3), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[70]_net_1\);
    
    \mdiclink_reg[123]\ : SLE
      port map(D => RX_FIFO_DOUT(1), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[123]_net_1\);
    
    \mdiclink_reg[77]\ : SLE
      port map(D => MANCH_OUT_P_c, CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[77]_net_1\);
    
    \mdiclink_reg[56]\ : SLE
      port map(D => int_reg(3), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[56]_net_1\);
    
    \mdiclink_reg[99]\ : SLE
      port map(D => un15(7), CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[99]_net_1\);
    
    \mdiclink_reg[42]\ : SLE
      port map(D => rx_FIFO_rst_reg, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[42]_net_1\);
    
    \mdiclink_reg[141]\ : SLE
      port map(D => RX_FIFO_DIN(6), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[141]_net_1\);
    
    \mdiclink_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PADDR(6), CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mdiclink_reg[7]_net_1\);
    
    \mdiclink_reg[161]\ : SLE
      port map(D => iup_EOP, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[161]_net_1\);
    
    \mdiclink_reg[119]\ : SLE
      port map(D => RX_FIFO_DOUT(5), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[119]_net_1\);
    
    \mdiclink_reg[44]\ : SLE
      port map(D => internal_loopback, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[44]_net_1\);
    
    \mdiclink_reg[125]\ : SLE
      port map(D => RX_FIFO_Empty, CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[125]_net_1\);
    
    \mdiclink_reg[95]\ : SLE
      port map(D => un15(3), CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[95]_net_1\);
    
    \mdiclink_reg[153]\ : SLE
      port map(D => TX_FIFO_Empty, CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[153]_net_1\);
    
    \mdiclink_reg[142]\ : SLE
      port map(D => RX_FIFO_DIN(5), CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mdiclink_reg[142]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b9_ORbIwXaEF_32s_2497421375_0s_x_0 is

    port( b6_uS_MrX           : in    std_logic_vector(1 downto 0);
          b3_ORb_0            : out   std_logic;
          N_39                : in    std_logic;
          b9_PLF_6lNa2_0_a2_0 : in    std_logic;
          b7_nFG0rDY          : in    std_logic;
          b12_ORbIwXaEF_bd    : in    std_logic;
          b5_OvyH3            : in    std_logic;
          b6_nv_0CC           : in    std_logic;
          tck                 : in    std_logic
        );

end b9_ORbIwXaEF_32s_2497421375_0s_x_0;

architecture DEF_ARCH of b9_ORbIwXaEF_32s_2497421375_0s_x_0 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal N_65, N_65_i, \b3_ORb[32]_net_1\, VCC_net_1, 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, GND_net_1, 
        \b3_ORb[31]_net_1\, \b3_ORb[30]_net_1\, 
        \b3_ORb[29]_net_1\, \b3_ORb[28]_net_1\, 
        \b3_ORb[27]_net_1\, \b3_ORb[26]_net_1\, 
        \b3_ORb[25]_net_1\, \b3_ORb[24]_net_1\, 
        \b3_ORb[23]_net_1\, \b3_ORb[22]_net_1\, 
        \b3_ORb[21]_net_1\, \b3_ORb[20]_net_1\, 
        \b3_ORb[19]_net_1\, \b3_ORb[18]_net_1\, 
        \b3_ORb[17]_net_1\, \b3_ORb[16]_net_1\, 
        \b3_ORb[15]_net_1\, \b3_ORb[14]_net_1\, 
        \b3_ORb[13]_net_1\, \b3_ORb[12]_net_1\, 
        \b3_ORb[11]_net_1\, \b3_ORb[10]_net_1\, \b3_ORb[9]_net_1\, 
        \b3_ORb[8]_net_1\, \b3_ORb[7]_net_1\, \b3_ORb[6]_net_1\, 
        \b3_ORb[5]_net_1\, \b3_ORb[4]_net_1\, \b3_ORb[3]_net_1\, 
        \b3_ORb[2]_net_1\, un1_b3_ORb9_1_or, 
        \un1_b3_ORb9_1_or_0_a2_0\ : std_logic;

begin 


    \b3_ORb[7]\ : SLE
      port map(D => \b3_ORb[8]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[7]_net_1\);
    
    b3_ORb_0_sqmuxa_0_a2 : CFG2
      generic map(INIT => x"8")

      port map(A => N_39, B => b12_ORbIwXaEF_bd, Y => N_65);
    
    \b3_ORb[9]\ : SLE
      port map(D => \b3_ORb[10]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[9]_net_1\);
    
    \b3_ORb[3]\ : SLE
      port map(D => \b3_ORb[4]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => VCC_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[3]_net_1\);
    
    \b3_ORb[23]\ : SLE
      port map(D => \b3_ORb[24]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => VCC_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[23]_net_1\);
    
    \b3_ORb[22]\ : SLE
      port map(D => \b3_ORb[23]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[22]_net_1\);
    
    \b3_ORb[1]\ : SLE
      port map(D => \b3_ORb[2]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => VCC_net_1, LAT => 
        GND_net_1, Q => b3_ORb_0);
    
    \b3_ORb[10]\ : SLE
      port map(D => \b3_ORb[11]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[10]_net_1\);
    
    un1_b3_ORb9_1_or_0_a2_0 : CFG3
      generic map(INIT => x"C8")

      port map(A => b5_OvyH3, B => b12_ORbIwXaEF_bd, C => 
        b7_nFG0rDY, Y => \un1_b3_ORb9_1_or_0_a2_0\);
    
    \b3_ORb[16]\ : SLE
      port map(D => \b3_ORb[17]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => VCC_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[16]_net_1\);
    
    \b3_ORb[11]\ : SLE
      port map(D => \b3_ORb[12]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[11]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \b3_ORb[17]\ : SLE
      port map(D => \b3_ORb[18]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => VCC_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[17]_net_1\);
    
    \b3_ORb[5]\ : SLE
      port map(D => \b3_ORb[6]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => VCC_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[5]_net_1\);
    
    \b3_ORb[28]\ : SLE
      port map(D => \b3_ORb[29]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[28]_net_1\);
    
    \b3_ORb[6]\ : SLE
      port map(D => \b3_ORb[7]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => VCC_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[6]_net_1\);
    
    \b3_ORb[29]\ : SLE
      port map(D => \b3_ORb[30]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => VCC_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[29]_net_1\);
    
    \b3_ORb[13]\ : SLE
      port map(D => \b3_ORb[14]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[13]_net_1\);
    
    \b3_ORb[12]\ : SLE
      port map(D => \b3_ORb[13]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[12]_net_1\);
    
    \b3_ORb[24]\ : SLE
      port map(D => \b3_ORb[25]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => VCC_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[24]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \b3_ORb[2]\ : SLE
      port map(D => \b3_ORb[3]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => VCC_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[2]_net_1\);
    
    \b3_ORb[25]\ : SLE
      port map(D => \b3_ORb[26]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[25]_net_1\);
    
    \b3_ORb[30]\ : SLE
      port map(D => \b3_ORb[31]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[30]_net_1\);
    
    b3_ORb_0_sqmuxa_0_a2_RNIQN0L2 : CFG2
      generic map(INIT => x"E")

      port map(A => N_65, B => un1_b3_ORb9_1_or, Y => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\);
    
    \b3_ORb[18]\ : SLE
      port map(D => \b3_ORb[19]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => VCC_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[18]_net_1\);
    
    \b3_ORb[20]\ : SLE
      port map(D => \b3_ORb[21]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => VCC_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[20]_net_1\);
    
    \b3_ORb[19]\ : SLE
      port map(D => \b3_ORb[20]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[19]_net_1\);
    
    \b3_ORb[31]\ : SLE
      port map(D => \b3_ORb[32]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[31]_net_1\);
    
    \b3_ORb[14]\ : SLE
      port map(D => \b3_ORb[15]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => VCC_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[14]_net_1\);
    
    \b3_ORb[26]\ : SLE
      port map(D => \b3_ORb[27]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[26]_net_1\);
    
    \b3_ORb[4]\ : SLE
      port map(D => \b3_ORb[5]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => VCC_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[4]_net_1\);
    
    \b3_ORb[21]\ : SLE
      port map(D => \b3_ORb[22]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => VCC_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[21]_net_1\);
    
    \b3_ORb[8]\ : SLE
      port map(D => \b3_ORb[9]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[8]_net_1\);
    
    \b3_ORb[15]\ : SLE
      port map(D => \b3_ORb[16]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[15]_net_1\);
    
    un1_b3_ORb9_1_or_0_a2 : CFG4
      generic map(INIT => x"4000")

      port map(A => b6_uS_MrX(1), B => b6_uS_MrX(0), C => 
        \un1_b3_ORb9_1_or_0_a2_0\, D => b9_PLF_6lNa2_0_a2_0, Y
         => un1_b3_ORb9_1_or);
    
    \b3_ORb[27]\ : SLE
      port map(D => \b3_ORb[28]_net_1\, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => VCC_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[27]_net_1\);
    
    b3_ORb_0_sqmuxa_0_a2_RNI9O7A : CFG1
      generic map(INIT => "01")

      port map(A => N_65, Y => N_65_i);
    
    \b3_ORb[32]\ : SLE
      port map(D => b6_nv_0CC, CLK => tck, EN => 
        \b3_ORb_0_sqmuxa_0_a2_RNIQN0L2\, ALn => VCC_net_1, ADn
         => VCC_net_1, SLn => N_65_i, SD => VCC_net_1, LAT => 
        GND_net_1, Q => \b3_ORb[32]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity jtag_interface_x_0 is

    port( b6_uS_MrX           : out   std_logic_vector(1 downto 0);
          atck                : in    std_logic;
          atms                : in    std_logic;
          atdi                : in    std_logic;
          atdo                : out   std_logic;
          atrstb              : in    std_logic;
          b6_nv_0CC           : out   std_logic;
          ch_update           : out   std_logic;
          N_52                : out   std_logic;
          b5_OvyH3            : out   std_logic;
          N_39                : out   std_logic;
          b7_nFG0rDY          : out   std_logic;
          N_27                : in    std_logic;
          N_73                : out   std_logic;
          b9_PLF_6lNa2_0_a2_0 : out   std_logic;
          dr2_tck_i           : out   std_logic;
          hcr_update          : out   std_logic
        );

end jtag_interface_x_0;

architecture DEF_ARCH of jtag_interface_x_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component UJTAG
    port( UDRCAP : out   std_logic;
          UDRSH  : out   std_logic;
          UDRUPD : out   std_logic;
          UIREG  : out   std_logic_vector(7 downto 0);
          URSTB  : out   std_logic;
          UDRCK  : out   std_logic;
          UTDI   : out   std_logic;
          UTDO   : in    std_logic := 'U';
          TDI    : in    std_logic := 'U';
          TMS    : in    std_logic := 'U';
          TCK    : in    std_logic := 'U';
          TRSTB  : in    std_logic := 'U';
          TDO    : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal b10_8Kz_rKlrtX, identify_clk_int, \b6_uS_MrX[4]\, 
        \b6_uS_MrX[3]\, \b6_uS_MrX[2]\, b3_1Um, 
        b9_PLF_6lNa2_0_a2_0_net_1, \N_73\, 
        identify_clk2_no_clk_buffer_needed, \b6_uS_MrX[1]\, 
        \b6_uS_MrX[0]\, b9_PLF_6lNa2, \b7_nFG0rDY\, \b5_OvyH3\, 
        \UIREGdummy[0]\, \UIREGdummy[7]\, URSTBdummy, GND_net_1, 
        VCC_net_1 : std_logic;

begin 

    b6_uS_MrX(1) <= \b6_uS_MrX[1]\;
    b6_uS_MrX(0) <= \b6_uS_MrX[0]\;
    b5_OvyH3 <= \b5_OvyH3\;
    b7_nFG0rDY <= \b7_nFG0rDY\;
    N_73 <= \N_73\;
    b9_PLF_6lNa2_0_a2_0 <= b9_PLF_6lNa2_0_a2_0_net_1;

    b10_nv_ywKMm9X_0_a2 : CFG4
      generic map(INIT => x"2000")

      port map(A => \b7_nFG0rDY\, B => \b6_uS_MrX[1]\, C => 
        \b6_uS_MrX[0]\, D => b9_PLF_6lNa2_0_a2_0_net_1, Y => N_39);
    
    b10_8Kz_fFfsjX_0_a2 : CFG3
      generic map(INIT => x"20")

      port map(A => \b6_uS_MrX[1]\, B => \b6_uS_MrX[0]\, C => 
        b9_PLF_6lNa2_0_a2_0_net_1, Y => \N_73\);
    
    b9_nv_oQwfYF_3_0_a2 : CFG4
      generic map(INIT => x"2000")

      port map(A => identify_clk2_no_clk_buffer_needed, B => 
        \b6_uS_MrX[1]\, C => \b6_uS_MrX[0]\, D => 
        b9_PLF_6lNa2_0_a2_0_net_1, Y => ch_update);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \b9_PLF_6lNa2_0_a2_0\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \b6_uS_MrX[4]\, B => \b6_uS_MrX[3]\, C => 
        \b6_uS_MrX[2]\, D => b3_1Um, Y => 
        b9_PLF_6lNa2_0_a2_0_net_1);
    
    b9_Rcmi_KsDw : UJTAG
      port map(UDRCAP => \b7_nFG0rDY\, UDRSH => \b5_OvyH3\, 
        UDRUPD => identify_clk2_no_clk_buffer_needed, UIREG(7)
         => \UIREGdummy[7]\, UIREG(6) => b3_1Um, UIREG(5) => 
        \b6_uS_MrX[4]\, UIREG(4) => \b6_uS_MrX[3]\, UIREG(3) => 
        \b6_uS_MrX[2]\, UIREG(2) => \b6_uS_MrX[1]\, UIREG(1) => 
        \b6_uS_MrX[0]\, UIREG(0) => \UIREGdummy[0]\, URSTB => 
        URSTBdummy, UDRCK => identify_clk_int, UTDI => b6_nv_0CC, 
        UTDO => b9_PLF_6lNa2, TDI => atdi, TMS => atms, TCK => 
        atck, TRSTB => atrstb, TDO => atdo);
    
    b8_nv_ZmCtY_0_a2 : CFG4
      generic map(INIT => x"4000")

      port map(A => \b6_uS_MrX[1]\, B => \b5_OvyH3\, C => 
        b9_PLF_6lNa2_0_a2_0_net_1, D => \b6_uS_MrX[0]\, Y => N_52);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b9_PLF_6lNa2_0_a2 : CFG4
      generic map(INIT => x"6000")

      port map(A => \b6_uS_MrX[1]\, B => \b6_uS_MrX[0]\, C => 
        b9_PLF_6lNa2_0_a2_0_net_1, D => N_27, Y => b9_PLF_6lNa2);
    
    b10_8Kz_rKlrtX_RNI2P6B : CLKINT
      port map(A => b10_8Kz_rKlrtX, Y => hcr_update);
    
    jtag_clkint_prim : CLKINT
      port map(A => identify_clk_int, Y => dr2_tck_i);
    
    b10_8Kz_rKlrtX_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => \N_73\, B => 
        identify_clk2_no_clk_buffer_needed, Y => b10_8Kz_rKlrtX);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity b16_Rcmi_qlx9_yHpm7y_6s_1s_0s_0s_8s_0s_0s_1s_6s_7s_x_0 is

    port( b13_nvmFL_fx2rbuQ : out   std_logic_vector(5 downto 0);
          b11_uRrc_WYOFjZ_0 : out   std_logic;
          b5_OvyH3          : in    std_logic;
          b7_nFG0rDY        : in    std_logic;
          tdo_sig           : in    std_logic;
          N_27              : out   std_logic;
          IICE_iice2comm    : in    std_logic;
          b6_nv_0CC         : in    std_logic;
          dr2_tck           : in    std_logic;
          b12_ORbIwXaEF_bd  : out   std_logic;
          N_73              : in    std_logic;
          hcr_update        : in    std_logic
        );

end b16_Rcmi_qlx9_yHpm7y_6s_1s_0s_0s_8s_0s_0s_1s_6s_7s_x_0;

architecture DEF_ARCH of 
        b16_Rcmi_qlx9_yHpm7y_6s_1s_0s_0s_8s_0s_0s_1s_6s_7s_x_0 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \b9_OvyH3_saL[5]_net_1\, GND_net_1, 
        \b9_OvyH3_saL[6]_net_1\, \b12_ORbIwXaEF_bd\, 
        b10_dZst39_EF3_18, \b9_OvyH3_saL[0]_net_1\, 
        \b9_OvyH3_saL[1]_net_1\, b9_OvyH3_saL_0_sqmuxa, 
        \b9_OvyH3_saL[2]_net_1\, \b9_OvyH3_saL[3]_net_1\, 
        \b9_OvyH3_saL[4]_net_1\, \b9_OvyH3_saL[7]_net_1\, 
        \b3_PLF_u_i_m2_1\ : std_logic;

begin 

    b12_ORbIwXaEF_bd <= \b12_ORbIwXaEF_bd\;

    \genblk1.b10_dZst39_EF3[5]\ : SLE
      port map(D => \b9_OvyH3_saL[5]_net_1\, CLK => hcr_update, 
        EN => N_73, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b13_nvmFL_fx2rbuQ(4));
    
    \genblk1.b10_dZst39_EF3[4]\ : SLE
      port map(D => \b9_OvyH3_saL[4]_net_1\, CLK => hcr_update, 
        EN => N_73, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b13_nvmFL_fx2rbuQ(3));
    
    b9_OvyH3_saL_0_sqmuxa_0_a2 : CFG3
      generic map(INIT => x"40")

      port map(A => b7_nFG0rDY, B => b5_OvyH3, C => N_73, Y => 
        b9_OvyH3_saL_0_sqmuxa);
    
    \genblk1.b10_dZst39_EF3[3]\ : SLE
      port map(D => \b9_OvyH3_saL[3]_net_1\, CLK => hcr_update, 
        EN => N_73, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b13_nvmFL_fx2rbuQ(2));
    
    \genblk1.b10_dZst39_EF3[1]\ : SLE
      port map(D => \b9_OvyH3_saL[1]_net_1\, CLK => hcr_update, 
        EN => N_73, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b13_nvmFL_fx2rbuQ(0));
    
    \b9_OvyH3_saL[6]\ : SLE
      port map(D => \b9_OvyH3_saL[7]_net_1\, CLK => dr2_tck, EN
         => b9_OvyH3_saL_0_sqmuxa, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b9_OvyH3_saL[6]_net_1\);
    
    \b9_OvyH3_saL[3]\ : SLE
      port map(D => \b9_OvyH3_saL[4]_net_1\, CLK => dr2_tck, EN
         => b9_OvyH3_saL_0_sqmuxa, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b9_OvyH3_saL[3]_net_1\);
    
    \genblk1.b10_dZst39_EF3[0]\ : SLE
      port map(D => \b9_OvyH3_saL[0]_net_1\, CLK => hcr_update, 
        EN => N_73, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b11_uRrc_WYOFjZ_0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b3_PLF_u_i_m2 : CFG4
      generic map(INIT => x"1F0E")

      port map(A => \b12_ORbIwXaEF_bd\, B => N_73, C => 
        \b3_PLF_u_i_m2_1\, D => IICE_iice2comm, Y => N_27);
    
    \genblk1.b10_dZst39_EF3_18\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \b12_ORbIwXaEF_bd\, B => N_73, C => 
        \b9_OvyH3_saL[7]_net_1\, Y => b10_dZst39_EF3_18);
    
    \genblk1.b10_dZst39_EF3[7]\ : SLE
      port map(D => b10_dZst39_EF3_18, CLK => hcr_update, EN => 
        VCC_net_1, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \b12_ORbIwXaEF_bd\);
    
    \b9_OvyH3_saL[5]\ : SLE
      port map(D => \b9_OvyH3_saL[6]_net_1\, CLK => dr2_tck, EN
         => b9_OvyH3_saL_0_sqmuxa, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b9_OvyH3_saL[5]_net_1\);
    
    \genblk1.b10_dZst39_EF3[6]\ : SLE
      port map(D => \b9_OvyH3_saL[6]_net_1\, CLK => hcr_update, 
        EN => N_73, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b13_nvmFL_fx2rbuQ(5));
    
    \genblk1.b10_dZst39_EF3[2]\ : SLE
      port map(D => \b9_OvyH3_saL[2]_net_1\, CLK => hcr_update, 
        EN => N_73, ALn => VCC_net_1, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        b13_nvmFL_fx2rbuQ(1));
    
    b3_PLF_u_i_m2_1 : CFG3
      generic map(INIT => x"1D")

      port map(A => tdo_sig, B => N_73, C => 
        \b9_OvyH3_saL[0]_net_1\, Y => \b3_PLF_u_i_m2_1\);
    
    \b9_OvyH3_saL[7]\ : SLE
      port map(D => b6_nv_0CC, CLK => dr2_tck, EN => 
        b9_OvyH3_saL_0_sqmuxa, ALn => VCC_net_1, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \b9_OvyH3_saL[7]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \b9_OvyH3_saL[1]\ : SLE
      port map(D => \b9_OvyH3_saL[2]_net_1\, CLK => dr2_tck, EN
         => b9_OvyH3_saL_0_sqmuxa, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b9_OvyH3_saL[1]_net_1\);
    
    \b9_OvyH3_saL[0]\ : SLE
      port map(D => \b9_OvyH3_saL[1]_net_1\, CLK => dr2_tck, EN
         => b9_OvyH3_saL_0_sqmuxa, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b9_OvyH3_saL[0]_net_1\);
    
    \b9_OvyH3_saL[4]\ : SLE
      port map(D => \b9_OvyH3_saL[5]_net_1\, CLK => dr2_tck, EN
         => b9_OvyH3_saL_0_sqmuxa, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b9_OvyH3_saL[4]_net_1\);
    
    \b9_OvyH3_saL[2]\ : SLE
      port map(D => \b9_OvyH3_saL[3]_net_1\, CLK => dr2_tck, EN
         => b9_OvyH3_saL_0_sqmuxa, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \b9_OvyH3_saL[2]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity comm_block_x is

    port( IICE_comm2iice : out   std_logic_vector(0 to 11);
          IICE_iice2comm : in    std_logic;
          atck           : in    std_logic;
          atdi           : in    std_logic;
          atdo           : out   std_logic;
          atms           : in    std_logic;
          atrstb         : in    std_logic
        );

end comm_block_x;

architecture DEF_ARCH of comm_block_x is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component b9_ORbIwXaEF_32s_2497421375_0s_x_0
    port( b6_uS_MrX           : in    std_logic_vector(1 downto 0) := (others => 'U');
          b3_ORb_0            : out   std_logic;
          N_39                : in    std_logic := 'U';
          b9_PLF_6lNa2_0_a2_0 : in    std_logic := 'U';
          b7_nFG0rDY          : in    std_logic := 'U';
          b12_ORbIwXaEF_bd    : in    std_logic := 'U';
          b5_OvyH3            : in    std_logic := 'U';
          b6_nv_0CC           : in    std_logic := 'U';
          tck                 : in    std_logic := 'U'
        );
  end component;

  component jtag_interface_x_0
    port( b6_uS_MrX           : out   std_logic_vector(1 downto 0);
          atck                : in    std_logic := 'U';
          atms                : in    std_logic := 'U';
          atdi                : in    std_logic := 'U';
          atdo                : out   std_logic;
          atrstb              : in    std_logic := 'U';
          b6_nv_0CC           : out   std_logic;
          ch_update           : out   std_logic;
          N_52                : out   std_logic;
          b5_OvyH3            : out   std_logic;
          N_39                : out   std_logic;
          b7_nFG0rDY          : out   std_logic;
          N_27                : in    std_logic := 'U';
          N_73                : out   std_logic;
          b9_PLF_6lNa2_0_a2_0 : out   std_logic;
          dr2_tck_i           : out   std_logic;
          hcr_update          : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component 
        b16_Rcmi_qlx9_yHpm7y_6s_1s_0s_0s_8s_0s_0s_1s_6s_7s_x_0
    port( b13_nvmFL_fx2rbuQ : out   std_logic_vector(5 downto 0);
          b11_uRrc_WYOFjZ_0 : out   std_logic;
          b5_OvyH3          : in    std_logic := 'U';
          b7_nFG0rDY        : in    std_logic := 'U';
          tdo_sig           : in    std_logic := 'U';
          N_27              : out   std_logic;
          IICE_iice2comm    : in    std_logic := 'U';
          b6_nv_0CC         : in    std_logic := 'U';
          dr2_tck           : in    std_logic := 'U';
          b12_ORbIwXaEF_bd  : out   std_logic;
          N_73              : in    std_logic := 'U';
          hcr_update        : in    std_logic := 'U'
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \IICE_comm2iice[11]\, \IICE_comm2iice[7]\, hcr_update, 
        \b11_uRrc_WYOFjZ[0]\, VCC_net_1, GND_net_1, tdo_sig, 
        \jtagi.b6_uS_MrX[0]\, \jtagi.b6_uS_MrX[1]\, 
        \jtagi.b7_nFG0rDY\, \jtagi.b5_OvyH3\, \IICE_comm2iice[9]\, 
        b12_ORbIwXaEF_bd, N_73, N_27, b9_PLF_6lNa2_0_a2_0
         : std_logic;

    for all : b9_ORbIwXaEF_32s_2497421375_0s_x_0
	Use entity work.b9_ORbIwXaEF_32s_2497421375_0s_x_0(DEF_ARCH);
    for all : jtag_interface_x_0
	Use entity work.jtag_interface_x_0(DEF_ARCH);
    for all : b16_Rcmi_qlx9_yHpm7y_6s_1s_0s_0s_8s_0s_0s_1s_6s_7s_x_0
	Use entity work.
        b16_Rcmi_qlx9_yHpm7y_6s_1s_0s_0s_8s_0s_0s_1s_6s_7s_x_0(DEF_ARCH);
begin 

    IICE_comm2iice(7) <= \IICE_comm2iice[7]\;
    IICE_comm2iice(9) <= \IICE_comm2iice[9]\;
    IICE_comm2iice(11) <= \IICE_comm2iice[11]\;

    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    b9_ORb_xNywD : b9_ORbIwXaEF_32s_2497421375_0s_x_0
      port map(b6_uS_MrX(1) => \jtagi.b6_uS_MrX[1]\, b6_uS_MrX(0)
         => \jtagi.b6_uS_MrX[0]\, b3_ORb_0 => tdo_sig, N_39 => 
        \IICE_comm2iice[9]\, b9_PLF_6lNa2_0_a2_0 => 
        b9_PLF_6lNa2_0_a2_0, b7_nFG0rDY => \jtagi.b7_nFG0rDY\, 
        b12_ORbIwXaEF_bd => b12_ORbIwXaEF_bd, b5_OvyH3 => 
        \jtagi.b5_OvyH3\, b6_nv_0CC => \IICE_comm2iice[7]\, tck
         => \IICE_comm2iice[11]\);
    
    jtagi : jtag_interface_x_0
      port map(b6_uS_MrX(1) => \jtagi.b6_uS_MrX[1]\, b6_uS_MrX(0)
         => \jtagi.b6_uS_MrX[0]\, atck => atck, atms => atms, 
        atdi => atdi, atdo => atdo, atrstb => atrstb, b6_nv_0CC
         => \IICE_comm2iice[7]\, ch_update => IICE_comm2iice(8), 
        N_52 => IICE_comm2iice(10), b5_OvyH3 => \jtagi.b5_OvyH3\, 
        N_39 => \IICE_comm2iice[9]\, b7_nFG0rDY => 
        \jtagi.b7_nFG0rDY\, N_27 => N_27, N_73 => N_73, 
        b9_PLF_6lNa2_0_a2_0 => b9_PLF_6lNa2_0_a2_0, dr2_tck_i => 
        \IICE_comm2iice[11]\, hcr_update => hcr_update);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    b7_Rcmi_ql : 
        b16_Rcmi_qlx9_yHpm7y_6s_1s_0s_0s_8s_0s_0s_1s_6s_7s_x_0
      port map(b13_nvmFL_fx2rbuQ(5) => IICE_comm2iice(0), 
        b13_nvmFL_fx2rbuQ(4) => IICE_comm2iice(1), 
        b13_nvmFL_fx2rbuQ(3) => IICE_comm2iice(2), 
        b13_nvmFL_fx2rbuQ(2) => IICE_comm2iice(3), 
        b13_nvmFL_fx2rbuQ(1) => IICE_comm2iice(4), 
        b13_nvmFL_fx2rbuQ(0) => IICE_comm2iice(5), 
        b11_uRrc_WYOFjZ_0 => \b11_uRrc_WYOFjZ[0]\, b5_OvyH3 => 
        \jtagi.b5_OvyH3\, b7_nFG0rDY => \jtagi.b7_nFG0rDY\, 
        tdo_sig => tdo_sig, N_27 => N_27, IICE_iice2comm => 
        IICE_iice2comm, b6_nv_0CC => \IICE_comm2iice[7]\, dr2_tck
         => \IICE_comm2iice[11]\, b12_ORbIwXaEF_bd => 
        b12_ORbIwXaEF_bd, N_73 => N_73, hcr_update => hcr_update);
    
    \b11_uRrc_9urXBb[0]\ : CFG4
      generic map(INIT => x"4000")

      port map(A => \jtagi.b6_uS_MrX[1]\, B => 
        \b11_uRrc_WYOFjZ[0]\, C => b9_PLF_6lNa2_0_a2_0, D => 
        \jtagi.b6_uS_MrX[0]\, Y => IICE_comm2iice(6));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity syn_identify_core0_0 is

    port( un6                              : in    std_logic_vector(5 downto 0);
          CoreAPB3_0_APBmslave0_PRDATA     : in    std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PADDR      : in    std_logic_vector(7 downto 0);
          clkdiv                           : in    std_logic_vector(3 downto 0);
          CoreAPB3_0_APBmslave0_PWDATA     : in    std_logic_vector(7 downto 0);
          manches_in_dly                   : in    std_logic_vector(1 downto 0);
          iRX_FIFO_Full                    : in    std_logic_vector(3 downto 0);
          iRX_FIFO_Empty                   : in    std_logic_vector(3 downto 0);
          int_reg                          : in    std_logic_vector(7 downto 1);
          iRX_FIFO_UNDERRUN                : in    std_logic_vector(3 downto 0);
          ReadFIFO_Read_Ptr                : in    std_logic_vector(1 downto 0);
          packet_available_clear_reg       : in    std_logic_vector(2 downto 0);
          p2s_data                         : in    std_logic_vector(7 downto 0);
          RX_FIFO_DIN_pipe                 : in    std_logic_vector(8 downto 0);
          ReadFIFO_Write_Ptr               : in    std_logic_vector(1 downto 0);
          un15                             : in    std_logic_vector(10 downto 0);
          RX_FIFO_DOUT                     : in    std_logic_vector(8 downto 0);
          RX_packet_depth                  : in    std_logic_vector(7 downto 0);
          RX_FIFO_DIN                      : in    std_logic_vector(7 downto 0);
          up_EOP_del                       : in    std_logic_vector(5 downto 0);
          control_reg_0                    : in    std_logic;
          control_reg_2                    : in    std_logic;
          control_reg_3                    : in    std_logic;
          CommsFPGA_CCC_0_GL0              : in    std_logic;
          long_reset                       : in    std_logic;
          CoreAPB3_0_APBmslave0_PREADY     : in    std_logic;
          block_int_until_rd               : in    std_logic;
          m2s010_som_sb_0_POWER_ON_RESET_N : in    std_logic;
          bd_reset                         : in    std_logic;
          CoreAPB3_0_APBmslave0_PWRITE     : in    std_logic;
          iNRZ_data                        : in    std_logic;
          external_loopback                : in    std_logic;
          internal_loopback                : in    std_logic;
          start_tx_FIFO                    : in    std_logic;
          rx_FIFO_rst_reg                  : in    std_logic;
          TX_FIFO_RST                      : in    std_logic;
          irx_center_sample                : in    std_logic;
          int_reg_clr                      : in    std_logic;
          MANCHESTER_IN_c                  : in    std_logic;
          MANCH_OUT_P_c                    : in    std_logic;
          CommsFPGA_CCC_0_LOCK             : in    std_logic;
          TX_FIFO_Empty                    : in    std_logic;
          rx_packet_avail_int              : in    std_logic;
          rx_CRC_error_int                 : in    std_logic;
          RESET                            : in    std_logic;
          rx_packet_complt                 : in    std_logic;
          rx_FIFO_UNDERRUN_int             : in    std_logic;
          RX_FIFO_rd_en                    : in    std_logic;
          rx_FIFO_OVERFLOW_int             : in    std_logic;
          RX_FIFO_Full                     : in    std_logic;
          RX_FIFO_Empty                    : in    std_logic;
          RX_packet_depth_status           : in    std_logic;
          tx_packet_complt                 : in    std_logic;
          TX_FIFO_wr_en                    : in    std_logic;
          TX_FIFO_Full                     : in    std_logic;
          m2s010_som_sb_0_GPIO_28_SW_RESET : in    std_logic;
          iup_EOP                          : in    std_logic;
          atrstb                           : in    std_logic;
          atms                             : in    std_logic;
          atdo                             : out   std_logic;
          atdi                             : in    std_logic;
          atck                             : in    std_logic
        );

end syn_identify_core0_0;

architecture DEF_ARCH of syn_identify_core0_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component IICE_x
    port( IICE_comm2iice                   : in    std_logic_vector(11 downto 0) := (others => 'U');
          up_EOP_del                       : in    std_logic_vector(5 downto 0) := (others => 'U');
          RX_FIFO_DIN                      : in    std_logic_vector(7 downto 0) := (others => 'U');
          RX_packet_depth                  : in    std_logic_vector(7 downto 0) := (others => 'U');
          RX_FIFO_DOUT                     : in    std_logic_vector(8 downto 0) := (others => 'U');
          un15                             : in    std_logic_vector(10 downto 0) := (others => 'U');
          ReadFIFO_Write_Ptr               : in    std_logic_vector(1 downto 0) := (others => 'U');
          RX_FIFO_DIN_pipe                 : in    std_logic_vector(8 downto 0) := (others => 'U');
          p2s_data                         : in    std_logic_vector(7 downto 0) := (others => 'U');
          packet_available_clear_reg       : in    std_logic_vector(2 downto 0) := (others => 'U');
          ReadFIFO_Read_Ptr                : in    std_logic_vector(1 downto 0) := (others => 'U');
          iRX_FIFO_UNDERRUN                : in    std_logic_vector(3 downto 0) := (others => 'U');
          int_reg                          : in    std_logic_vector(7 downto 1) := (others => 'U');
          iRX_FIFO_Empty                   : in    std_logic_vector(3 downto 0) := (others => 'U');
          iRX_FIFO_Full                    : in    std_logic_vector(3 downto 0) := (others => 'U');
          manches_in_dly                   : in    std_logic_vector(1 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PWDATA     : in    std_logic_vector(7 downto 0) := (others => 'U');
          clkdiv                           : in    std_logic_vector(3 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PADDR      : in    std_logic_vector(7 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PRDATA     : in    std_logic_vector(7 downto 0) := (others => 'U');
          un6                              : in    std_logic_vector(5 downto 0) := (others => 'U');
          control_reg_0                    : in    std_logic := 'U';
          control_reg_2                    : in    std_logic := 'U';
          control_reg_3                    : in    std_logic := 'U';
          IICE_iice2comm                   : out   std_logic;
          iup_EOP                          : in    std_logic := 'U';
          m2s010_som_sb_0_GPIO_28_SW_RESET : in    std_logic := 'U';
          TX_FIFO_Full                     : in    std_logic := 'U';
          TX_FIFO_wr_en                    : in    std_logic := 'U';
          tx_packet_complt                 : in    std_logic := 'U';
          RX_packet_depth_status           : in    std_logic := 'U';
          RX_FIFO_Empty                    : in    std_logic := 'U';
          RX_FIFO_Full                     : in    std_logic := 'U';
          rx_FIFO_OVERFLOW_int             : in    std_logic := 'U';
          RX_FIFO_rd_en                    : in    std_logic := 'U';
          rx_FIFO_UNDERRUN_int             : in    std_logic := 'U';
          rx_packet_complt                 : in    std_logic := 'U';
          RESET                            : in    std_logic := 'U';
          rx_CRC_error_int                 : in    std_logic := 'U';
          rx_packet_avail_int              : in    std_logic := 'U';
          TX_FIFO_Empty                    : in    std_logic := 'U';
          CommsFPGA_CCC_0_LOCK             : in    std_logic := 'U';
          MANCH_OUT_P_c                    : in    std_logic := 'U';
          MANCHESTER_IN_c                  : in    std_logic := 'U';
          int_reg_clr                      : in    std_logic := 'U';
          irx_center_sample                : in    std_logic := 'U';
          TX_FIFO_RST                      : in    std_logic := 'U';
          rx_FIFO_rst_reg                  : in    std_logic := 'U';
          start_tx_FIFO                    : in    std_logic := 'U';
          internal_loopback                : in    std_logic := 'U';
          external_loopback                : in    std_logic := 'U';
          iNRZ_data                        : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PWRITE     : in    std_logic := 'U';
          bd_reset                         : in    std_logic := 'U';
          m2s010_som_sb_0_POWER_ON_RESET_N : in    std_logic := 'U';
          block_int_until_rd               : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PREADY     : in    std_logic := 'U';
          long_reset                       : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0              : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component comm_block_x
    port( IICE_comm2iice : out   std_logic_vector(0 to 11);
          IICE_iice2comm : in    std_logic := 'U';
          atck           : in    std_logic := 'U';
          atdi           : in    std_logic := 'U';
          atdo           : out   std_logic;
          atms           : in    std_logic := 'U';
          atrstb         : in    std_logic := 'U'
        );
  end component;

    signal \IICE_comm2iice[11]\, \IICE_comm2iice[10]\, 
        \IICE_comm2iice[9]\, \IICE_comm2iice[8]\, 
        \IICE_comm2iice[7]\, \IICE_comm2iice[6]\, 
        \IICE_comm2iice[5]\, \IICE_comm2iice[4]\, 
        \IICE_comm2iice[3]\, \IICE_comm2iice[2]\, 
        \IICE_comm2iice[1]\, \IICE_comm2iice[0]\, IICE_iice2comm, 
        GND_net_1, VCC_net_1 : std_logic;
    signal nc2, nc1 : std_logic;

    for all : IICE_x
	Use entity work.IICE_x(DEF_ARCH);
    for all : comm_block_x
	Use entity work.comm_block_x(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    IICE_INST : IICE_x
      port map(IICE_comm2iice(11) => \IICE_comm2iice[11]\, 
        IICE_comm2iice(10) => \IICE_comm2iice[10]\, 
        IICE_comm2iice(9) => \IICE_comm2iice[9]\, 
        IICE_comm2iice(8) => \IICE_comm2iice[8]\, 
        IICE_comm2iice(7) => \IICE_comm2iice[7]\, 
        IICE_comm2iice(6) => \IICE_comm2iice[6]\, 
        IICE_comm2iice(5) => \IICE_comm2iice[5]\, 
        IICE_comm2iice(4) => \IICE_comm2iice[4]\, 
        IICE_comm2iice(3) => \IICE_comm2iice[3]\, 
        IICE_comm2iice(2) => \IICE_comm2iice[2]\, 
        IICE_comm2iice(1) => \IICE_comm2iice[1]\, 
        IICE_comm2iice(0) => \IICE_comm2iice[0]\, up_EOP_del(5)
         => up_EOP_del(5), up_EOP_del(4) => up_EOP_del(4), 
        up_EOP_del(3) => up_EOP_del(3), up_EOP_del(2) => 
        up_EOP_del(2), up_EOP_del(1) => up_EOP_del(1), 
        up_EOP_del(0) => up_EOP_del(0), RX_FIFO_DIN(7) => 
        RX_FIFO_DIN(7), RX_FIFO_DIN(6) => RX_FIFO_DIN(6), 
        RX_FIFO_DIN(5) => RX_FIFO_DIN(5), RX_FIFO_DIN(4) => 
        RX_FIFO_DIN(4), RX_FIFO_DIN(3) => RX_FIFO_DIN(3), 
        RX_FIFO_DIN(2) => RX_FIFO_DIN(2), RX_FIFO_DIN(1) => 
        RX_FIFO_DIN(1), RX_FIFO_DIN(0) => RX_FIFO_DIN(0), 
        RX_packet_depth(7) => RX_packet_depth(7), 
        RX_packet_depth(6) => RX_packet_depth(6), 
        RX_packet_depth(5) => RX_packet_depth(5), 
        RX_packet_depth(4) => RX_packet_depth(4), 
        RX_packet_depth(3) => RX_packet_depth(3), 
        RX_packet_depth(2) => RX_packet_depth(2), 
        RX_packet_depth(1) => RX_packet_depth(1), 
        RX_packet_depth(0) => RX_packet_depth(0), RX_FIFO_DOUT(8)
         => RX_FIFO_DOUT(8), RX_FIFO_DOUT(7) => RX_FIFO_DOUT(7), 
        RX_FIFO_DOUT(6) => RX_FIFO_DOUT(6), RX_FIFO_DOUT(5) => 
        RX_FIFO_DOUT(5), RX_FIFO_DOUT(4) => RX_FIFO_DOUT(4), 
        RX_FIFO_DOUT(3) => RX_FIFO_DOUT(3), RX_FIFO_DOUT(2) => 
        RX_FIFO_DOUT(2), RX_FIFO_DOUT(1) => RX_FIFO_DOUT(1), 
        RX_FIFO_DOUT(0) => RX_FIFO_DOUT(0), un15(10) => un15(10), 
        un15(9) => un15(9), un15(8) => un15(8), un15(7) => 
        un15(7), un15(6) => nc2, un15(5) => un15(5), un15(4) => 
        un15(4), un15(3) => un15(3), un15(2) => un15(2), un15(1)
         => un15(1), un15(0) => un15(0), ReadFIFO_Write_Ptr(1)
         => ReadFIFO_Write_Ptr(1), ReadFIFO_Write_Ptr(0) => 
        ReadFIFO_Write_Ptr(0), RX_FIFO_DIN_pipe(8) => 
        RX_FIFO_DIN_pipe(8), RX_FIFO_DIN_pipe(7) => 
        RX_FIFO_DIN_pipe(7), RX_FIFO_DIN_pipe(6) => 
        RX_FIFO_DIN_pipe(6), RX_FIFO_DIN_pipe(5) => 
        RX_FIFO_DIN_pipe(5), RX_FIFO_DIN_pipe(4) => 
        RX_FIFO_DIN_pipe(4), RX_FIFO_DIN_pipe(3) => 
        RX_FIFO_DIN_pipe(3), RX_FIFO_DIN_pipe(2) => 
        RX_FIFO_DIN_pipe(2), RX_FIFO_DIN_pipe(1) => 
        RX_FIFO_DIN_pipe(1), RX_FIFO_DIN_pipe(0) => 
        RX_FIFO_DIN_pipe(0), p2s_data(7) => p2s_data(7), 
        p2s_data(6) => p2s_data(6), p2s_data(5) => p2s_data(5), 
        p2s_data(4) => p2s_data(4), p2s_data(3) => p2s_data(3), 
        p2s_data(2) => p2s_data(2), p2s_data(1) => p2s_data(1), 
        p2s_data(0) => p2s_data(0), packet_available_clear_reg(2)
         => packet_available_clear_reg(2), 
        packet_available_clear_reg(1) => 
        packet_available_clear_reg(1), 
        packet_available_clear_reg(0) => 
        packet_available_clear_reg(0), ReadFIFO_Read_Ptr(1) => 
        ReadFIFO_Read_Ptr(1), ReadFIFO_Read_Ptr(0) => 
        ReadFIFO_Read_Ptr(0), iRX_FIFO_UNDERRUN(3) => 
        iRX_FIFO_UNDERRUN(3), iRX_FIFO_UNDERRUN(2) => 
        iRX_FIFO_UNDERRUN(2), iRX_FIFO_UNDERRUN(1) => 
        iRX_FIFO_UNDERRUN(1), iRX_FIFO_UNDERRUN(0) => 
        iRX_FIFO_UNDERRUN(0), int_reg(7) => int_reg(7), 
        int_reg(6) => int_reg(6), int_reg(5) => int_reg(5), 
        int_reg(4) => int_reg(4), int_reg(3) => int_reg(3), 
        int_reg(2) => int_reg(2), int_reg(1) => int_reg(1), 
        iRX_FIFO_Empty(3) => iRX_FIFO_Empty(3), iRX_FIFO_Empty(2)
         => iRX_FIFO_Empty(2), iRX_FIFO_Empty(1) => 
        iRX_FIFO_Empty(1), iRX_FIFO_Empty(0) => iRX_FIFO_Empty(0), 
        iRX_FIFO_Full(3) => iRX_FIFO_Full(3), iRX_FIFO_Full(2)
         => iRX_FIFO_Full(2), iRX_FIFO_Full(1) => 
        iRX_FIFO_Full(1), iRX_FIFO_Full(0) => iRX_FIFO_Full(0), 
        manches_in_dly(1) => manches_in_dly(1), manches_in_dly(0)
         => manches_in_dly(0), CoreAPB3_0_APBmslave0_PWDATA(7)
         => CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), clkdiv(3) => clkdiv(3), 
        clkdiv(2) => clkdiv(2), clkdiv(1) => clkdiv(1), clkdiv(0)
         => clkdiv(0), CoreAPB3_0_APBmslave0_PADDR(7) => 
        CoreAPB3_0_APBmslave0_PADDR(7), 
        CoreAPB3_0_APBmslave0_PADDR(6) => 
        CoreAPB3_0_APBmslave0_PADDR(6), 
        CoreAPB3_0_APBmslave0_PADDR(5) => 
        CoreAPB3_0_APBmslave0_PADDR(5), 
        CoreAPB3_0_APBmslave0_PADDR(4) => 
        CoreAPB3_0_APBmslave0_PADDR(4), 
        CoreAPB3_0_APBmslave0_PADDR(3) => 
        CoreAPB3_0_APBmslave0_PADDR(3), 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        CoreAPB3_0_APBmslave0_PADDR(2), 
        CoreAPB3_0_APBmslave0_PADDR(1) => 
        CoreAPB3_0_APBmslave0_PADDR(1), 
        CoreAPB3_0_APBmslave0_PADDR(0) => 
        CoreAPB3_0_APBmslave0_PADDR(0), 
        CoreAPB3_0_APBmslave0_PRDATA(7) => 
        CoreAPB3_0_APBmslave0_PRDATA(7), 
        CoreAPB3_0_APBmslave0_PRDATA(6) => 
        CoreAPB3_0_APBmslave0_PRDATA(6), 
        CoreAPB3_0_APBmslave0_PRDATA(5) => 
        CoreAPB3_0_APBmslave0_PRDATA(5), 
        CoreAPB3_0_APBmslave0_PRDATA(4) => 
        CoreAPB3_0_APBmslave0_PRDATA(4), 
        CoreAPB3_0_APBmslave0_PRDATA(3) => 
        CoreAPB3_0_APBmslave0_PRDATA(3), 
        CoreAPB3_0_APBmslave0_PRDATA(2) => 
        CoreAPB3_0_APBmslave0_PRDATA(2), 
        CoreAPB3_0_APBmslave0_PRDATA(1) => 
        CoreAPB3_0_APBmslave0_PRDATA(1), 
        CoreAPB3_0_APBmslave0_PRDATA(0) => 
        CoreAPB3_0_APBmslave0_PRDATA(0), un6(5) => un6(5), un6(4)
         => un6(4), un6(3) => un6(3), un6(2) => un6(2), un6(1)
         => nc1, un6(0) => un6(0), control_reg_0 => control_reg_0, 
        control_reg_2 => control_reg_2, control_reg_3 => 
        control_reg_3, IICE_iice2comm => IICE_iice2comm, iup_EOP
         => iup_EOP, m2s010_som_sb_0_GPIO_28_SW_RESET => 
        m2s010_som_sb_0_GPIO_28_SW_RESET, TX_FIFO_Full => 
        TX_FIFO_Full, TX_FIFO_wr_en => TX_FIFO_wr_en, 
        tx_packet_complt => tx_packet_complt, 
        RX_packet_depth_status => RX_packet_depth_status, 
        RX_FIFO_Empty => RX_FIFO_Empty, RX_FIFO_Full => 
        RX_FIFO_Full, rx_FIFO_OVERFLOW_int => 
        rx_FIFO_OVERFLOW_int, RX_FIFO_rd_en => RX_FIFO_rd_en, 
        rx_FIFO_UNDERRUN_int => rx_FIFO_UNDERRUN_int, 
        rx_packet_complt => rx_packet_complt, RESET => RESET, 
        rx_CRC_error_int => rx_CRC_error_int, rx_packet_avail_int
         => rx_packet_avail_int, TX_FIFO_Empty => TX_FIFO_Empty, 
        CommsFPGA_CCC_0_LOCK => CommsFPGA_CCC_0_LOCK, 
        MANCH_OUT_P_c => MANCH_OUT_P_c, MANCHESTER_IN_c => 
        MANCHESTER_IN_c, int_reg_clr => int_reg_clr, 
        irx_center_sample => irx_center_sample, TX_FIFO_RST => 
        TX_FIFO_RST, rx_FIFO_rst_reg => rx_FIFO_rst_reg, 
        start_tx_FIFO => start_tx_FIFO, internal_loopback => 
        internal_loopback, external_loopback => external_loopback, 
        iNRZ_data => iNRZ_data, CoreAPB3_0_APBmslave0_PWRITE => 
        CoreAPB3_0_APBmslave0_PWRITE, bd_reset => bd_reset, 
        m2s010_som_sb_0_POWER_ON_RESET_N => 
        m2s010_som_sb_0_POWER_ON_RESET_N, block_int_until_rd => 
        block_int_until_rd, CoreAPB3_0_APBmslave0_PREADY => 
        CoreAPB3_0_APBmslave0_PREADY, long_reset => long_reset, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    comm_block_INST : comm_block_x
      port map(IICE_comm2iice(0) => \IICE_comm2iice[0]\, 
        IICE_comm2iice(1) => \IICE_comm2iice[1]\, 
        IICE_comm2iice(2) => \IICE_comm2iice[2]\, 
        IICE_comm2iice(3) => \IICE_comm2iice[3]\, 
        IICE_comm2iice(4) => \IICE_comm2iice[4]\, 
        IICE_comm2iice(5) => \IICE_comm2iice[5]\, 
        IICE_comm2iice(6) => \IICE_comm2iice[6]\, 
        IICE_comm2iice(7) => \IICE_comm2iice[7]\, 
        IICE_comm2iice(8) => \IICE_comm2iice[8]\, 
        IICE_comm2iice(9) => \IICE_comm2iice[9]\, 
        IICE_comm2iice(10) => \IICE_comm2iice[10]\, 
        IICE_comm2iice(11) => \IICE_comm2iice[11]\, 
        IICE_iice2comm => IICE_iice2comm, atck => atck, atdi => 
        atdi, atdo => atdo, atms => atms, atrstb => atrstb);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreAPB3 is

    port( m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR : in    std_logic_vector(15 downto 12);
          CoreAPB3_0_APBmslave0_PSELx            : out   std_logic;
          m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx : in    std_logic
        );

end CoreAPB3;

architecture DEF_ARCH of CoreAPB3 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \iPSELS_raw_1[0]_net_1\, GND_net_1, VCC_net_1
         : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \iPSELS_raw_1[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(15), B
         => m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(14), Y => 
        \iPSELS_raw_1[0]_net_1\);
    
    \iPSELS_raw[0]\ : CFG4
      generic map(INIT => x"0008")

      port map(A => m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx, B => 
        \iPSELS_raw_1[0]_net_1\, C => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(13), D => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(12), Y => 
        CoreAPB3_0_APBmslave0_PSELx);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_CommsFPGA_CCC_0_FCCC is

    port( m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC : in    std_logic;
          CommsFPGA_CCC_0_LOCK                      : out   std_logic;
          CommsFPGA_CCC_0_GL1                       : out   std_logic;
          CommsFPGA_CCC_0_GL0                       : out   std_logic
        );

end m2s010_som_CommsFPGA_CCC_0_FCCC;

architecture DEF_ARCH of m2s010_som_CommsFPGA_CCC_0_FCCC is 

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CCC

            generic (INIT:std_logic_vector(209 downto 0) := "00" & x"0000000000000000000000000000000000000000000000000000"; 
        VCOFREQUENCY:real := 0.0);

    port( Y0              : out   std_logic;
          Y1              : out   std_logic;
          Y2              : out   std_logic;
          Y3              : out   std_logic;
          PRDATA          : out   std_logic_vector(7 downto 0);
          LOCK            : out   std_logic;
          BUSY            : out   std_logic;
          CLK0            : in    std_logic := 'U';
          CLK1            : in    std_logic := 'U';
          CLK2            : in    std_logic := 'U';
          CLK3            : in    std_logic := 'U';
          NGMUX0_SEL      : in    std_logic := 'U';
          NGMUX1_SEL      : in    std_logic := 'U';
          NGMUX2_SEL      : in    std_logic := 'U';
          NGMUX3_SEL      : in    std_logic := 'U';
          NGMUX0_HOLD_N   : in    std_logic := 'U';
          NGMUX1_HOLD_N   : in    std_logic := 'U';
          NGMUX2_HOLD_N   : in    std_logic := 'U';
          NGMUX3_HOLD_N   : in    std_logic := 'U';
          NGMUX0_ARST_N   : in    std_logic := 'U';
          NGMUX1_ARST_N   : in    std_logic := 'U';
          NGMUX2_ARST_N   : in    std_logic := 'U';
          NGMUX3_ARST_N   : in    std_logic := 'U';
          PLL_BYPASS_N    : in    std_logic := 'U';
          PLL_ARST_N      : in    std_logic := 'U';
          PLL_POWERDOWN_N : in    std_logic := 'U';
          GPD0_ARST_N     : in    std_logic := 'U';
          GPD1_ARST_N     : in    std_logic := 'U';
          GPD2_ARST_N     : in    std_logic := 'U';
          GPD3_ARST_N     : in    std_logic := 'U';
          PRESET_N        : in    std_logic := 'U';
          PCLK            : in    std_logic := 'U';
          PSEL            : in    std_logic := 'U';
          PENABLE         : in    std_logic := 'U';
          PWRITE          : in    std_logic := 'U';
          PADDR           : in    std_logic_vector(7 downto 2) := (others => 'U');
          PWDATA          : in    std_logic_vector(7 downto 0) := (others => 'U');
          CLK0_PAD        : in    std_logic := 'U';
          CLK1_PAD        : in    std_logic := 'U';
          CLK2_PAD        : in    std_logic := 'U';
          CLK3_PAD        : in    std_logic := 'U';
          GL0             : out   std_logic;
          GL1             : out   std_logic;
          GL2             : out   std_logic;
          GL3             : out   std_logic;
          RCOSC_25_50MHZ  : in    std_logic := 'U';
          RCOSC_1MHZ      : in    std_logic := 'U';
          XTLOSC          : in    std_logic := 'U'
        );
  end component;

    signal GL0_net, GL1_net, VCC_net_1, GND_net_1 : std_logic;
    signal nc8, nc7, nc6, nc2, nc5, nc4, nc3, nc1 : std_logic;

begin 


    GL1_INST : CLKINT
      port map(A => GL1_net, Y => CommsFPGA_CCC_0_GL1);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    GL0_INST : CLKINT
      port map(A => GL0_net, Y => CommsFPGA_CCC_0_GL0);
    
    CCC_INST : CCC

              generic map(INIT => "00" & x"000007FB8000044164000F18C6309C231839DE40404C41803000",
         VCOFREQUENCY => 980.0)

      port map(Y0 => OPEN, Y1 => OPEN, Y2 => OPEN, Y3 => OPEN, 
        PRDATA(7) => nc8, PRDATA(6) => nc7, PRDATA(5) => nc6, 
        PRDATA(4) => nc2, PRDATA(3) => nc5, PRDATA(2) => nc4, 
        PRDATA(1) => nc3, PRDATA(0) => nc1, LOCK => 
        CommsFPGA_CCC_0_LOCK, BUSY => OPEN, CLK0 => VCC_net_1, 
        CLK1 => VCC_net_1, CLK2 => VCC_net_1, CLK3 => VCC_net_1, 
        NGMUX0_SEL => GND_net_1, NGMUX1_SEL => GND_net_1, 
        NGMUX2_SEL => GND_net_1, NGMUX3_SEL => GND_net_1, 
        NGMUX0_HOLD_N => VCC_net_1, NGMUX1_HOLD_N => VCC_net_1, 
        NGMUX2_HOLD_N => VCC_net_1, NGMUX3_HOLD_N => VCC_net_1, 
        NGMUX0_ARST_N => VCC_net_1, NGMUX1_ARST_N => VCC_net_1, 
        NGMUX2_ARST_N => VCC_net_1, NGMUX3_ARST_N => VCC_net_1, 
        PLL_BYPASS_N => VCC_net_1, PLL_ARST_N => VCC_net_1, 
        PLL_POWERDOWN_N => VCC_net_1, GPD0_ARST_N => VCC_net_1, 
        GPD1_ARST_N => VCC_net_1, GPD2_ARST_N => VCC_net_1, 
        GPD3_ARST_N => VCC_net_1, PRESET_N => GND_net_1, PCLK => 
        VCC_net_1, PSEL => VCC_net_1, PENABLE => VCC_net_1, 
        PWRITE => VCC_net_1, PADDR(7) => VCC_net_1, PADDR(6) => 
        VCC_net_1, PADDR(5) => VCC_net_1, PADDR(4) => VCC_net_1, 
        PADDR(3) => VCC_net_1, PADDR(2) => VCC_net_1, PWDATA(7)
         => VCC_net_1, PWDATA(6) => VCC_net_1, PWDATA(5) => 
        VCC_net_1, PWDATA(4) => VCC_net_1, PWDATA(3) => VCC_net_1, 
        PWDATA(2) => VCC_net_1, PWDATA(1) => VCC_net_1, PWDATA(0)
         => VCC_net_1, CLK0_PAD => GND_net_1, CLK1_PAD => 
        GND_net_1, CLK2_PAD => GND_net_1, CLK3_PAD => GND_net_1, 
        GL0 => GL0_net, GL1 => GL1_net, GL2 => OPEN, GL3 => OPEN, 
        RCOSC_25_50MHZ => GND_net_1, RCOSC_1MHZ => GND_net_1, 
        XTLOSC => m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_ID_RES_0_IO is

    port( ID_RES  : in    std_logic_vector(3 downto 0);
          Y_net_0 : out   std_logic_vector(3 downto 0)
        );

end m2s010_som_ID_RES_0_IO;

architecture DEF_ARCH of m2s010_som_ID_RES_0_IO is 

  component INBUF
    generic (IOSTD:string := "");

    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    U0_0 : INBUF
      port map(PAD => ID_RES(0), Y => Y_net_0(0));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    U0_3 : INBUF
      port map(PAD => ID_RES(3), Y => Y_net_0(3));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    U0_2 : INBUF
      port map(PAD => ID_RES(2), Y => Y_net_0(2));
    
    U0_1 : INBUF
      port map(PAD => ID_RES(1), Y => Y_net_0(1));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb_GPIO_1_IO is

    port( GPIO_1_BI_0                       : inout std_logic := 'Z';
          GPIO_1_in_0                       : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_1_M2F_OE : in    std_logic;
          GPIO_1_M2F                        : in    std_logic
        );

end m2s010_som_sb_GPIO_1_IO;

architecture DEF_ARCH of m2s010_som_sb_GPIO_1_IO is 

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    U0_0 : BIBUF
      generic map(IOSTD => "LVCMOS33")

      port map(PAD => GPIO_1_BI_0, D => GPIO_1_M2F, E => 
        m2s010_som_sb_MSS_0_GPIO_1_M2F_OE, Y => GPIO_1_in_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb_CAM_SPI_1_CLK_IO is

    port( CAM_SPI_1_CLK_Y_0                    : out   std_logic;
          SPI_1_CLK_0                          : inout std_logic := 'Z';
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE : in    std_logic;
          m2s010_som_sb_MSS_0_SPI_1_CLK_M2F    : in    std_logic
        );

end m2s010_som_sb_CAM_SPI_1_CLK_IO;

architecture DEF_ARCH of m2s010_som_sb_CAM_SPI_1_CLK_IO is 

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    U0_0 : BIBUF
      port map(PAD => SPI_1_CLK_0, D => 
        m2s010_som_sb_MSS_0_SPI_1_CLK_M2F, E => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE, Y => 
        CAM_SPI_1_CLK_Y_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb_GPIO_7_IO is

    port( GPIO_7_PADI_0                     : inout std_logic := 'Z';
          GPIO_7_Y_0                        : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_7_M2F_OE : in    std_logic;
          m2s010_som_sb_MSS_0_GPIO_7_M2F    : in    std_logic
        );

end m2s010_som_sb_GPIO_7_IO;

architecture DEF_ARCH of m2s010_som_sb_GPIO_7_IO is 

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    U0_0 : BIBUF
      port map(PAD => GPIO_7_PADI_0, D => 
        m2s010_som_sb_MSS_0_GPIO_7_M2F, E => 
        m2s010_som_sb_MSS_0_GPIO_7_M2F_OE, Y => GPIO_7_Y_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb_CAM_SPI_1_SS0_IO is

    port( SPI_1_SS0_CAM_0                      : inout std_logic := 'Z';
          CAM_SPI_1_SS0_Y_0                    : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE : in    std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F    : in    std_logic
        );

end m2s010_som_sb_CAM_SPI_1_SS0_IO;

architecture DEF_ARCH of m2s010_som_sb_CAM_SPI_1_SS0_IO is 

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    U0_0 : BIBUF
      port map(PAD => SPI_1_SS0_CAM_0, D => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F, E => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE, Y => 
        CAM_SPI_1_SS0_Y_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb_MSS is

    port( CORECONFIGP_0_MDDR_APBmslave_PWDATA              : in    std_logic_vector(15 downto 0);
          CORECONFIGP_0_MDDR_APBmslave_PADDR               : in    std_logic_vector(10 downto 2);
          MAC_MII_RXD_c                                    : in    std_logic_vector(3 downto 0);
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA  : in    std_logic_vector(17 downto 0);
          Y_net_0                                          : in    std_logic_vector(3 downto 0);
          CoreAPB3_0_APBmslave0_PRDATA_m                   : in    std_logic_vector(7 downto 0);
          CORECONFIGP_0_MDDR_APBmslave_PRDATA              : out   std_logic_vector(15 downto 0);
          MAC_MII_TXD_c                                    : out   std_logic_vector(3 downto 0);
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA  : out   std_logic_vector(16 downto 0);
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR   : out   std_logic_vector(15 downto 2);
          CoreAPB3_0_APBmslave0_PWDATA                     : out   std_logic_vector(7 downto 0);
          m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR           : out   std_logic_vector(15 downto 12);
          CoreAPB3_0_APBmslave0_PADDR                      : out   std_logic_vector(7 downto 0);
          MDDR_ADDR                                        : out   std_logic_vector(15 downto 0);
          MDDR_BA                                          : out   std_logic_vector(2 downto 0);
          MDDR_DM_RDQS                                     : inout std_logic_vector(1 downto 0) := (others => 'Z');
          MDDR_DQ                                          : inout std_logic_vector(15 downto 0) := (others => 'Z');
          MDDR_DQS                                         : inout std_logic_vector(1 downto 0) := (others => 'Z');
          CAM_SPI_1_CLK_Y_0                                : in    std_logic;
          GPIO_7_Y_0                                       : in    std_logic;
          GPIO_6_Y_0                                       : in    std_logic;
          DEBOUNCE_OUT_net_0_0                             : in    std_logic;
          GPIO_1_in_0                                      : in    std_logic;
          MDDR_CLK                                         : out   std_logic;
          MDDR_CLK_N                                       : out   std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PWRITE              : in    std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PSELx               : in    std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PENABLE             : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz                        : in    std_logic;
          MAC_MII_TX_CLK_c                                 : in    std_logic;
          SPI_1_SS0_MX_Y                                   : in    std_logic;
          SPI_1_DI                                         : in    std_logic;
          MAC_MII_RX_ER_c                                  : in    std_logic;
          MAC_MII_RX_DV_c                                  : in    std_logic;
          MAC_MII_RX_CLK_c                                 : in    std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR : in    std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY  : in    std_logic;
          MMUART_0_RXD_F2M_c                               : in    std_logic;
          DEBOUNCE_OUT_2_c                                 : in    std_logic;
          DEBOUNCE_OUT_1_c                                 : in    std_logic;
          BIBUF_0_Y                                        : in    std_logic;
          FAB_CCC_LOCK                                     : in    std_logic;
          CoreAPB3_0_APBmslave0_PREADY_i_m_i               : in    std_logic;
          CommsFPGA_top_0_INT                              : in    std_logic;
          MAC_MII_CRS_c                                    : in    std_logic;
          MAC_MII_COL_c                                    : in    std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PSLVERR             : out   std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PREADY              : out   std_logic;
          MAC_MII_TX_EN_c                                  : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE             : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F                : out   std_logic;
          SPI_1_DO_CAM_c                                   : out   std_logic;
          GPIO_11_M2F_c                                    : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_CLK_M2F                : out   std_logic;
          GPIO_8_M2F_c                                     : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_7_M2F                   : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_7_M2F_OE                : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_6_M2F                   : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_6_M2F_OE                : out   std_logic;
          GPIO_5_M2F_c                                     : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE  : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx   : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE : out   std_logic;
          GPIO_24_M2F_c                                    : out   std_logic;
          MMUART_0_TXD_M2F_c                               : out   std_logic;
          m2s010_som_sb_0_GPIO_28_SW_RESET                 : out   std_logic;
          GPIO_21_M2F_c                                    : out   std_logic;
          GPIO_22_M2F_c                                    : out   std_logic;
          m2s010_som_sb_MSS_0_MAC_MII_MDO                  : out   std_logic;
          m2s010_som_sb_MSS_0_MAC_MII_MDO_EN               : out   std_logic;
          MAC_MII_MDC_c                                    : out   std_logic;
          GPIO_1_M2F                                       : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_1_M2F_OE                : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F          : out   std_logic;
          CoreAPB3_0_APBmslave0_PWRITE                     : out   std_logic;
          m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx           : out   std_logic;
          CoreAPB3_0_APBmslave0_PENABLE                    : out   std_logic;
          GPIO_0_BI                                        : inout std_logic := 'Z';
          GPIO_3_BI                                        : inout std_logic := 'Z';
          GPIO_4_BI                                        : inout std_logic := 'Z';
          GPIO_12_BI                                       : inout std_logic := 'Z';
          GPIO_14_BI                                       : inout std_logic := 'Z';
          GPIO_15_BI                                       : inout std_logic := 'Z';
          GPIO_16_BI                                       : inout std_logic := 'Z';
          GPIO_17_BI                                       : inout std_logic := 'Z';
          GPIO_18_BI                                       : inout std_logic := 'Z';
          GPIO_20_OUT                                      : out   std_logic;
          GPIO_25_BI                                       : inout std_logic := 'Z';
          GPIO_26_BI                                       : inout std_logic := 'Z';
          GPIO_31_BI                                       : inout std_logic := 'Z';
          I2C_1_SCL                                        : inout std_logic := 'Z';
          I2C_1_SDA                                        : inout std_logic := 'Z';
          MDDR_CAS_N                                       : out   std_logic;
          MDDR_CKE                                         : out   std_logic;
          MDDR_CS_N                                        : out   std_logic;
          MDDR_DQS_TMATCH_0_IN                             : in    std_logic;
          MDDR_DQS_TMATCH_0_OUT                            : out   std_logic;
          MDDR_ODT                                         : out   std_logic;
          MDDR_RAS_N                                       : out   std_logic;
          MDDR_RESET_N                                     : out   std_logic;
          MDDR_WE_N                                        : out   std_logic;
          MMUART_1_RXD                                     : in    std_logic;
          MMUART_1_TXD                                     : out   std_logic;
          SPI_0_CLK                                        : inout std_logic := 'Z';
          SPI_0_DI                                         : in    std_logic;
          SPI_0_DO                                         : out   std_logic;
          SPI_0_SS0                                        : inout std_logic := 'Z';
          SPI_0_SS1                                        : out   std_logic;
          CORECONFIGP_0_APB_S_PCLK_i                       : out   std_logic;
          CORECONFIGP_0_APB_S_PRESET_N                     : out   std_logic;
          CORECONFIGP_0_APB_S_PCLK                         : out   std_logic
        );

end m2s010_som_sb_MSS;

architecture DEF_ARCH of m2s010_som_sb_MSS is 

  component OUTBUF
    generic (IOSTD:string := "");

    port( D   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component TRIBUFF
    generic (IOSTD:string := "");

    port( D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component INBUF
    generic (IOSTD:string := "");

    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component MSS_060

            generic (INIT:std_logic_vector(1437 downto 0) := "00" & x"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"; 
        ACT_UBITS:std_logic_vector(55 downto 0) := x"FFFFFFFFFFFFFF"; 
        MEMORYFILE:string := ""; RTC_MAIN_XTL_FREQ:real := 0.0; 
        RTC_MAIN_XTL_MODE:string := "1"; DDR_CLK_FREQ:real := 0.0
        );

    port( CAN_RXBUS_MGPIO3A_H2F_A                 : out   std_logic;
          CAN_RXBUS_MGPIO3A_H2F_B                 : out   std_logic;
          CAN_TX_EBL_MGPIO4A_H2F_A                : out   std_logic;
          CAN_TX_EBL_MGPIO4A_H2F_B                : out   std_logic;
          CAN_TXBUS_MGPIO2A_H2F_A                 : out   std_logic;
          CAN_TXBUS_MGPIO2A_H2F_B                 : out   std_logic;
          CLK_CONFIG_APB                          : out   std_logic;
          COMMS_INT                               : out   std_logic;
          CONFIG_PRESET_N                         : out   std_logic;
          EDAC_ERROR                              : out   std_logic_vector(7 downto 0);
          F_FM0_RDATA                             : out   std_logic_vector(31 downto 0);
          F_FM0_READYOUT                          : out   std_logic;
          F_FM0_RESP                              : out   std_logic;
          F_HM0_ADDR                              : out   std_logic_vector(31 downto 0);
          F_HM0_ENABLE                            : out   std_logic;
          F_HM0_SEL                               : out   std_logic;
          F_HM0_SIZE                              : out   std_logic_vector(1 downto 0);
          F_HM0_TRANS1                            : out   std_logic;
          F_HM0_WDATA                             : out   std_logic_vector(31 downto 0);
          F_HM0_WRITE                             : out   std_logic;
          FAB_CHRGVBUS                            : out   std_logic;
          FAB_DISCHRGVBUS                         : out   std_logic;
          FAB_DMPULLDOWN                          : out   std_logic;
          FAB_DPPULLDOWN                          : out   std_logic;
          FAB_DRVVBUS                             : out   std_logic;
          FAB_IDPULLUP                            : out   std_logic;
          FAB_OPMODE                              : out   std_logic_vector(1 downto 0);
          FAB_SUSPENDM                            : out   std_logic;
          FAB_TERMSEL                             : out   std_logic;
          FAB_TXVALID                             : out   std_logic;
          FAB_VCONTROL                            : out   std_logic_vector(3 downto 0);
          FAB_VCONTROLLOADM                       : out   std_logic;
          FAB_XCVRSEL                             : out   std_logic_vector(1 downto 0);
          FAB_XDATAOUT                            : out   std_logic_vector(7 downto 0);
          FACC_GLMUX_SEL                          : out   std_logic;
          FIC32_0_MASTER                          : out   std_logic_vector(1 downto 0);
          FIC32_1_MASTER                          : out   std_logic_vector(1 downto 0);
          FPGA_RESET_N                            : out   std_logic;
          GTX_CLK                                 : out   std_logic;
          H2F_INTERRUPT                           : out   std_logic_vector(15 downto 0);
          H2F_NMI                                 : out   std_logic;
          H2FCALIB                                : out   std_logic;
          I2C0_SCL_MGPIO31B_H2F_A                 : out   std_logic;
          I2C0_SCL_MGPIO31B_H2F_B                 : out   std_logic;
          I2C0_SDA_MGPIO30B_H2F_A                 : out   std_logic;
          I2C0_SDA_MGPIO30B_H2F_B                 : out   std_logic;
          I2C1_SCL_MGPIO1A_H2F_A                  : out   std_logic;
          I2C1_SCL_MGPIO1A_H2F_B                  : out   std_logic;
          I2C1_SDA_MGPIO0A_H2F_A                  : out   std_logic;
          I2C1_SDA_MGPIO0A_H2F_B                  : out   std_logic;
          MDCF                                    : out   std_logic;
          MDOENF                                  : out   std_logic;
          MDOF                                    : out   std_logic;
          MMUART0_CTS_MGPIO19B_H2F_A              : out   std_logic;
          MMUART0_CTS_MGPIO19B_H2F_B              : out   std_logic;
          MMUART0_DCD_MGPIO22B_H2F_A              : out   std_logic;
          MMUART0_DCD_MGPIO22B_H2F_B              : out   std_logic;
          MMUART0_DSR_MGPIO20B_H2F_A              : out   std_logic;
          MMUART0_DSR_MGPIO20B_H2F_B              : out   std_logic;
          MMUART0_DTR_MGPIO18B_H2F_A              : out   std_logic;
          MMUART0_DTR_MGPIO18B_H2F_B              : out   std_logic;
          MMUART0_RI_MGPIO21B_H2F_A               : out   std_logic;
          MMUART0_RI_MGPIO21B_H2F_B               : out   std_logic;
          MMUART0_RTS_MGPIO17B_H2F_A              : out   std_logic;
          MMUART0_RTS_MGPIO17B_H2F_B              : out   std_logic;
          MMUART0_RXD_MGPIO28B_H2F_A              : out   std_logic;
          MMUART0_RXD_MGPIO28B_H2F_B              : out   std_logic;
          MMUART0_SCK_MGPIO29B_H2F_A              : out   std_logic;
          MMUART0_SCK_MGPIO29B_H2F_B              : out   std_logic;
          MMUART0_TXD_MGPIO27B_H2F_A              : out   std_logic;
          MMUART0_TXD_MGPIO27B_H2F_B              : out   std_logic;
          MMUART1_DTR_MGPIO12B_H2F_A              : out   std_logic;
          MMUART1_RTS_MGPIO11B_H2F_A              : out   std_logic;
          MMUART1_RTS_MGPIO11B_H2F_B              : out   std_logic;
          MMUART1_RXD_MGPIO26B_H2F_A              : out   std_logic;
          MMUART1_RXD_MGPIO26B_H2F_B              : out   std_logic;
          MMUART1_SCK_MGPIO25B_H2F_A              : out   std_logic;
          MMUART1_SCK_MGPIO25B_H2F_B              : out   std_logic;
          MMUART1_TXD_MGPIO24B_H2F_A              : out   std_logic;
          MMUART1_TXD_MGPIO24B_H2F_B              : out   std_logic;
          MPLL_LOCK                               : out   std_logic;
          PER2_FABRIC_PADDR                       : out   std_logic_vector(15 downto 2);
          PER2_FABRIC_PENABLE                     : out   std_logic;
          PER2_FABRIC_PSEL                        : out   std_logic;
          PER2_FABRIC_PWDATA                      : out   std_logic_vector(31 downto 0);
          PER2_FABRIC_PWRITE                      : out   std_logic;
          RTC_MATCH                               : out   std_logic;
          SLEEPDEEP                               : out   std_logic;
          SLEEPHOLDACK                            : out   std_logic;
          SLEEPING                                : out   std_logic;
          SMBALERT_NO0                            : out   std_logic;
          SMBALERT_NO1                            : out   std_logic;
          SMBSUS_NO0                              : out   std_logic;
          SMBSUS_NO1                              : out   std_logic;
          SPI0_CLK_OUT                            : out   std_logic;
          SPI0_SDI_MGPIO5A_H2F_A                  : out   std_logic;
          SPI0_SDI_MGPIO5A_H2F_B                  : out   std_logic;
          SPI0_SDO_MGPIO6A_H2F_A                  : out   std_logic;
          SPI0_SDO_MGPIO6A_H2F_B                  : out   std_logic;
          SPI0_SS0_MGPIO7A_H2F_A                  : out   std_logic;
          SPI0_SS0_MGPIO7A_H2F_B                  : out   std_logic;
          SPI0_SS1_MGPIO8A_H2F_A                  : out   std_logic;
          SPI0_SS1_MGPIO8A_H2F_B                  : out   std_logic;
          SPI0_SS2_MGPIO9A_H2F_A                  : out   std_logic;
          SPI0_SS2_MGPIO9A_H2F_B                  : out   std_logic;
          SPI0_SS3_MGPIO10A_H2F_A                 : out   std_logic;
          SPI0_SS3_MGPIO10A_H2F_B                 : out   std_logic;
          SPI0_SS4_MGPIO19A_H2F_A                 : out   std_logic;
          SPI0_SS5_MGPIO20A_H2F_A                 : out   std_logic;
          SPI0_SS6_MGPIO21A_H2F_A                 : out   std_logic;
          SPI0_SS7_MGPIO22A_H2F_A                 : out   std_logic;
          SPI1_CLK_OUT                            : out   std_logic;
          SPI1_SDI_MGPIO11A_H2F_A                 : out   std_logic;
          SPI1_SDI_MGPIO11A_H2F_B                 : out   std_logic;
          SPI1_SDO_MGPIO12A_H2F_A                 : out   std_logic;
          SPI1_SDO_MGPIO12A_H2F_B                 : out   std_logic;
          SPI1_SS0_MGPIO13A_H2F_A                 : out   std_logic;
          SPI1_SS0_MGPIO13A_H2F_B                 : out   std_logic;
          SPI1_SS1_MGPIO14A_H2F_A                 : out   std_logic;
          SPI1_SS1_MGPIO14A_H2F_B                 : out   std_logic;
          SPI1_SS2_MGPIO15A_H2F_A                 : out   std_logic;
          SPI1_SS2_MGPIO15A_H2F_B                 : out   std_logic;
          SPI1_SS3_MGPIO16A_H2F_A                 : out   std_logic;
          SPI1_SS3_MGPIO16A_H2F_B                 : out   std_logic;
          SPI1_SS4_MGPIO17A_H2F_A                 : out   std_logic;
          SPI1_SS5_MGPIO18A_H2F_A                 : out   std_logic;
          SPI1_SS6_MGPIO23A_H2F_A                 : out   std_logic;
          SPI1_SS7_MGPIO24A_H2F_A                 : out   std_logic;
          TCGF                                    : out   std_logic_vector(9 downto 0);
          TRACECLK                                : out   std_logic;
          TRACEDATA                               : out   std_logic_vector(3 downto 0);
          TX_CLK                                  : out   std_logic;
          TX_ENF                                  : out   std_logic;
          TX_ERRF                                 : out   std_logic;
          TXCTL_EN_RIF                            : out   std_logic;
          TXD_RIF                                 : out   std_logic_vector(3 downto 0);
          TXDF                                    : out   std_logic_vector(7 downto 0);
          TXEV                                    : out   std_logic;
          WDOGTIMEOUT                             : out   std_logic;
          F_ARREADY_HREADYOUT1                    : out   std_logic;
          F_AWREADY_HREADYOUT0                    : out   std_logic;
          F_BID                                   : out   std_logic_vector(3 downto 0);
          F_BRESP_HRESP0                          : out   std_logic_vector(1 downto 0);
          F_BVALID                                : out   std_logic;
          F_RDATA_HRDATA01                        : out   std_logic_vector(63 downto 0);
          F_RID                                   : out   std_logic_vector(3 downto 0);
          F_RLAST                                 : out   std_logic;
          F_RRESP_HRESP1                          : out   std_logic_vector(1 downto 0);
          F_RVALID                                : out   std_logic;
          F_WREADY                                : out   std_logic;
          MDDR_FABRIC_PRDATA                      : out   std_logic_vector(15 downto 0);
          MDDR_FABRIC_PREADY                      : out   std_logic;
          MDDR_FABRIC_PSLVERR                     : out   std_logic;
          CAN_RXBUS_F2H_SCP                       : in    std_logic := 'U';
          CAN_TX_EBL_F2H_SCP                      : in    std_logic := 'U';
          CAN_TXBUS_F2H_SCP                       : in    std_logic := 'U';
          COLF                                    : in    std_logic := 'U';
          CRSF                                    : in    std_logic := 'U';
          F2_DMAREADY                             : in    std_logic_vector(1 downto 0) := (others => 'U');
          F2H_INTERRUPT                           : in    std_logic_vector(15 downto 0) := (others => 'U');
          F2HCALIB                                : in    std_logic := 'U';
          F_DMAREADY                              : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_FM0_ADDR                              : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_FM0_ENABLE                            : in    std_logic := 'U';
          F_FM0_MASTLOCK                          : in    std_logic := 'U';
          F_FM0_READY                             : in    std_logic := 'U';
          F_FM0_SEL                               : in    std_logic := 'U';
          F_FM0_SIZE                              : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_FM0_TRANS1                            : in    std_logic := 'U';
          F_FM0_WDATA                             : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_FM0_WRITE                             : in    std_logic := 'U';
          F_HM0_RDATA                             : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_HM0_READY                             : in    std_logic := 'U';
          F_HM0_RESP                              : in    std_logic := 'U';
          FAB_AVALID                              : in    std_logic := 'U';
          FAB_HOSTDISCON                          : in    std_logic := 'U';
          FAB_IDDIG                               : in    std_logic := 'U';
          FAB_LINESTATE                           : in    std_logic_vector(1 downto 0) := (others => 'U');
          FAB_M3_RESET_N                          : in    std_logic := 'U';
          FAB_PLL_LOCK                            : in    std_logic := 'U';
          FAB_RXACTIVE                            : in    std_logic := 'U';
          FAB_RXERROR                             : in    std_logic := 'U';
          FAB_RXVALID                             : in    std_logic := 'U';
          FAB_RXVALIDH                            : in    std_logic := 'U';
          FAB_SESSEND                             : in    std_logic := 'U';
          FAB_TXREADY                             : in    std_logic := 'U';
          FAB_VBUSVALID                           : in    std_logic := 'U';
          FAB_VSTATUS                             : in    std_logic_vector(7 downto 0) := (others => 'U');
          FAB_XDATAIN                             : in    std_logic_vector(7 downto 0) := (others => 'U');
          GTX_CLKPF                               : in    std_logic := 'U';
          I2C0_BCLK                               : in    std_logic := 'U';
          I2C0_SCL_F2H_SCP                        : in    std_logic := 'U';
          I2C0_SDA_F2H_SCP                        : in    std_logic := 'U';
          I2C1_BCLK                               : in    std_logic := 'U';
          I2C1_SCL_F2H_SCP                        : in    std_logic := 'U';
          I2C1_SDA_F2H_SCP                        : in    std_logic := 'U';
          MDIF                                    : in    std_logic := 'U';
          MGPIO0A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO10A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO11A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO11B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO12A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO13A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO14A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO15A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO16A_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO17B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO18B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO19B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO1A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO20B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO21B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO22B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO24B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO25B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO26B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO27B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO28B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO29B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO2A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO30B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO31B_F2H_GPIN                       : in    std_logic := 'U';
          MGPIO3A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO4A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO5A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO6A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO7A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO8A_F2H_GPIN                        : in    std_logic := 'U';
          MGPIO9A_F2H_GPIN                        : in    std_logic := 'U';
          MMUART0_CTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DCD_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DSR_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_DTR_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_RI_F2H_SCP                      : in    std_logic := 'U';
          MMUART0_RTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_RXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_SCK_F2H_SCP                     : in    std_logic := 'U';
          MMUART0_TXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_CTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_DCD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_DSR_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_RI_F2H_SCP                      : in    std_logic := 'U';
          MMUART1_RTS_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_RXD_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_SCK_F2H_SCP                     : in    std_logic := 'U';
          MMUART1_TXD_F2H_SCP                     : in    std_logic := 'U';
          PER2_FABRIC_PRDATA                      : in    std_logic_vector(31 downto 0) := (others => 'U');
          PER2_FABRIC_PREADY                      : in    std_logic := 'U';
          PER2_FABRIC_PSLVERR                     : in    std_logic := 'U';
          RCGF                                    : in    std_logic_vector(9 downto 0) := (others => 'U');
          RX_CLKPF                                : in    std_logic := 'U';
          RX_DVF                                  : in    std_logic := 'U';
          RX_ERRF                                 : in    std_logic := 'U';
          RX_EV                                   : in    std_logic := 'U';
          RXDF                                    : in    std_logic_vector(7 downto 0) := (others => 'U');
          SLEEPHOLDREQ                            : in    std_logic := 'U';
          SMBALERT_NI0                            : in    std_logic := 'U';
          SMBALERT_NI1                            : in    std_logic := 'U';
          SMBSUS_NI0                              : in    std_logic := 'U';
          SMBSUS_NI1                              : in    std_logic := 'U';
          SPI0_CLK_IN                             : in    std_logic := 'U';
          SPI0_SDI_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SDO_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS0_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS1_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS2_F2H_SCP                        : in    std_logic := 'U';
          SPI0_SS3_F2H_SCP                        : in    std_logic := 'U';
          SPI1_CLK_IN                             : in    std_logic := 'U';
          SPI1_SDI_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SDO_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS0_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS1_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS2_F2H_SCP                        : in    std_logic := 'U';
          SPI1_SS3_F2H_SCP                        : in    std_logic := 'U';
          TX_CLKPF                                : in    std_logic := 'U';
          USER_MSS_GPIO_RESET_N                   : in    std_logic := 'U';
          USER_MSS_RESET_N                        : in    std_logic := 'U';
          XCLK_FAB                                : in    std_logic := 'U';
          CLK_BASE                                : in    std_logic := 'U';
          CLK_MDDR_APB                            : in    std_logic := 'U';
          F_ARADDR_HADDR1                         : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_ARBURST_HTRANS1                       : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARID_HSEL1                            : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_ARLEN_HBURST1                         : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_ARLOCK_HMASTLOCK1                     : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARSIZE_HSIZE1                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_ARVALID_HWRITE1                       : in    std_logic := 'U';
          F_AWADDR_HADDR0                         : in    std_logic_vector(31 downto 0) := (others => 'U');
          F_AWBURST_HTRANS0                       : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWID_HSEL0                            : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_AWLEN_HBURST0                         : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_AWLOCK_HMASTLOCK0                     : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWSIZE_HSIZE0                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          F_AWVALID_HWRITE0                       : in    std_logic := 'U';
          F_BREADY                                : in    std_logic := 'U';
          F_RMW_AXI                               : in    std_logic := 'U';
          F_RREADY                                : in    std_logic := 'U';
          F_WDATA_HWDATA01                        : in    std_logic_vector(63 downto 0) := (others => 'U');
          F_WID_HREADY01                          : in    std_logic_vector(3 downto 0) := (others => 'U');
          F_WLAST                                 : in    std_logic := 'U';
          F_WSTRB                                 : in    std_logic_vector(7 downto 0) := (others => 'U');
          F_WVALID                                : in    std_logic := 'U';
          FPGA_MDDR_ARESET_N                      : in    std_logic := 'U';
          MDDR_FABRIC_PADDR                       : in    std_logic_vector(10 downto 2) := (others => 'U');
          MDDR_FABRIC_PENABLE                     : in    std_logic := 'U';
          MDDR_FABRIC_PSEL                        : in    std_logic := 'U';
          MDDR_FABRIC_PWDATA                      : in    std_logic_vector(15 downto 0) := (others => 'U');
          MDDR_FABRIC_PWRITE                      : in    std_logic := 'U';
          PRESET_N                                : in    std_logic := 'U';
          CAN_RXBUS_USBA_DATA1_MGPIO3A_IN         : in    std_logic := 'U';
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN        : in    std_logic := 'U';
          CAN_TXBUS_USBA_DATA0_MGPIO2A_IN         : in    std_logic := 'U';
          DM_IN                                   : in    std_logic_vector(2 downto 0) := (others => 'U');
          DRAM_DQ_IN                              : in    std_logic_vector(17 downto 0) := (others => 'U');
          DRAM_DQS_IN                             : in    std_logic_vector(2 downto 0) := (others => 'U');
          DRAM_FIFO_WE_IN                         : in    std_logic_vector(1 downto 0) := (others => 'U');
          I2C0_SCL_USBC_DATA1_MGPIO31B_IN         : in    std_logic := 'U';
          I2C0_SDA_USBC_DATA0_MGPIO30B_IN         : in    std_logic := 'U';
          I2C1_SCL_USBA_DATA4_MGPIO1A_IN          : in    std_logic := 'U';
          I2C1_SDA_USBA_DATA3_MGPIO0A_IN          : in    std_logic := 'U';
          MGPIO0B_IN                              : in    std_logic := 'U';
          MGPIO10B_IN                             : in    std_logic := 'U';
          MGPIO1B_IN                              : in    std_logic := 'U';
          MGPIO25A_IN                             : in    std_logic := 'U';
          MGPIO26A_IN                             : in    std_logic := 'U';
          MGPIO27A_IN                             : in    std_logic := 'U';
          MGPIO28A_IN                             : in    std_logic := 'U';
          MGPIO29A_IN                             : in    std_logic := 'U';
          MGPIO2B_IN                              : in    std_logic := 'U';
          MGPIO30A_IN                             : in    std_logic := 'U';
          MGPIO31A_IN                             : in    std_logic := 'U';
          MGPIO3B_IN                              : in    std_logic := 'U';
          MGPIO4B_IN                              : in    std_logic := 'U';
          MGPIO5B_IN                              : in    std_logic := 'U';
          MGPIO6B_IN                              : in    std_logic := 'U';
          MGPIO7B_IN                              : in    std_logic := 'U';
          MGPIO8B_IN                              : in    std_logic := 'U';
          MGPIO9B_IN                              : in    std_logic := 'U';
          MMUART0_CTS_USBC_DATA7_MGPIO19B_IN      : in    std_logic := 'U';
          MMUART0_DCD_MGPIO22B_IN                 : in    std_logic := 'U';
          MMUART0_DSR_MGPIO20B_IN                 : in    std_logic := 'U';
          MMUART0_DTR_USBC_DATA6_MGPIO18B_IN      : in    std_logic := 'U';
          MMUART0_RI_MGPIO21B_IN                  : in    std_logic := 'U';
          MMUART0_RTS_USBC_DATA5_MGPIO17B_IN      : in    std_logic := 'U';
          MMUART0_RXD_USBC_STP_MGPIO28B_IN        : in    std_logic := 'U';
          MMUART0_SCK_USBC_NXT_MGPIO29B_IN        : in    std_logic := 'U';
          MMUART0_TXD_USBC_DIR_MGPIO27B_IN        : in    std_logic := 'U';
          MMUART1_CTS_MGPIO13B_IN                 : in    std_logic := 'U';
          MMUART1_DCD_MGPIO16B_IN                 : in    std_logic := 'U';
          MMUART1_DSR_MGPIO14B_IN                 : in    std_logic := 'U';
          MMUART1_DTR_MGPIO12B_IN                 : in    std_logic := 'U';
          MMUART1_RI_MGPIO15B_IN                  : in    std_logic := 'U';
          MMUART1_RTS_MGPIO11B_IN                 : in    std_logic := 'U';
          MMUART1_RXD_USBC_DATA3_MGPIO26B_IN      : in    std_logic := 'U';
          MMUART1_SCK_USBC_DATA4_MGPIO25B_IN      : in    std_logic := 'U';
          MMUART1_TXD_USBC_DATA2_MGPIO24B_IN      : in    std_logic := 'U';
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN     : in    std_logic := 'U';
          RGMII_MDC_RMII_MDC_IN                   : in    std_logic := 'U';
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN      : in    std_logic := 'U';
          RGMII_RX_CLK_IN                         : in    std_logic := 'U';
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN  : in    std_logic := 'U';
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN      : in    std_logic := 'U';
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN      : in    std_logic := 'U';
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN     : in    std_logic := 'U';
          RGMII_RXD3_USBB_DATA4_IN                : in    std_logic := 'U';
          RGMII_TX_CLK_IN                         : in    std_logic := 'U';
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN     : in    std_logic := 'U';
          RGMII_TXD0_RMII_TXD0_USBB_DIR_IN        : in    std_logic := 'U';
          RGMII_TXD1_RMII_TXD1_USBB_STP_IN        : in    std_logic := 'U';
          RGMII_TXD2_USBB_DATA5_IN                : in    std_logic := 'U';
          RGMII_TXD3_USBB_DATA6_IN                : in    std_logic := 'U';
          SPI0_SCK_USBA_XCLK_IN                   : in    std_logic := 'U';
          SPI0_SDI_USBA_DIR_MGPIO5A_IN            : in    std_logic := 'U';
          SPI0_SDO_USBA_STP_MGPIO6A_IN            : in    std_logic := 'U';
          SPI0_SS0_USBA_NXT_MGPIO7A_IN            : in    std_logic := 'U';
          SPI0_SS1_USBA_DATA5_MGPIO8A_IN          : in    std_logic := 'U';
          SPI0_SS2_USBA_DATA6_MGPIO9A_IN          : in    std_logic := 'U';
          SPI0_SS3_USBA_DATA7_MGPIO10A_IN         : in    std_logic := 'U';
          SPI0_SS4_MGPIO19A_IN                    : in    std_logic := 'U';
          SPI0_SS5_MGPIO20A_IN                    : in    std_logic := 'U';
          SPI0_SS6_MGPIO21A_IN                    : in    std_logic := 'U';
          SPI0_SS7_MGPIO22A_IN                    : in    std_logic := 'U';
          SPI1_SCK_IN                             : in    std_logic := 'U';
          SPI1_SDI_MGPIO11A_IN                    : in    std_logic := 'U';
          SPI1_SDO_MGPIO12A_IN                    : in    std_logic := 'U';
          SPI1_SS0_MGPIO13A_IN                    : in    std_logic := 'U';
          SPI1_SS1_MGPIO14A_IN                    : in    std_logic := 'U';
          SPI1_SS2_MGPIO15A_IN                    : in    std_logic := 'U';
          SPI1_SS3_MGPIO16A_IN                    : in    std_logic := 'U';
          SPI1_SS4_MGPIO17A_IN                    : in    std_logic := 'U';
          SPI1_SS5_MGPIO18A_IN                    : in    std_logic := 'U';
          SPI1_SS6_MGPIO23A_IN                    : in    std_logic := 'U';
          SPI1_SS7_MGPIO24A_IN                    : in    std_logic := 'U';
          USBC_XCLK_IN                            : in    std_logic := 'U';
          USBD_DATA0_IN                           : in    std_logic := 'U';
          USBD_DATA1_IN                           : in    std_logic := 'U';
          USBD_DATA2_IN                           : in    std_logic := 'U';
          USBD_DATA3_IN                           : in    std_logic := 'U';
          USBD_DATA4_IN                           : in    std_logic := 'U';
          USBD_DATA5_IN                           : in    std_logic := 'U';
          USBD_DATA6_IN                           : in    std_logic := 'U';
          USBD_DATA7_MGPIO23B_IN                  : in    std_logic := 'U';
          USBD_DIR_IN                             : in    std_logic := 'U';
          USBD_NXT_IN                             : in    std_logic := 'U';
          USBD_STP_IN                             : in    std_logic := 'U';
          USBD_XCLK_IN                            : in    std_logic := 'U';
          CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT        : out   std_logic;
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT       : out   std_logic;
          CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT        : out   std_logic;
          DRAM_ADDR                               : out   std_logic_vector(15 downto 0);
          DRAM_BA                                 : out   std_logic_vector(2 downto 0);
          DRAM_CASN                               : out   std_logic;
          DRAM_CKE                                : out   std_logic;
          DRAM_CLK                                : out   std_logic;
          DRAM_CSN                                : out   std_logic;
          DRAM_DM_RDQS_OUT                        : out   std_logic_vector(2 downto 0);
          DRAM_DQ_OUT                             : out   std_logic_vector(17 downto 0);
          DRAM_DQS_OUT                            : out   std_logic_vector(2 downto 0);
          DRAM_FIFO_WE_OUT                        : out   std_logic_vector(1 downto 0);
          DRAM_ODT                                : out   std_logic;
          DRAM_RASN                               : out   std_logic;
          DRAM_RSTN                               : out   std_logic;
          DRAM_WEN                                : out   std_logic;
          I2C0_SCL_USBC_DATA1_MGPIO31B_OUT        : out   std_logic;
          I2C0_SDA_USBC_DATA0_MGPIO30B_OUT        : out   std_logic;
          I2C1_SCL_USBA_DATA4_MGPIO1A_OUT         : out   std_logic;
          I2C1_SDA_USBA_DATA3_MGPIO0A_OUT         : out   std_logic;
          MGPIO0B_OUT                             : out   std_logic;
          MGPIO10B_OUT                            : out   std_logic;
          MGPIO1B_OUT                             : out   std_logic;
          MGPIO25A_OUT                            : out   std_logic;
          MGPIO26A_OUT                            : out   std_logic;
          MGPIO27A_OUT                            : out   std_logic;
          MGPIO28A_OUT                            : out   std_logic;
          MGPIO29A_OUT                            : out   std_logic;
          MGPIO2B_OUT                             : out   std_logic;
          MGPIO30A_OUT                            : out   std_logic;
          MGPIO31A_OUT                            : out   std_logic;
          MGPIO3B_OUT                             : out   std_logic;
          MGPIO4B_OUT                             : out   std_logic;
          MGPIO5B_OUT                             : out   std_logic;
          MGPIO6B_OUT                             : out   std_logic;
          MGPIO7B_OUT                             : out   std_logic;
          MGPIO8B_OUT                             : out   std_logic;
          MGPIO9B_OUT                             : out   std_logic;
          MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT     : out   std_logic;
          MMUART0_DCD_MGPIO22B_OUT                : out   std_logic;
          MMUART0_DSR_MGPIO20B_OUT                : out   std_logic;
          MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT     : out   std_logic;
          MMUART0_RI_MGPIO21B_OUT                 : out   std_logic;
          MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT     : out   std_logic;
          MMUART0_RXD_USBC_STP_MGPIO28B_OUT       : out   std_logic;
          MMUART0_SCK_USBC_NXT_MGPIO29B_OUT       : out   std_logic;
          MMUART0_TXD_USBC_DIR_MGPIO27B_OUT       : out   std_logic;
          MMUART1_CTS_MGPIO13B_OUT                : out   std_logic;
          MMUART1_DCD_MGPIO16B_OUT                : out   std_logic;
          MMUART1_DSR_MGPIO14B_OUT                : out   std_logic;
          MMUART1_DTR_MGPIO12B_OUT                : out   std_logic;
          MMUART1_RI_MGPIO15B_OUT                 : out   std_logic;
          MMUART1_RTS_MGPIO11B_OUT                : out   std_logic;
          MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT     : out   std_logic;
          MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT     : out   std_logic;
          MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT     : out   std_logic;
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT    : out   std_logic;
          RGMII_MDC_RMII_MDC_OUT                  : out   std_logic;
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT     : out   std_logic;
          RGMII_RX_CLK_OUT                        : out   std_logic;
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT : out   std_logic;
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT     : out   std_logic;
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT     : out   std_logic;
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT    : out   std_logic;
          RGMII_RXD3_USBB_DATA4_OUT               : out   std_logic;
          RGMII_TX_CLK_OUT                        : out   std_logic;
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT    : out   std_logic;
          RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT       : out   std_logic;
          RGMII_TXD1_RMII_TXD1_USBB_STP_OUT       : out   std_logic;
          RGMII_TXD2_USBB_DATA5_OUT               : out   std_logic;
          RGMII_TXD3_USBB_DATA6_OUT               : out   std_logic;
          SPI0_SCK_USBA_XCLK_OUT                  : out   std_logic;
          SPI0_SDI_USBA_DIR_MGPIO5A_OUT           : out   std_logic;
          SPI0_SDO_USBA_STP_MGPIO6A_OUT           : out   std_logic;
          SPI0_SS0_USBA_NXT_MGPIO7A_OUT           : out   std_logic;
          SPI0_SS1_USBA_DATA5_MGPIO8A_OUT         : out   std_logic;
          SPI0_SS2_USBA_DATA6_MGPIO9A_OUT         : out   std_logic;
          SPI0_SS3_USBA_DATA7_MGPIO10A_OUT        : out   std_logic;
          SPI0_SS4_MGPIO19A_OUT                   : out   std_logic;
          SPI0_SS5_MGPIO20A_OUT                   : out   std_logic;
          SPI0_SS6_MGPIO21A_OUT                   : out   std_logic;
          SPI0_SS7_MGPIO22A_OUT                   : out   std_logic;
          SPI1_SCK_OUT                            : out   std_logic;
          SPI1_SDI_MGPIO11A_OUT                   : out   std_logic;
          SPI1_SDO_MGPIO12A_OUT                   : out   std_logic;
          SPI1_SS0_MGPIO13A_OUT                   : out   std_logic;
          SPI1_SS1_MGPIO14A_OUT                   : out   std_logic;
          SPI1_SS2_MGPIO15A_OUT                   : out   std_logic;
          SPI1_SS3_MGPIO16A_OUT                   : out   std_logic;
          SPI1_SS4_MGPIO17A_OUT                   : out   std_logic;
          SPI1_SS5_MGPIO18A_OUT                   : out   std_logic;
          SPI1_SS6_MGPIO23A_OUT                   : out   std_logic;
          SPI1_SS7_MGPIO24A_OUT                   : out   std_logic;
          USBC_XCLK_OUT                           : out   std_logic;
          USBD_DATA0_OUT                          : out   std_logic;
          USBD_DATA1_OUT                          : out   std_logic;
          USBD_DATA2_OUT                          : out   std_logic;
          USBD_DATA3_OUT                          : out   std_logic;
          USBD_DATA4_OUT                          : out   std_logic;
          USBD_DATA5_OUT                          : out   std_logic;
          USBD_DATA6_OUT                          : out   std_logic;
          USBD_DATA7_MGPIO23B_OUT                 : out   std_logic;
          USBD_DIR_OUT                            : out   std_logic;
          USBD_NXT_OUT                            : out   std_logic;
          USBD_STP_OUT                            : out   std_logic;
          USBD_XCLK_OUT                           : out   std_logic;
          CAN_RXBUS_USBA_DATA1_MGPIO3A_OE         : out   std_logic;
          CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE        : out   std_logic;
          CAN_TXBUS_USBA_DATA0_MGPIO2A_OE         : out   std_logic;
          DM_OE                                   : out   std_logic_vector(2 downto 0);
          DRAM_DQ_OE                              : out   std_logic_vector(17 downto 0);
          DRAM_DQS_OE                             : out   std_logic_vector(2 downto 0);
          I2C0_SCL_USBC_DATA1_MGPIO31B_OE         : out   std_logic;
          I2C0_SDA_USBC_DATA0_MGPIO30B_OE         : out   std_logic;
          I2C1_SCL_USBA_DATA4_MGPIO1A_OE          : out   std_logic;
          I2C1_SDA_USBA_DATA3_MGPIO0A_OE          : out   std_logic;
          MGPIO0B_OE                              : out   std_logic;
          MGPIO10B_OE                             : out   std_logic;
          MGPIO1B_OE                              : out   std_logic;
          MGPIO25A_OE                             : out   std_logic;
          MGPIO26A_OE                             : out   std_logic;
          MGPIO27A_OE                             : out   std_logic;
          MGPIO28A_OE                             : out   std_logic;
          MGPIO29A_OE                             : out   std_logic;
          MGPIO2B_OE                              : out   std_logic;
          MGPIO30A_OE                             : out   std_logic;
          MGPIO31A_OE                             : out   std_logic;
          MGPIO3B_OE                              : out   std_logic;
          MGPIO4B_OE                              : out   std_logic;
          MGPIO5B_OE                              : out   std_logic;
          MGPIO6B_OE                              : out   std_logic;
          MGPIO7B_OE                              : out   std_logic;
          MGPIO8B_OE                              : out   std_logic;
          MGPIO9B_OE                              : out   std_logic;
          MMUART0_CTS_USBC_DATA7_MGPIO19B_OE      : out   std_logic;
          MMUART0_DCD_MGPIO22B_OE                 : out   std_logic;
          MMUART0_DSR_MGPIO20B_OE                 : out   std_logic;
          MMUART0_DTR_USBC_DATA6_MGPIO18B_OE      : out   std_logic;
          MMUART0_RI_MGPIO21B_OE                  : out   std_logic;
          MMUART0_RTS_USBC_DATA5_MGPIO17B_OE      : out   std_logic;
          MMUART0_RXD_USBC_STP_MGPIO28B_OE        : out   std_logic;
          MMUART0_SCK_USBC_NXT_MGPIO29B_OE        : out   std_logic;
          MMUART0_TXD_USBC_DIR_MGPIO27B_OE        : out   std_logic;
          MMUART1_CTS_MGPIO13B_OE                 : out   std_logic;
          MMUART1_DCD_MGPIO16B_OE                 : out   std_logic;
          MMUART1_DSR_MGPIO14B_OE                 : out   std_logic;
          MMUART1_DTR_MGPIO12B_OE                 : out   std_logic;
          MMUART1_RI_MGPIO15B_OE                  : out   std_logic;
          MMUART1_RTS_MGPIO11B_OE                 : out   std_logic;
          MMUART1_RXD_USBC_DATA3_MGPIO26B_OE      : out   std_logic;
          MMUART1_SCK_USBC_DATA4_MGPIO25B_OE      : out   std_logic;
          MMUART1_TXD_USBC_DATA2_MGPIO24B_OE      : out   std_logic;
          RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE     : out   std_logic;
          RGMII_MDC_RMII_MDC_OE                   : out   std_logic;
          RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE      : out   std_logic;
          RGMII_RX_CLK_OE                         : out   std_logic;
          RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE  : out   std_logic;
          RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE      : out   std_logic;
          RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE      : out   std_logic;
          RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE     : out   std_logic;
          RGMII_RXD3_USBB_DATA4_OE                : out   std_logic;
          RGMII_TX_CLK_OE                         : out   std_logic;
          RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE     : out   std_logic;
          RGMII_TXD0_RMII_TXD0_USBB_DIR_OE        : out   std_logic;
          RGMII_TXD1_RMII_TXD1_USBB_STP_OE        : out   std_logic;
          RGMII_TXD2_USBB_DATA5_OE                : out   std_logic;
          RGMII_TXD3_USBB_DATA6_OE                : out   std_logic;
          SPI0_SCK_USBA_XCLK_OE                   : out   std_logic;
          SPI0_SDI_USBA_DIR_MGPIO5A_OE            : out   std_logic;
          SPI0_SDO_USBA_STP_MGPIO6A_OE            : out   std_logic;
          SPI0_SS0_USBA_NXT_MGPIO7A_OE            : out   std_logic;
          SPI0_SS1_USBA_DATA5_MGPIO8A_OE          : out   std_logic;
          SPI0_SS2_USBA_DATA6_MGPIO9A_OE          : out   std_logic;
          SPI0_SS3_USBA_DATA7_MGPIO10A_OE         : out   std_logic;
          SPI0_SS4_MGPIO19A_OE                    : out   std_logic;
          SPI0_SS5_MGPIO20A_OE                    : out   std_logic;
          SPI0_SS6_MGPIO21A_OE                    : out   std_logic;
          SPI0_SS7_MGPIO22A_OE                    : out   std_logic;
          SPI1_SCK_OE                             : out   std_logic;
          SPI1_SDI_MGPIO11A_OE                    : out   std_logic;
          SPI1_SDO_MGPIO12A_OE                    : out   std_logic;
          SPI1_SS0_MGPIO13A_OE                    : out   std_logic;
          SPI1_SS1_MGPIO14A_OE                    : out   std_logic;
          SPI1_SS2_MGPIO15A_OE                    : out   std_logic;
          SPI1_SS3_MGPIO16A_OE                    : out   std_logic;
          SPI1_SS4_MGPIO17A_OE                    : out   std_logic;
          SPI1_SS5_MGPIO18A_OE                    : out   std_logic;
          SPI1_SS6_MGPIO23A_OE                    : out   std_logic;
          SPI1_SS7_MGPIO24A_OE                    : out   std_logic;
          USBC_XCLK_OE                            : out   std_logic;
          USBD_DATA0_OE                           : out   std_logic;
          USBD_DATA1_OE                           : out   std_logic;
          USBD_DATA2_OE                           : out   std_logic;
          USBD_DATA3_OE                           : out   std_logic;
          USBD_DATA4_OE                           : out   std_logic;
          USBD_DATA5_OE                           : out   std_logic;
          USBD_DATA6_OE                           : out   std_logic;
          USBD_DATA7_MGPIO23B_OE                  : out   std_logic;
          USBD_DIR_OE                             : out   std_logic;
          USBD_NXT_OE                             : out   std_logic;
          USBD_STP_OE                             : out   std_logic;
          USBD_XCLK_OE                            : out   std_logic
        );
  end component;

  component OUTBUF_DIFF
    generic (IOSTD:string := "");

    port( D    : in    std_logic := 'U';
          PADP : out   std_logic;
          PADN : out   std_logic
        );
  end component;

    signal \CORECONFIGP_0_APB_S_PCLK\, FIC_2_APB_M_PCLK, 
        \CORECONFIGP_0_APB_S_PRESET_N\, CONFIG_PRESET_N, 
        MSS_ADLIB_INST_SPI0_SS1_USBA_DATA5_MGPIO8A_OUT, 
        MSS_ADLIB_INST_SPI0_SS1_USBA_DATA5_MGPIO8A_OE, 
        SPI_0_SS0_PAD_Y, 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT, 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE, 
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT, 
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE, 
        SPI_0_DI_PAD_Y, SPI_0_CLK_PAD_Y, 
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT, 
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE, 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT, 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE, 
        MMUART_1_RXD_PAD_Y, MSS_ADLIB_INST_DRAM_WEN, 
        MSS_ADLIB_INST_DRAM_RSTN, MSS_ADLIB_INST_DRAM_RASN, 
        MSS_ADLIB_INST_DRAM_ODT, \DRAM_FIFO_WE_OUT_net_0[0]\, 
        MDDR_DQS_TMATCH_0_IN_PAD_Y, MDDR_DQS_1_PAD_Y, 
        \DRAM_DQS_OUT_net_0[1]\, \DRAM_DQS_OE_net_0[1]\, 
        MDDR_DQS_0_PAD_Y, \DRAM_DQS_OUT_net_0[0]\, 
        \DRAM_DQS_OE_net_0[0]\, MDDR_DQ_15_PAD_Y, 
        \DRAM_DQ_OUT_net_0[15]\, \DRAM_DQ_OE_net_0[15]\, 
        MDDR_DQ_14_PAD_Y, \DRAM_DQ_OUT_net_0[14]\, 
        \DRAM_DQ_OE_net_0[14]\, MDDR_DQ_13_PAD_Y, 
        \DRAM_DQ_OUT_net_0[13]\, \DRAM_DQ_OE_net_0[13]\, 
        MDDR_DQ_12_PAD_Y, \DRAM_DQ_OUT_net_0[12]\, 
        \DRAM_DQ_OE_net_0[12]\, MDDR_DQ_11_PAD_Y, 
        \DRAM_DQ_OUT_net_0[11]\, \DRAM_DQ_OE_net_0[11]\, 
        MDDR_DQ_10_PAD_Y, \DRAM_DQ_OUT_net_0[10]\, 
        \DRAM_DQ_OE_net_0[10]\, MDDR_DQ_9_PAD_Y, 
        \DRAM_DQ_OUT_net_0[9]\, \DRAM_DQ_OE_net_0[9]\, 
        MDDR_DQ_8_PAD_Y, \DRAM_DQ_OUT_net_0[8]\, 
        \DRAM_DQ_OE_net_0[8]\, MDDR_DQ_7_PAD_Y, 
        \DRAM_DQ_OUT_net_0[7]\, \DRAM_DQ_OE_net_0[7]\, 
        MDDR_DQ_6_PAD_Y, \DRAM_DQ_OUT_net_0[6]\, 
        \DRAM_DQ_OE_net_0[6]\, MDDR_DQ_5_PAD_Y, 
        \DRAM_DQ_OUT_net_0[5]\, \DRAM_DQ_OE_net_0[5]\, 
        MDDR_DQ_4_PAD_Y, \DRAM_DQ_OUT_net_0[4]\, 
        \DRAM_DQ_OE_net_0[4]\, MDDR_DQ_3_PAD_Y, 
        \DRAM_DQ_OUT_net_0[3]\, \DRAM_DQ_OE_net_0[3]\, 
        MDDR_DQ_2_PAD_Y, \DRAM_DQ_OUT_net_0[2]\, 
        \DRAM_DQ_OE_net_0[2]\, MDDR_DQ_1_PAD_Y, 
        \DRAM_DQ_OUT_net_0[1]\, \DRAM_DQ_OE_net_0[1]\, 
        MDDR_DQ_0_PAD_Y, \DRAM_DQ_OUT_net_0[0]\, 
        \DRAM_DQ_OE_net_0[0]\, MDDR_DM_RDQS_1_PAD_Y, 
        \DRAM_DM_RDQS_OUT_net_0[1]\, \DM_OE_net_0[1]\, 
        MDDR_DM_RDQS_0_PAD_Y, \DRAM_DM_RDQS_OUT_net_0[0]\, 
        \DM_OE_net_0[0]\, MSS_ADLIB_INST_DRAM_CSN, 
        MSS_ADLIB_INST_DRAM_CKE, MSS_ADLIB_INST_DRAM_CASN, 
        \DRAM_BA_net_0[2]\, \DRAM_BA_net_0[1]\, 
        \DRAM_BA_net_0[0]\, \DRAM_ADDR_net_0[15]\, 
        \DRAM_ADDR_net_0[14]\, \DRAM_ADDR_net_0[13]\, 
        \DRAM_ADDR_net_0[12]\, \DRAM_ADDR_net_0[11]\, 
        \DRAM_ADDR_net_0[10]\, \DRAM_ADDR_net_0[9]\, 
        \DRAM_ADDR_net_0[8]\, \DRAM_ADDR_net_0[7]\, 
        \DRAM_ADDR_net_0[6]\, \DRAM_ADDR_net_0[5]\, 
        \DRAM_ADDR_net_0[4]\, \DRAM_ADDR_net_0[3]\, 
        \DRAM_ADDR_net_0[2]\, \DRAM_ADDR_net_0[1]\, 
        \DRAM_ADDR_net_0[0]\, I2C_1_SDA_PAD_Y, 
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OUT, 
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OE, 
        I2C_1_SCL_PAD_Y, 
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OUT, 
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OE, 
        GPIO_GPIO_31_BI_PAD_Y, MSS_ADLIB_INST_MGPIO31A_OUT, 
        MSS_ADLIB_INST_MGPIO31A_OE, GPIO_GPIO_26_BI_PAD_Y, 
        MSS_ADLIB_INST_MGPIO26A_OUT, MSS_ADLIB_INST_MGPIO26A_OE, 
        GPIO_GPIO_25_BI_PAD_Y, MSS_ADLIB_INST_MGPIO25A_OUT, 
        MSS_ADLIB_INST_MGPIO25A_OE, 
        MSS_ADLIB_INST_SPI0_SS5_MGPIO20A_OUT, 
        GPIO_GPIO_18_BI_PAD_Y, 
        MSS_ADLIB_INST_SPI1_SS5_MGPIO18A_OUT, 
        MSS_ADLIB_INST_SPI1_SS5_MGPIO18A_OE, 
        GPIO_GPIO_17_BI_PAD_Y, 
        MSS_ADLIB_INST_SPI1_SS4_MGPIO17A_OUT, 
        MSS_ADLIB_INST_SPI1_SS4_MGPIO17A_OE, 
        GPIO_GPIO_16_BI_PAD_Y, 
        MSS_ADLIB_INST_MMUART1_DCD_MGPIO16B_OUT, 
        MSS_ADLIB_INST_MMUART1_DCD_MGPIO16B_OE, 
        GPIO_GPIO_15_BI_PAD_Y, 
        MSS_ADLIB_INST_MMUART1_RI_MGPIO15B_OUT, 
        MSS_ADLIB_INST_MMUART1_RI_MGPIO15B_OE, 
        GPIO_GPIO_14_BI_PAD_Y, 
        MSS_ADLIB_INST_MMUART1_DSR_MGPIO14B_OUT, 
        MSS_ADLIB_INST_MMUART1_DSR_MGPIO14B_OE, 
        GPIO_GPIO_12_BI_PAD_Y, 
        MSS_ADLIB_INST_MMUART1_DTR_MGPIO12B_OUT, 
        MSS_ADLIB_INST_MMUART1_DTR_MGPIO12B_OE, 
        GPIO_GPIO_4_BI_PAD_Y, 
        MSS_ADLIB_INST_CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT, 
        MSS_ADLIB_INST_CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE, 
        GPIO_GPIO_3_BI_PAD_Y, 
        MSS_ADLIB_INST_CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT, 
        MSS_ADLIB_INST_CAN_RXBUS_USBA_DATA1_MGPIO3A_OE, 
        GPIO_GPIO_0_BI_PAD_Y, MSS_ADLIB_INST_MGPIO0B_OUT, 
        MSS_ADLIB_INST_MGPIO0B_OE, VCC_net_1, GND_net_1, 
        MSS_ADLIB_INST_DRAM_CLK : std_logic;
    signal nc228, nc203, nc216, nc194, nc151, nc23, nc175, nc58, 
        nc116, nc74, nc133, nc238, nc167, nc84, nc39, nc72, nc212, 
        nc205, nc82, nc145, nc181, nc160, nc57, nc156, nc125, 
        nc211, nc73, nc107, nc66, nc83, nc9, nc171, nc54, nc135, 
        nc41, nc100, nc52, nc186, nc29, nc118, nc60, nc141, nc193, 
        nc214, nc240, nc45, nc53, nc121, nc176, nc220, nc158, 
        nc209, nc246, nc162, nc11, nc131, nc96, nc79, nc226, 
        nc146, nc230, nc89, nc119, nc48, nc213, nc126, nc195, 
        nc188, nc242, nc15, nc236, nc102, nc3, nc207, nc47, nc90, 
        nc222, nc159, nc136, nc241, nc178, nc215, nc59, nc221, 
        nc232, nc18, nc44, nc117, nc189, nc164, nc148, nc42, 
        nc231, nc191, nc17, nc2, nc110, nc128, nc244, nc43, nc179, 
        nc157, nc36, nc224, nc61, nc104, nc138, nc14, nc150, 
        nc196, nc234, nc149, nc12, nc219, nc30, nc243, nc187, 
        nc65, nc7, nc129, nc8, nc223, nc13, nc180, nc26, nc177, 
        nc139, nc245, nc233, nc163, nc112, nc68, nc49, nc217, 
        nc170, nc91, nc225, nc5, nc20, nc198, nc147, nc67, nc152, 
        nc127, nc103, nc235, nc76, nc208, nc140, nc86, nc95, 
        nc120, nc165, nc137, nc64, nc19, nc70, nc182, nc62, nc199, 
        nc80, nc130, nc98, nc114, nc56, nc105, nc63, nc172, nc229, 
        nc97, nc161, nc31, nc154, nc50, nc239, nc142, nc94, nc197, 
        nc122, nc35, nc4, nc227, nc92, nc101, nc184, nc200, nc190, 
        nc166, nc132, nc21, nc237, nc93, nc69, nc206, nc174, nc38, 
        nc113, nc218, nc106, nc25, nc1, nc37, nc202, nc144, nc153, 
        nc46, nc71, nc124, nc81, nc201, nc168, nc34, nc28, nc115, 
        nc192, nc134, nc32, nc40, nc99, nc75, nc183, nc85, nc27, 
        nc108, nc16, nc155, nc51, nc33, nc204, nc173, nc169, nc78, 
        nc24, nc88, nc111, nc55, nc10, nc22, nc210, nc185, nc143, 
        nc77, nc6, nc109, nc87, nc123 : std_logic;

begin 

    CORECONFIGP_0_APB_S_PRESET_N <= 
        \CORECONFIGP_0_APB_S_PRESET_N\;
    CORECONFIGP_0_APB_S_PCLK <= \CORECONFIGP_0_APB_S_PCLK\;

    MDDR_ADDR_6_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[6]\, PAD => MDDR_ADDR(6));
    
    MDDR_CAS_N_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => MSS_ADLIB_INST_DRAM_CASN, PAD => MDDR_CAS_N);
    
    MDDR_RESET_N_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => MSS_ADLIB_INST_DRAM_RSTN, PAD => MDDR_RESET_N);
    
    MDDR_ODT_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => MSS_ADLIB_INST_DRAM_ODT, PAD => MDDR_ODT);
    
    GPIO_GPIO_31_BI_PAD : BIBUF
      port map(PAD => GPIO_31_BI, D => 
        MSS_ADLIB_INST_MGPIO31A_OUT, E => 
        MSS_ADLIB_INST_MGPIO31A_OE, Y => GPIO_GPIO_31_BI_PAD_Y);
    
    MDDR_ADDR_11_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[11]\, PAD => MDDR_ADDR(11));
    
    MMUART_1_TXD_PAD : TRIBUFF
      port map(D => 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT, E => 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE, PAD
         => MMUART_1_TXD);
    
    MDDR_DQ_10_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(10), D => \DRAM_DQ_OUT_net_0[10]\, 
        E => \DRAM_DQ_OE_net_0[10]\, Y => MDDR_DQ_10_PAD_Y);
    
    MDDR_DQ_1_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(1), D => \DRAM_DQ_OUT_net_0[1]\, E
         => \DRAM_DQ_OE_net_0[1]\, Y => MDDR_DQ_1_PAD_Y);
    
    MDDR_ADDR_7_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[7]\, PAD => MDDR_ADDR(7));
    
    MDDR_DQ_11_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(11), D => \DRAM_DQ_OUT_net_0[11]\, 
        E => \DRAM_DQ_OE_net_0[11]\, Y => MDDR_DQ_11_PAD_Y);
    
    MDDR_DQ_9_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(9), D => \DRAM_DQ_OUT_net_0[9]\, E
         => \DRAM_DQ_OE_net_0[9]\, Y => MDDR_DQ_9_PAD_Y);
    
    MSS_ADLIB_INST_RNI1CJ7 : CLKINT
      port map(A => CONFIG_PRESET_N, Y => 
        \CORECONFIGP_0_APB_S_PRESET_N\);
    
    MDDR_DQ_3_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(3), D => \DRAM_DQ_OUT_net_0[3]\, E
         => \DRAM_DQ_OE_net_0[3]\, Y => MDDR_DQ_3_PAD_Y);
    
    GPIO_GPIO_25_BI_PAD : BIBUF
      port map(PAD => GPIO_25_BI, D => 
        MSS_ADLIB_INST_MGPIO25A_OUT, E => 
        MSS_ADLIB_INST_MGPIO25A_OE, Y => GPIO_GPIO_25_BI_PAD_Y);
    
    MDDR_DQ_0_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(0), D => \DRAM_DQ_OUT_net_0[0]\, E
         => \DRAM_DQ_OE_net_0[0]\, Y => MDDR_DQ_0_PAD_Y);
    
    MDDR_ADDR_12_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[12]\, PAD => MDDR_ADDR(12));
    
    GPIO_GPIO_17_BI_PAD : BIBUF
      port map(PAD => GPIO_17_BI, D => 
        MSS_ADLIB_INST_SPI1_SS4_MGPIO17A_OUT, E => 
        MSS_ADLIB_INST_SPI1_SS4_MGPIO17A_OE, Y => 
        GPIO_GPIO_17_BI_PAD_Y);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    MDDR_DQ_2_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(2), D => \DRAM_DQ_OUT_net_0[2]\, E
         => \DRAM_DQ_OE_net_0[2]\, Y => MDDR_DQ_2_PAD_Y);
    
    MDDR_DQ_12_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(12), D => \DRAM_DQ_OUT_net_0[12]\, 
        E => \DRAM_DQ_OE_net_0[12]\, Y => MDDR_DQ_12_PAD_Y);
    
    MDDR_CKE_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => MSS_ADLIB_INST_DRAM_CKE, PAD => MDDR_CKE);
    
    MDDR_ADDR_2_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[2]\, PAD => MDDR_ADDR(2));
    
    GPIO_GPIO_0_BI_PAD : BIBUF
      port map(PAD => GPIO_0_BI, D => MSS_ADLIB_INST_MGPIO0B_OUT, 
        E => MSS_ADLIB_INST_MGPIO0B_OE, Y => GPIO_GPIO_0_BI_PAD_Y);
    
    FIC_2_APB_M_PCLK_inferred_clock_RNIPG5_0 : CFG1
      generic map(INIT => "01")

      port map(A => \CORECONFIGP_0_APB_S_PCLK\, Y => 
        CORECONFIGP_0_APB_S_PCLK_i);
    
    MDDR_ADDR_13_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[13]\, PAD => MDDR_ADDR(13));
    
    I2C_1_SDA_PAD : BIBUF
      port map(PAD => I2C_1_SDA, D => 
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OUT, E => 
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OE, Y => 
        I2C_1_SDA_PAD_Y);
    
    I2C_1_SCL_PAD : BIBUF
      port map(PAD => I2C_1_SCL, D => 
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OUT, E => 
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OE, Y => 
        I2C_1_SCL_PAD_Y);
    
    MDDR_ADDR_5_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[5]\, PAD => MDDR_ADDR(5));
    
    MDDR_DM_RDQS_1_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DM_RDQS(1), D => 
        \DRAM_DM_RDQS_OUT_net_0[1]\, E => \DM_OE_net_0[1]\, Y => 
        MDDR_DM_RDQS_1_PAD_Y);
    
    GPIO_GPIO_12_BI_PAD : BIBUF
      port map(PAD => GPIO_12_BI, D => 
        MSS_ADLIB_INST_MMUART1_DTR_MGPIO12B_OUT, E => 
        MSS_ADLIB_INST_MMUART1_DTR_MGPIO12B_OE, Y => 
        GPIO_GPIO_12_BI_PAD_Y);
    
    SPI_0_DO_PAD : TRIBUFF
      port map(D => MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT, 
        E => MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE, PAD => 
        SPI_0_DO);
    
    MDDR_DQS_0_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQS(0), D => \DRAM_DQS_OUT_net_0[0]\, 
        E => \DRAM_DQS_OE_net_0[0]\, Y => MDDR_DQS_0_PAD_Y);
    
    MDDR_DQS_1_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQS(1), D => \DRAM_DQS_OUT_net_0[1]\, 
        E => \DRAM_DQS_OE_net_0[1]\, Y => MDDR_DQS_1_PAD_Y);
    
    MDDR_DQ_15_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(15), D => \DRAM_DQ_OUT_net_0[15]\, 
        E => \DRAM_DQ_OE_net_0[15]\, Y => MDDR_DQ_15_PAD_Y);
    
    MDDR_DM_RDQS_0_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DM_RDQS(0), D => 
        \DRAM_DM_RDQS_OUT_net_0[0]\, E => \DM_OE_net_0[0]\, Y => 
        MDDR_DM_RDQS_0_PAD_Y);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    SPI_0_DI_PAD : INBUF
      port map(PAD => SPI_0_DI, Y => SPI_0_DI_PAD_Y);
    
    MDDR_DQ_8_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(8), D => \DRAM_DQ_OUT_net_0[8]\, E
         => \DRAM_DQ_OE_net_0[8]\, Y => MDDR_DQ_8_PAD_Y);
    
    GPIO_GPIO_14_BI_PAD : BIBUF
      port map(PAD => GPIO_14_BI, D => 
        MSS_ADLIB_INST_MMUART1_DSR_MGPIO14B_OUT, E => 
        MSS_ADLIB_INST_MMUART1_DSR_MGPIO14B_OE, Y => 
        GPIO_GPIO_14_BI_PAD_Y);
    
    GPIO_GPIO_4_BI_PAD : BIBUF
      port map(PAD => GPIO_4_BI, D => 
        MSS_ADLIB_INST_CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT, E => 
        MSS_ADLIB_INST_CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE, Y => 
        GPIO_GPIO_4_BI_PAD_Y);
    
    MDDR_ADDR_9_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[9]\, PAD => MDDR_ADDR(9));
    
    MDDR_BA_2_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_BA_net_0[2]\, PAD => MDDR_BA(2));
    
    MDDR_ADDR_14_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[14]\, PAD => MDDR_ADDR(14));
    
    MSS_ADLIB_INST : MSS_060

              generic map(INIT => "00" & x"000000000000030000000000000003610008090A4290800908000000090A42000000000C03000000009000000000200012036190A4200001004000000000000000000000000000000000000F000000000000000000000000000000007FFFFFFFB000001007C35C804248006090801041A3FFFFE400000000000846809D001F0F41C000000025A00010842108421000001FE34001FF8000000400000000020CD1007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
         ACT_UBITS => x"FFFFFFFFFFFFFF",
         MEMORYFILE => "ENVM_init.mem", RTC_MAIN_XTL_FREQ => 0.0,
         DDR_CLK_FREQ => 142.0)

      port map(CAN_RXBUS_MGPIO3A_H2F_A => OPEN, 
        CAN_RXBUS_MGPIO3A_H2F_B => OPEN, CAN_TX_EBL_MGPIO4A_H2F_A
         => OPEN, CAN_TX_EBL_MGPIO4A_H2F_B => OPEN, 
        CAN_TXBUS_MGPIO2A_H2F_A => OPEN, CAN_TXBUS_MGPIO2A_H2F_B
         => OPEN, CLK_CONFIG_APB => FIC_2_APB_M_PCLK, COMMS_INT
         => OPEN, CONFIG_PRESET_N => CONFIG_PRESET_N, 
        EDAC_ERROR(7) => nc228, EDAC_ERROR(6) => nc203, 
        EDAC_ERROR(5) => nc216, EDAC_ERROR(4) => nc194, 
        EDAC_ERROR(3) => nc151, EDAC_ERROR(2) => nc23, 
        EDAC_ERROR(1) => nc175, EDAC_ERROR(0) => nc58, 
        F_FM0_RDATA(31) => nc116, F_FM0_RDATA(30) => nc74, 
        F_FM0_RDATA(29) => nc133, F_FM0_RDATA(28) => nc238, 
        F_FM0_RDATA(27) => nc167, F_FM0_RDATA(26) => nc84, 
        F_FM0_RDATA(25) => nc39, F_FM0_RDATA(24) => nc72, 
        F_FM0_RDATA(23) => nc212, F_FM0_RDATA(22) => nc205, 
        F_FM0_RDATA(21) => nc82, F_FM0_RDATA(20) => nc145, 
        F_FM0_RDATA(19) => nc181, F_FM0_RDATA(18) => nc160, 
        F_FM0_RDATA(17) => nc57, F_FM0_RDATA(16) => nc156, 
        F_FM0_RDATA(15) => nc125, F_FM0_RDATA(14) => nc211, 
        F_FM0_RDATA(13) => nc73, F_FM0_RDATA(12) => nc107, 
        F_FM0_RDATA(11) => nc66, F_FM0_RDATA(10) => nc83, 
        F_FM0_RDATA(9) => nc9, F_FM0_RDATA(8) => nc171, 
        F_FM0_RDATA(7) => nc54, F_FM0_RDATA(6) => nc135, 
        F_FM0_RDATA(5) => nc41, F_FM0_RDATA(4) => nc100, 
        F_FM0_RDATA(3) => nc52, F_FM0_RDATA(2) => nc186, 
        F_FM0_RDATA(1) => nc29, F_FM0_RDATA(0) => nc118, 
        F_FM0_READYOUT => OPEN, F_FM0_RESP => OPEN, 
        F_HM0_ADDR(31) => nc60, F_HM0_ADDR(30) => nc141, 
        F_HM0_ADDR(29) => nc193, F_HM0_ADDR(28) => nc214, 
        F_HM0_ADDR(27) => nc240, F_HM0_ADDR(26) => nc45, 
        F_HM0_ADDR(25) => nc53, F_HM0_ADDR(24) => nc121, 
        F_HM0_ADDR(23) => nc176, F_HM0_ADDR(22) => nc220, 
        F_HM0_ADDR(21) => nc158, F_HM0_ADDR(20) => nc209, 
        F_HM0_ADDR(19) => nc246, F_HM0_ADDR(18) => nc162, 
        F_HM0_ADDR(17) => nc11, F_HM0_ADDR(16) => nc131, 
        F_HM0_ADDR(15) => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(15), 
        F_HM0_ADDR(14) => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(14), 
        F_HM0_ADDR(13) => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(13), 
        F_HM0_ADDR(12) => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(12), 
        F_HM0_ADDR(11) => nc96, F_HM0_ADDR(10) => nc79, 
        F_HM0_ADDR(9) => nc226, F_HM0_ADDR(8) => nc146, 
        F_HM0_ADDR(7) => CoreAPB3_0_APBmslave0_PADDR(7), 
        F_HM0_ADDR(6) => CoreAPB3_0_APBmslave0_PADDR(6), 
        F_HM0_ADDR(5) => CoreAPB3_0_APBmslave0_PADDR(5), 
        F_HM0_ADDR(4) => CoreAPB3_0_APBmslave0_PADDR(4), 
        F_HM0_ADDR(3) => CoreAPB3_0_APBmslave0_PADDR(3), 
        F_HM0_ADDR(2) => CoreAPB3_0_APBmslave0_PADDR(2), 
        F_HM0_ADDR(1) => CoreAPB3_0_APBmslave0_PADDR(1), 
        F_HM0_ADDR(0) => CoreAPB3_0_APBmslave0_PADDR(0), 
        F_HM0_ENABLE => CoreAPB3_0_APBmslave0_PENABLE, F_HM0_SEL
         => m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx, F_HM0_SIZE(1)
         => nc230, F_HM0_SIZE(0) => nc89, F_HM0_TRANS1 => OPEN, 
        F_HM0_WDATA(31) => nc119, F_HM0_WDATA(30) => nc48, 
        F_HM0_WDATA(29) => nc213, F_HM0_WDATA(28) => nc126, 
        F_HM0_WDATA(27) => nc195, F_HM0_WDATA(26) => nc188, 
        F_HM0_WDATA(25) => nc242, F_HM0_WDATA(24) => nc15, 
        F_HM0_WDATA(23) => nc236, F_HM0_WDATA(22) => nc102, 
        F_HM0_WDATA(21) => nc3, F_HM0_WDATA(20) => nc207, 
        F_HM0_WDATA(19) => nc47, F_HM0_WDATA(18) => nc90, 
        F_HM0_WDATA(17) => nc222, F_HM0_WDATA(16) => nc159, 
        F_HM0_WDATA(15) => nc136, F_HM0_WDATA(14) => nc241, 
        F_HM0_WDATA(13) => nc178, F_HM0_WDATA(12) => nc215, 
        F_HM0_WDATA(11) => nc59, F_HM0_WDATA(10) => nc221, 
        F_HM0_WDATA(9) => nc232, F_HM0_WDATA(8) => nc18, 
        F_HM0_WDATA(7) => CoreAPB3_0_APBmslave0_PWDATA(7), 
        F_HM0_WDATA(6) => CoreAPB3_0_APBmslave0_PWDATA(6), 
        F_HM0_WDATA(5) => CoreAPB3_0_APBmslave0_PWDATA(5), 
        F_HM0_WDATA(4) => CoreAPB3_0_APBmslave0_PWDATA(4), 
        F_HM0_WDATA(3) => CoreAPB3_0_APBmslave0_PWDATA(3), 
        F_HM0_WDATA(2) => CoreAPB3_0_APBmslave0_PWDATA(2), 
        F_HM0_WDATA(1) => CoreAPB3_0_APBmslave0_PWDATA(1), 
        F_HM0_WDATA(0) => CoreAPB3_0_APBmslave0_PWDATA(0), 
        F_HM0_WRITE => CoreAPB3_0_APBmslave0_PWRITE, FAB_CHRGVBUS
         => OPEN, FAB_DISCHRGVBUS => OPEN, FAB_DMPULLDOWN => OPEN, 
        FAB_DPPULLDOWN => OPEN, FAB_DRVVBUS => OPEN, FAB_IDPULLUP
         => OPEN, FAB_OPMODE(1) => nc44, FAB_OPMODE(0) => nc117, 
        FAB_SUSPENDM => OPEN, FAB_TERMSEL => OPEN, FAB_TXVALID
         => OPEN, FAB_VCONTROL(3) => nc189, FAB_VCONTROL(2) => 
        nc164, FAB_VCONTROL(1) => nc148, FAB_VCONTROL(0) => nc42, 
        FAB_VCONTROLLOADM => OPEN, FAB_XCVRSEL(1) => nc231, 
        FAB_XCVRSEL(0) => nc191, FAB_XDATAOUT(7) => nc17, 
        FAB_XDATAOUT(6) => nc2, FAB_XDATAOUT(5) => nc110, 
        FAB_XDATAOUT(4) => nc128, FAB_XDATAOUT(3) => nc244, 
        FAB_XDATAOUT(2) => nc43, FAB_XDATAOUT(1) => nc179, 
        FAB_XDATAOUT(0) => nc157, FACC_GLMUX_SEL => OPEN, 
        FIC32_0_MASTER(1) => nc36, FIC32_0_MASTER(0) => nc224, 
        FIC32_1_MASTER(1) => nc61, FIC32_1_MASTER(0) => nc104, 
        FPGA_RESET_N => m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        GTX_CLK => OPEN, H2F_INTERRUPT(15) => nc138, 
        H2F_INTERRUPT(14) => nc14, H2F_INTERRUPT(13) => nc150, 
        H2F_INTERRUPT(12) => nc196, H2F_INTERRUPT(11) => nc234, 
        H2F_INTERRUPT(10) => nc149, H2F_INTERRUPT(9) => nc12, 
        H2F_INTERRUPT(8) => nc219, H2F_INTERRUPT(7) => nc30, 
        H2F_INTERRUPT(6) => nc243, H2F_INTERRUPT(5) => nc187, 
        H2F_INTERRUPT(4) => nc65, H2F_INTERRUPT(3) => nc7, 
        H2F_INTERRUPT(2) => nc129, H2F_INTERRUPT(1) => nc8, 
        H2F_INTERRUPT(0) => nc223, H2F_NMI => OPEN, H2FCALIB => 
        OPEN, I2C0_SCL_MGPIO31B_H2F_A => OPEN, 
        I2C0_SCL_MGPIO31B_H2F_B => OPEN, I2C0_SDA_MGPIO30B_H2F_A
         => OPEN, I2C0_SDA_MGPIO30B_H2F_B => OPEN, 
        I2C1_SCL_MGPIO1A_H2F_A => 
        m2s010_som_sb_MSS_0_GPIO_1_M2F_OE, I2C1_SCL_MGPIO1A_H2F_B
         => GPIO_1_M2F, I2C1_SDA_MGPIO0A_H2F_A => OPEN, 
        I2C1_SDA_MGPIO0A_H2F_B => OPEN, MDCF => MAC_MII_MDC_c, 
        MDOENF => m2s010_som_sb_MSS_0_MAC_MII_MDO_EN, MDOF => 
        m2s010_som_sb_MSS_0_MAC_MII_MDO, 
        MMUART0_CTS_MGPIO19B_H2F_A => OPEN, 
        MMUART0_CTS_MGPIO19B_H2F_B => OPEN, 
        MMUART0_DCD_MGPIO22B_H2F_A => OPEN, 
        MMUART0_DCD_MGPIO22B_H2F_B => GPIO_22_M2F_c, 
        MMUART0_DSR_MGPIO20B_H2F_A => OPEN, 
        MMUART0_DSR_MGPIO20B_H2F_B => OPEN, 
        MMUART0_DTR_MGPIO18B_H2F_A => OPEN, 
        MMUART0_DTR_MGPIO18B_H2F_B => OPEN, 
        MMUART0_RI_MGPIO21B_H2F_A => OPEN, 
        MMUART0_RI_MGPIO21B_H2F_B => GPIO_21_M2F_c, 
        MMUART0_RTS_MGPIO17B_H2F_A => OPEN, 
        MMUART0_RTS_MGPIO17B_H2F_B => OPEN, 
        MMUART0_RXD_MGPIO28B_H2F_A => OPEN, 
        MMUART0_RXD_MGPIO28B_H2F_B => 
        m2s010_som_sb_0_GPIO_28_SW_RESET, 
        MMUART0_SCK_MGPIO29B_H2F_A => OPEN, 
        MMUART0_SCK_MGPIO29B_H2F_B => OPEN, 
        MMUART0_TXD_MGPIO27B_H2F_A => MMUART_0_TXD_M2F_c, 
        MMUART0_TXD_MGPIO27B_H2F_B => OPEN, 
        MMUART1_DTR_MGPIO12B_H2F_A => OPEN, 
        MMUART1_RTS_MGPIO11B_H2F_A => OPEN, 
        MMUART1_RTS_MGPIO11B_H2F_B => OPEN, 
        MMUART1_RXD_MGPIO26B_H2F_A => OPEN, 
        MMUART1_RXD_MGPIO26B_H2F_B => OPEN, 
        MMUART1_SCK_MGPIO25B_H2F_A => OPEN, 
        MMUART1_SCK_MGPIO25B_H2F_B => OPEN, 
        MMUART1_TXD_MGPIO24B_H2F_A => OPEN, 
        MMUART1_TXD_MGPIO24B_H2F_B => GPIO_24_M2F_c, MPLL_LOCK
         => OPEN, PER2_FABRIC_PADDR(15) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(15), 
        PER2_FABRIC_PADDR(14) => nc13, PER2_FABRIC_PADDR(13) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(13), 
        PER2_FABRIC_PADDR(12) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(12), 
        PER2_FABRIC_PADDR(11) => nc180, PER2_FABRIC_PADDR(10) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(10), 
        PER2_FABRIC_PADDR(9) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(9), 
        PER2_FABRIC_PADDR(8) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(8), 
        PER2_FABRIC_PADDR(7) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(7), 
        PER2_FABRIC_PADDR(6) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(6), 
        PER2_FABRIC_PADDR(5) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(5), 
        PER2_FABRIC_PADDR(4) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), 
        PER2_FABRIC_PADDR(3) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), 
        PER2_FABRIC_PADDR(2) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), 
        PER2_FABRIC_PENABLE => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE, 
        PER2_FABRIC_PSEL => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx, 
        PER2_FABRIC_PWDATA(31) => nc26, PER2_FABRIC_PWDATA(30)
         => nc177, PER2_FABRIC_PWDATA(29) => nc139, 
        PER2_FABRIC_PWDATA(28) => nc245, PER2_FABRIC_PWDATA(27)
         => nc233, PER2_FABRIC_PWDATA(26) => nc163, 
        PER2_FABRIC_PWDATA(25) => nc112, PER2_FABRIC_PWDATA(24)
         => nc68, PER2_FABRIC_PWDATA(23) => nc49, 
        PER2_FABRIC_PWDATA(22) => nc217, PER2_FABRIC_PWDATA(21)
         => nc170, PER2_FABRIC_PWDATA(20) => nc91, 
        PER2_FABRIC_PWDATA(19) => nc225, PER2_FABRIC_PWDATA(18)
         => nc5, PER2_FABRIC_PWDATA(17) => nc20, 
        PER2_FABRIC_PWDATA(16) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(16), 
        PER2_FABRIC_PWDATA(15) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(15), 
        PER2_FABRIC_PWDATA(14) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(14), 
        PER2_FABRIC_PWDATA(13) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(13), 
        PER2_FABRIC_PWDATA(12) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(12), 
        PER2_FABRIC_PWDATA(11) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(11), 
        PER2_FABRIC_PWDATA(10) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(10), 
        PER2_FABRIC_PWDATA(9) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(9), 
        PER2_FABRIC_PWDATA(8) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(8), 
        PER2_FABRIC_PWDATA(7) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(7), 
        PER2_FABRIC_PWDATA(6) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(6), 
        PER2_FABRIC_PWDATA(5) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(5), 
        PER2_FABRIC_PWDATA(4) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(4), 
        PER2_FABRIC_PWDATA(3) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(3), 
        PER2_FABRIC_PWDATA(2) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(2), 
        PER2_FABRIC_PWDATA(1) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(1), 
        PER2_FABRIC_PWDATA(0) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(0), 
        PER2_FABRIC_PWRITE => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE, 
        RTC_MATCH => OPEN, SLEEPDEEP => OPEN, SLEEPHOLDACK => 
        OPEN, SLEEPING => OPEN, SMBALERT_NO0 => OPEN, 
        SMBALERT_NO1 => OPEN, SMBSUS_NO0 => OPEN, SMBSUS_NO1 => 
        OPEN, SPI0_CLK_OUT => OPEN, SPI0_SDI_MGPIO5A_H2F_A => 
        OPEN, SPI0_SDI_MGPIO5A_H2F_B => GPIO_5_M2F_c, 
        SPI0_SDO_MGPIO6A_H2F_A => 
        m2s010_som_sb_MSS_0_GPIO_6_M2F_OE, SPI0_SDO_MGPIO6A_H2F_B
         => m2s010_som_sb_MSS_0_GPIO_6_M2F, 
        SPI0_SS0_MGPIO7A_H2F_A => 
        m2s010_som_sb_MSS_0_GPIO_7_M2F_OE, SPI0_SS0_MGPIO7A_H2F_B
         => m2s010_som_sb_MSS_0_GPIO_7_M2F, 
        SPI0_SS1_MGPIO8A_H2F_A => OPEN, SPI0_SS1_MGPIO8A_H2F_B
         => GPIO_8_M2F_c, SPI0_SS2_MGPIO9A_H2F_A => OPEN, 
        SPI0_SS2_MGPIO9A_H2F_B => OPEN, SPI0_SS3_MGPIO10A_H2F_A
         => OPEN, SPI0_SS3_MGPIO10A_H2F_B => OPEN, 
        SPI0_SS4_MGPIO19A_H2F_A => OPEN, SPI0_SS5_MGPIO20A_H2F_A
         => OPEN, SPI0_SS6_MGPIO21A_H2F_A => OPEN, 
        SPI0_SS7_MGPIO22A_H2F_A => OPEN, SPI1_CLK_OUT => 
        m2s010_som_sb_MSS_0_SPI_1_CLK_M2F, 
        SPI1_SDI_MGPIO11A_H2F_A => OPEN, SPI1_SDI_MGPIO11A_H2F_B
         => GPIO_11_M2F_c, SPI1_SDO_MGPIO12A_H2F_A => 
        SPI_1_DO_CAM_c, SPI1_SDO_MGPIO12A_H2F_B => OPEN, 
        SPI1_SS0_MGPIO13A_H2F_A => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F, 
        SPI1_SS0_MGPIO13A_H2F_B => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE, 
        SPI1_SS1_MGPIO14A_H2F_A => OPEN, SPI1_SS1_MGPIO14A_H2F_B
         => OPEN, SPI1_SS2_MGPIO15A_H2F_A => OPEN, 
        SPI1_SS2_MGPIO15A_H2F_B => OPEN, SPI1_SS3_MGPIO16A_H2F_A
         => OPEN, SPI1_SS3_MGPIO16A_H2F_B => OPEN, 
        SPI1_SS4_MGPIO17A_H2F_A => OPEN, SPI1_SS5_MGPIO18A_H2F_A
         => OPEN, SPI1_SS6_MGPIO23A_H2F_A => OPEN, 
        SPI1_SS7_MGPIO24A_H2F_A => OPEN, TCGF(9) => nc198, 
        TCGF(8) => nc147, TCGF(7) => nc67, TCGF(6) => nc152, 
        TCGF(5) => nc127, TCGF(4) => nc103, TCGF(3) => nc235, 
        TCGF(2) => nc76, TCGF(1) => nc208, TCGF(0) => nc140, 
        TRACECLK => OPEN, TRACEDATA(3) => nc86, TRACEDATA(2) => 
        nc95, TRACEDATA(1) => nc120, TRACEDATA(0) => nc165, 
        TX_CLK => OPEN, TX_ENF => MAC_MII_TX_EN_c, TX_ERRF => 
        OPEN, TXCTL_EN_RIF => OPEN, TXD_RIF(3) => nc137, 
        TXD_RIF(2) => nc64, TXD_RIF(1) => nc19, TXD_RIF(0) => 
        nc70, TXDF(7) => nc182, TXDF(6) => nc62, TXDF(5) => nc199, 
        TXDF(4) => nc80, TXDF(3) => MAC_MII_TXD_c(3), TXDF(2) => 
        MAC_MII_TXD_c(2), TXDF(1) => MAC_MII_TXD_c(1), TXDF(0)
         => MAC_MII_TXD_c(0), TXEV => OPEN, WDOGTIMEOUT => OPEN, 
        F_ARREADY_HREADYOUT1 => OPEN, F_AWREADY_HREADYOUT0 => 
        OPEN, F_BID(3) => nc130, F_BID(2) => nc98, F_BID(1) => 
        nc114, F_BID(0) => nc56, F_BRESP_HRESP0(1) => nc105, 
        F_BRESP_HRESP0(0) => nc63, F_BVALID => OPEN, 
        F_RDATA_HRDATA01(63) => nc172, F_RDATA_HRDATA01(62) => 
        nc229, F_RDATA_HRDATA01(61) => nc97, F_RDATA_HRDATA01(60)
         => nc161, F_RDATA_HRDATA01(59) => nc31, 
        F_RDATA_HRDATA01(58) => nc154, F_RDATA_HRDATA01(57) => 
        nc50, F_RDATA_HRDATA01(56) => nc239, F_RDATA_HRDATA01(55)
         => nc142, F_RDATA_HRDATA01(54) => nc94, 
        F_RDATA_HRDATA01(53) => nc197, F_RDATA_HRDATA01(52) => 
        nc122, F_RDATA_HRDATA01(51) => nc35, F_RDATA_HRDATA01(50)
         => nc4, F_RDATA_HRDATA01(49) => nc227, 
        F_RDATA_HRDATA01(48) => nc92, F_RDATA_HRDATA01(47) => 
        nc101, F_RDATA_HRDATA01(46) => nc184, 
        F_RDATA_HRDATA01(45) => nc200, F_RDATA_HRDATA01(44) => 
        nc190, F_RDATA_HRDATA01(43) => nc166, 
        F_RDATA_HRDATA01(42) => nc132, F_RDATA_HRDATA01(41) => 
        nc21, F_RDATA_HRDATA01(40) => nc237, F_RDATA_HRDATA01(39)
         => nc93, F_RDATA_HRDATA01(38) => nc69, 
        F_RDATA_HRDATA01(37) => nc206, F_RDATA_HRDATA01(36) => 
        nc174, F_RDATA_HRDATA01(35) => nc38, F_RDATA_HRDATA01(34)
         => nc113, F_RDATA_HRDATA01(33) => nc218, 
        F_RDATA_HRDATA01(32) => nc106, F_RDATA_HRDATA01(31) => 
        nc25, F_RDATA_HRDATA01(30) => nc1, F_RDATA_HRDATA01(29)
         => nc37, F_RDATA_HRDATA01(28) => nc202, 
        F_RDATA_HRDATA01(27) => nc144, F_RDATA_HRDATA01(26) => 
        nc153, F_RDATA_HRDATA01(25) => nc46, F_RDATA_HRDATA01(24)
         => nc71, F_RDATA_HRDATA01(23) => nc124, 
        F_RDATA_HRDATA01(22) => nc81, F_RDATA_HRDATA01(21) => 
        nc201, F_RDATA_HRDATA01(20) => nc168, 
        F_RDATA_HRDATA01(19) => nc34, F_RDATA_HRDATA01(18) => 
        nc28, F_RDATA_HRDATA01(17) => nc115, F_RDATA_HRDATA01(16)
         => nc192, F_RDATA_HRDATA01(15) => nc134, 
        F_RDATA_HRDATA01(14) => nc32, F_RDATA_HRDATA01(13) => 
        nc40, F_RDATA_HRDATA01(12) => nc99, F_RDATA_HRDATA01(11)
         => nc75, F_RDATA_HRDATA01(10) => nc183, 
        F_RDATA_HRDATA01(9) => nc85, F_RDATA_HRDATA01(8) => nc27, 
        F_RDATA_HRDATA01(7) => nc108, F_RDATA_HRDATA01(6) => nc16, 
        F_RDATA_HRDATA01(5) => nc155, F_RDATA_HRDATA01(4) => nc51, 
        F_RDATA_HRDATA01(3) => nc33, F_RDATA_HRDATA01(2) => nc204, 
        F_RDATA_HRDATA01(1) => nc173, F_RDATA_HRDATA01(0) => 
        nc169, F_RID(3) => nc78, F_RID(2) => nc24, F_RID(1) => 
        nc88, F_RID(0) => nc111, F_RLAST => OPEN, 
        F_RRESP_HRESP1(1) => nc55, F_RRESP_HRESP1(0) => nc10, 
        F_RVALID => OPEN, F_WREADY => OPEN, 
        MDDR_FABRIC_PRDATA(15) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(15), 
        MDDR_FABRIC_PRDATA(14) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(14), 
        MDDR_FABRIC_PRDATA(13) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(13), 
        MDDR_FABRIC_PRDATA(12) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(12), 
        MDDR_FABRIC_PRDATA(11) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(11), 
        MDDR_FABRIC_PRDATA(10) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(10), 
        MDDR_FABRIC_PRDATA(9) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(9), 
        MDDR_FABRIC_PRDATA(8) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(8), 
        MDDR_FABRIC_PRDATA(7) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(7), 
        MDDR_FABRIC_PRDATA(6) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(6), 
        MDDR_FABRIC_PRDATA(5) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(5), 
        MDDR_FABRIC_PRDATA(4) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(4), 
        MDDR_FABRIC_PRDATA(3) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(3), 
        MDDR_FABRIC_PRDATA(2) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(2), 
        MDDR_FABRIC_PRDATA(1) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(1), 
        MDDR_FABRIC_PRDATA(0) => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(0), 
        MDDR_FABRIC_PREADY => CORECONFIGP_0_MDDR_APBmslave_PREADY, 
        MDDR_FABRIC_PSLVERR => 
        CORECONFIGP_0_MDDR_APBmslave_PSLVERR, CAN_RXBUS_F2H_SCP
         => VCC_net_1, CAN_TX_EBL_F2H_SCP => VCC_net_1, 
        CAN_TXBUS_F2H_SCP => VCC_net_1, COLF => MAC_MII_COL_c, 
        CRSF => MAC_MII_CRS_c, F2_DMAREADY(1) => VCC_net_1, 
        F2_DMAREADY(0) => VCC_net_1, F2H_INTERRUPT(15) => 
        GND_net_1, F2H_INTERRUPT(14) => GND_net_1, 
        F2H_INTERRUPT(13) => GND_net_1, F2H_INTERRUPT(12) => 
        GND_net_1, F2H_INTERRUPT(11) => GND_net_1, 
        F2H_INTERRUPT(10) => GND_net_1, F2H_INTERRUPT(9) => 
        GND_net_1, F2H_INTERRUPT(8) => GND_net_1, 
        F2H_INTERRUPT(7) => GND_net_1, F2H_INTERRUPT(6) => 
        GND_net_1, F2H_INTERRUPT(5) => GND_net_1, 
        F2H_INTERRUPT(4) => GND_net_1, F2H_INTERRUPT(3) => 
        GND_net_1, F2H_INTERRUPT(2) => GND_net_1, 
        F2H_INTERRUPT(1) => GND_net_1, F2H_INTERRUPT(0) => 
        CommsFPGA_top_0_INT, F2HCALIB => VCC_net_1, F_DMAREADY(1)
         => VCC_net_1, F_DMAREADY(0) => VCC_net_1, F_FM0_ADDR(31)
         => GND_net_1, F_FM0_ADDR(30) => GND_net_1, 
        F_FM0_ADDR(29) => GND_net_1, F_FM0_ADDR(28) => GND_net_1, 
        F_FM0_ADDR(27) => GND_net_1, F_FM0_ADDR(26) => GND_net_1, 
        F_FM0_ADDR(25) => GND_net_1, F_FM0_ADDR(24) => GND_net_1, 
        F_FM0_ADDR(23) => GND_net_1, F_FM0_ADDR(22) => GND_net_1, 
        F_FM0_ADDR(21) => GND_net_1, F_FM0_ADDR(20) => GND_net_1, 
        F_FM0_ADDR(19) => GND_net_1, F_FM0_ADDR(18) => GND_net_1, 
        F_FM0_ADDR(17) => GND_net_1, F_FM0_ADDR(16) => GND_net_1, 
        F_FM0_ADDR(15) => GND_net_1, F_FM0_ADDR(14) => GND_net_1, 
        F_FM0_ADDR(13) => GND_net_1, F_FM0_ADDR(12) => GND_net_1, 
        F_FM0_ADDR(11) => GND_net_1, F_FM0_ADDR(10) => GND_net_1, 
        F_FM0_ADDR(9) => GND_net_1, F_FM0_ADDR(8) => GND_net_1, 
        F_FM0_ADDR(7) => GND_net_1, F_FM0_ADDR(6) => GND_net_1, 
        F_FM0_ADDR(5) => GND_net_1, F_FM0_ADDR(4) => GND_net_1, 
        F_FM0_ADDR(3) => GND_net_1, F_FM0_ADDR(2) => GND_net_1, 
        F_FM0_ADDR(1) => GND_net_1, F_FM0_ADDR(0) => GND_net_1, 
        F_FM0_ENABLE => GND_net_1, F_FM0_MASTLOCK => GND_net_1, 
        F_FM0_READY => VCC_net_1, F_FM0_SEL => GND_net_1, 
        F_FM0_SIZE(1) => GND_net_1, F_FM0_SIZE(0) => GND_net_1, 
        F_FM0_TRANS1 => GND_net_1, F_FM0_WDATA(31) => GND_net_1, 
        F_FM0_WDATA(30) => GND_net_1, F_FM0_WDATA(29) => 
        GND_net_1, F_FM0_WDATA(28) => GND_net_1, F_FM0_WDATA(27)
         => GND_net_1, F_FM0_WDATA(26) => GND_net_1, 
        F_FM0_WDATA(25) => GND_net_1, F_FM0_WDATA(24) => 
        GND_net_1, F_FM0_WDATA(23) => GND_net_1, F_FM0_WDATA(22)
         => GND_net_1, F_FM0_WDATA(21) => GND_net_1, 
        F_FM0_WDATA(20) => GND_net_1, F_FM0_WDATA(19) => 
        GND_net_1, F_FM0_WDATA(18) => GND_net_1, F_FM0_WDATA(17)
         => GND_net_1, F_FM0_WDATA(16) => GND_net_1, 
        F_FM0_WDATA(15) => GND_net_1, F_FM0_WDATA(14) => 
        GND_net_1, F_FM0_WDATA(13) => GND_net_1, F_FM0_WDATA(12)
         => GND_net_1, F_FM0_WDATA(11) => GND_net_1, 
        F_FM0_WDATA(10) => GND_net_1, F_FM0_WDATA(9) => GND_net_1, 
        F_FM0_WDATA(8) => GND_net_1, F_FM0_WDATA(7) => GND_net_1, 
        F_FM0_WDATA(6) => GND_net_1, F_FM0_WDATA(5) => GND_net_1, 
        F_FM0_WDATA(4) => GND_net_1, F_FM0_WDATA(3) => GND_net_1, 
        F_FM0_WDATA(2) => GND_net_1, F_FM0_WDATA(1) => GND_net_1, 
        F_FM0_WDATA(0) => GND_net_1, F_FM0_WRITE => GND_net_1, 
        F_HM0_RDATA(31) => GND_net_1, F_HM0_RDATA(30) => 
        GND_net_1, F_HM0_RDATA(29) => GND_net_1, F_HM0_RDATA(28)
         => GND_net_1, F_HM0_RDATA(27) => GND_net_1, 
        F_HM0_RDATA(26) => GND_net_1, F_HM0_RDATA(25) => 
        GND_net_1, F_HM0_RDATA(24) => GND_net_1, F_HM0_RDATA(23)
         => GND_net_1, F_HM0_RDATA(22) => GND_net_1, 
        F_HM0_RDATA(21) => GND_net_1, F_HM0_RDATA(20) => 
        GND_net_1, F_HM0_RDATA(19) => GND_net_1, F_HM0_RDATA(18)
         => GND_net_1, F_HM0_RDATA(17) => GND_net_1, 
        F_HM0_RDATA(16) => GND_net_1, F_HM0_RDATA(15) => 
        GND_net_1, F_HM0_RDATA(14) => GND_net_1, F_HM0_RDATA(13)
         => GND_net_1, F_HM0_RDATA(12) => GND_net_1, 
        F_HM0_RDATA(11) => GND_net_1, F_HM0_RDATA(10) => 
        GND_net_1, F_HM0_RDATA(9) => GND_net_1, F_HM0_RDATA(8)
         => GND_net_1, F_HM0_RDATA(7) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(7), F_HM0_RDATA(6) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(6), F_HM0_RDATA(5) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(5), F_HM0_RDATA(4) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(4), F_HM0_RDATA(3) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(3), F_HM0_RDATA(2) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(2), F_HM0_RDATA(1) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(1), F_HM0_RDATA(0) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(0), F_HM0_READY => 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i, F_HM0_RESP => 
        GND_net_1, FAB_AVALID => VCC_net_1, FAB_HOSTDISCON => 
        VCC_net_1, FAB_IDDIG => VCC_net_1, FAB_LINESTATE(1) => 
        VCC_net_1, FAB_LINESTATE(0) => VCC_net_1, FAB_M3_RESET_N
         => VCC_net_1, FAB_PLL_LOCK => FAB_CCC_LOCK, FAB_RXACTIVE
         => VCC_net_1, FAB_RXERROR => VCC_net_1, FAB_RXVALID => 
        VCC_net_1, FAB_RXVALIDH => GND_net_1, FAB_SESSEND => 
        VCC_net_1, FAB_TXREADY => VCC_net_1, FAB_VBUSVALID => 
        VCC_net_1, FAB_VSTATUS(7) => VCC_net_1, FAB_VSTATUS(6)
         => VCC_net_1, FAB_VSTATUS(5) => VCC_net_1, 
        FAB_VSTATUS(4) => VCC_net_1, FAB_VSTATUS(3) => VCC_net_1, 
        FAB_VSTATUS(2) => VCC_net_1, FAB_VSTATUS(1) => VCC_net_1, 
        FAB_VSTATUS(0) => VCC_net_1, FAB_XDATAIN(7) => VCC_net_1, 
        FAB_XDATAIN(6) => VCC_net_1, FAB_XDATAIN(5) => VCC_net_1, 
        FAB_XDATAIN(4) => VCC_net_1, FAB_XDATAIN(3) => VCC_net_1, 
        FAB_XDATAIN(2) => VCC_net_1, FAB_XDATAIN(1) => VCC_net_1, 
        FAB_XDATAIN(0) => VCC_net_1, GTX_CLKPF => VCC_net_1, 
        I2C0_BCLK => VCC_net_1, I2C0_SCL_F2H_SCP => VCC_net_1, 
        I2C0_SDA_F2H_SCP => VCC_net_1, I2C1_BCLK => VCC_net_1, 
        I2C1_SCL_F2H_SCP => VCC_net_1, I2C1_SDA_F2H_SCP => 
        VCC_net_1, MDIF => BIBUF_0_Y, MGPIO0A_F2H_GPIN => 
        VCC_net_1, MGPIO10A_F2H_GPIN => Y_net_0(3), 
        MGPIO11A_F2H_GPIN => VCC_net_1, MGPIO11B_F2H_GPIN => 
        VCC_net_1, MGPIO12A_F2H_GPIN => VCC_net_1, 
        MGPIO13A_F2H_GPIN => VCC_net_1, MGPIO14A_F2H_GPIN => 
        VCC_net_1, MGPIO15A_F2H_GPIN => VCC_net_1, 
        MGPIO16A_F2H_GPIN => VCC_net_1, MGPIO17B_F2H_GPIN => 
        VCC_net_1, MGPIO18B_F2H_GPIN => VCC_net_1, 
        MGPIO19B_F2H_GPIN => Y_net_0(1), MGPIO1A_F2H_GPIN => 
        GPIO_1_in_0, MGPIO20B_F2H_GPIN => VCC_net_1, 
        MGPIO21B_F2H_GPIN => VCC_net_1, MGPIO22B_F2H_GPIN => 
        VCC_net_1, MGPIO24B_F2H_GPIN => VCC_net_1, 
        MGPIO25B_F2H_GPIN => VCC_net_1, MGPIO26B_F2H_GPIN => 
        VCC_net_1, MGPIO27B_F2H_GPIN => DEBOUNCE_OUT_1_c, 
        MGPIO28B_F2H_GPIN => VCC_net_1, MGPIO29B_F2H_GPIN => 
        DEBOUNCE_OUT_2_c, MGPIO2A_F2H_GPIN => Y_net_0(2), 
        MGPIO30B_F2H_GPIN => DEBOUNCE_OUT_net_0_0, 
        MGPIO31B_F2H_GPIN => VCC_net_1, MGPIO3A_F2H_GPIN => 
        VCC_net_1, MGPIO4A_F2H_GPIN => VCC_net_1, 
        MGPIO5A_F2H_GPIN => VCC_net_1, MGPIO6A_F2H_GPIN => 
        GPIO_6_Y_0, MGPIO7A_F2H_GPIN => GPIO_7_Y_0, 
        MGPIO8A_F2H_GPIN => VCC_net_1, MGPIO9A_F2H_GPIN => 
        Y_net_0(0), MMUART0_CTS_F2H_SCP => VCC_net_1, 
        MMUART0_DCD_F2H_SCP => VCC_net_1, MMUART0_DSR_F2H_SCP => 
        VCC_net_1, MMUART0_DTR_F2H_SCP => VCC_net_1, 
        MMUART0_RI_F2H_SCP => VCC_net_1, MMUART0_RTS_F2H_SCP => 
        VCC_net_1, MMUART0_RXD_F2H_SCP => MMUART_0_RXD_F2M_c, 
        MMUART0_SCK_F2H_SCP => VCC_net_1, MMUART0_TXD_F2H_SCP => 
        VCC_net_1, MMUART1_CTS_F2H_SCP => VCC_net_1, 
        MMUART1_DCD_F2H_SCP => VCC_net_1, MMUART1_DSR_F2H_SCP => 
        VCC_net_1, MMUART1_RI_F2H_SCP => VCC_net_1, 
        MMUART1_RTS_F2H_SCP => VCC_net_1, MMUART1_RXD_F2H_SCP => 
        VCC_net_1, MMUART1_SCK_F2H_SCP => VCC_net_1, 
        MMUART1_TXD_F2H_SCP => VCC_net_1, PER2_FABRIC_PRDATA(31)
         => GND_net_1, PER2_FABRIC_PRDATA(30) => GND_net_1, 
        PER2_FABRIC_PRDATA(29) => GND_net_1, 
        PER2_FABRIC_PRDATA(28) => GND_net_1, 
        PER2_FABRIC_PRDATA(27) => GND_net_1, 
        PER2_FABRIC_PRDATA(26) => GND_net_1, 
        PER2_FABRIC_PRDATA(25) => GND_net_1, 
        PER2_FABRIC_PRDATA(24) => GND_net_1, 
        PER2_FABRIC_PRDATA(23) => GND_net_1, 
        PER2_FABRIC_PRDATA(22) => GND_net_1, 
        PER2_FABRIC_PRDATA(21) => GND_net_1, 
        PER2_FABRIC_PRDATA(20) => GND_net_1, 
        PER2_FABRIC_PRDATA(19) => GND_net_1, 
        PER2_FABRIC_PRDATA(18) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(17), 
        PER2_FABRIC_PRDATA(17) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(17), 
        PER2_FABRIC_PRDATA(16) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(16), 
        PER2_FABRIC_PRDATA(15) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(15), 
        PER2_FABRIC_PRDATA(14) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(14), 
        PER2_FABRIC_PRDATA(13) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(13), 
        PER2_FABRIC_PRDATA(12) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(12), 
        PER2_FABRIC_PRDATA(11) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(11), 
        PER2_FABRIC_PRDATA(10) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(10), 
        PER2_FABRIC_PRDATA(9) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(9), 
        PER2_FABRIC_PRDATA(8) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(8), 
        PER2_FABRIC_PRDATA(7) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(7), 
        PER2_FABRIC_PRDATA(6) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(6), 
        PER2_FABRIC_PRDATA(5) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(5), 
        PER2_FABRIC_PRDATA(4) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(4), 
        PER2_FABRIC_PRDATA(3) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(3), 
        PER2_FABRIC_PRDATA(2) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(2), 
        PER2_FABRIC_PRDATA(1) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(1), 
        PER2_FABRIC_PRDATA(0) => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(0), 
        PER2_FABRIC_PREADY => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY, 
        PER2_FABRIC_PSLVERR => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR, RCGF(9)
         => VCC_net_1, RCGF(8) => VCC_net_1, RCGF(7) => VCC_net_1, 
        RCGF(6) => VCC_net_1, RCGF(5) => VCC_net_1, RCGF(4) => 
        VCC_net_1, RCGF(3) => VCC_net_1, RCGF(2) => VCC_net_1, 
        RCGF(1) => VCC_net_1, RCGF(0) => VCC_net_1, RX_CLKPF => 
        MAC_MII_RX_CLK_c, RX_DVF => MAC_MII_RX_DV_c, RX_ERRF => 
        MAC_MII_RX_ER_c, RX_EV => VCC_net_1, RXDF(7) => VCC_net_1, 
        RXDF(6) => VCC_net_1, RXDF(5) => VCC_net_1, RXDF(4) => 
        VCC_net_1, RXDF(3) => MAC_MII_RXD_c(3), RXDF(2) => 
        MAC_MII_RXD_c(2), RXDF(1) => MAC_MII_RXD_c(1), RXDF(0)
         => MAC_MII_RXD_c(0), SLEEPHOLDREQ => GND_net_1, 
        SMBALERT_NI0 => VCC_net_1, SMBALERT_NI1 => VCC_net_1, 
        SMBSUS_NI0 => VCC_net_1, SMBSUS_NI1 => VCC_net_1, 
        SPI0_CLK_IN => VCC_net_1, SPI0_SDI_F2H_SCP => VCC_net_1, 
        SPI0_SDO_F2H_SCP => VCC_net_1, SPI0_SS0_F2H_SCP => 
        VCC_net_1, SPI0_SS1_F2H_SCP => VCC_net_1, 
        SPI0_SS2_F2H_SCP => VCC_net_1, SPI0_SS3_F2H_SCP => 
        VCC_net_1, SPI1_CLK_IN => CAM_SPI_1_CLK_Y_0, 
        SPI1_SDI_F2H_SCP => SPI_1_DI, SPI1_SDO_F2H_SCP => 
        VCC_net_1, SPI1_SS0_F2H_SCP => SPI_1_SS0_MX_Y, 
        SPI1_SS1_F2H_SCP => VCC_net_1, SPI1_SS2_F2H_SCP => 
        VCC_net_1, SPI1_SS3_F2H_SCP => VCC_net_1, TX_CLKPF => 
        MAC_MII_TX_CLK_c, USER_MSS_GPIO_RESET_N => VCC_net_1, 
        USER_MSS_RESET_N => VCC_net_1, XCLK_FAB => VCC_net_1, 
        CLK_BASE => m2s010_som_sb_0_CCC_71MHz, CLK_MDDR_APB => 
        \CORECONFIGP_0_APB_S_PCLK\, F_ARADDR_HADDR1(31) => 
        VCC_net_1, F_ARADDR_HADDR1(30) => VCC_net_1, 
        F_ARADDR_HADDR1(29) => VCC_net_1, F_ARADDR_HADDR1(28) => 
        VCC_net_1, F_ARADDR_HADDR1(27) => VCC_net_1, 
        F_ARADDR_HADDR1(26) => VCC_net_1, F_ARADDR_HADDR1(25) => 
        VCC_net_1, F_ARADDR_HADDR1(24) => VCC_net_1, 
        F_ARADDR_HADDR1(23) => VCC_net_1, F_ARADDR_HADDR1(22) => 
        VCC_net_1, F_ARADDR_HADDR1(21) => VCC_net_1, 
        F_ARADDR_HADDR1(20) => VCC_net_1, F_ARADDR_HADDR1(19) => 
        VCC_net_1, F_ARADDR_HADDR1(18) => VCC_net_1, 
        F_ARADDR_HADDR1(17) => VCC_net_1, F_ARADDR_HADDR1(16) => 
        VCC_net_1, F_ARADDR_HADDR1(15) => VCC_net_1, 
        F_ARADDR_HADDR1(14) => VCC_net_1, F_ARADDR_HADDR1(13) => 
        VCC_net_1, F_ARADDR_HADDR1(12) => VCC_net_1, 
        F_ARADDR_HADDR1(11) => VCC_net_1, F_ARADDR_HADDR1(10) => 
        VCC_net_1, F_ARADDR_HADDR1(9) => VCC_net_1, 
        F_ARADDR_HADDR1(8) => VCC_net_1, F_ARADDR_HADDR1(7) => 
        VCC_net_1, F_ARADDR_HADDR1(6) => VCC_net_1, 
        F_ARADDR_HADDR1(5) => VCC_net_1, F_ARADDR_HADDR1(4) => 
        VCC_net_1, F_ARADDR_HADDR1(3) => VCC_net_1, 
        F_ARADDR_HADDR1(2) => VCC_net_1, F_ARADDR_HADDR1(1) => 
        VCC_net_1, F_ARADDR_HADDR1(0) => VCC_net_1, 
        F_ARBURST_HTRANS1(1) => GND_net_1, F_ARBURST_HTRANS1(0)
         => GND_net_1, F_ARID_HSEL1(3) => GND_net_1, 
        F_ARID_HSEL1(2) => GND_net_1, F_ARID_HSEL1(1) => 
        GND_net_1, F_ARID_HSEL1(0) => GND_net_1, 
        F_ARLEN_HBURST1(3) => GND_net_1, F_ARLEN_HBURST1(2) => 
        GND_net_1, F_ARLEN_HBURST1(1) => GND_net_1, 
        F_ARLEN_HBURST1(0) => GND_net_1, F_ARLOCK_HMASTLOCK1(1)
         => GND_net_1, F_ARLOCK_HMASTLOCK1(0) => GND_net_1, 
        F_ARSIZE_HSIZE1(1) => GND_net_1, F_ARSIZE_HSIZE1(0) => 
        GND_net_1, F_ARVALID_HWRITE1 => GND_net_1, 
        F_AWADDR_HADDR0(31) => VCC_net_1, F_AWADDR_HADDR0(30) => 
        VCC_net_1, F_AWADDR_HADDR0(29) => VCC_net_1, 
        F_AWADDR_HADDR0(28) => VCC_net_1, F_AWADDR_HADDR0(27) => 
        VCC_net_1, F_AWADDR_HADDR0(26) => VCC_net_1, 
        F_AWADDR_HADDR0(25) => VCC_net_1, F_AWADDR_HADDR0(24) => 
        VCC_net_1, F_AWADDR_HADDR0(23) => VCC_net_1, 
        F_AWADDR_HADDR0(22) => VCC_net_1, F_AWADDR_HADDR0(21) => 
        VCC_net_1, F_AWADDR_HADDR0(20) => VCC_net_1, 
        F_AWADDR_HADDR0(19) => VCC_net_1, F_AWADDR_HADDR0(18) => 
        VCC_net_1, F_AWADDR_HADDR0(17) => VCC_net_1, 
        F_AWADDR_HADDR0(16) => VCC_net_1, F_AWADDR_HADDR0(15) => 
        VCC_net_1, F_AWADDR_HADDR0(14) => VCC_net_1, 
        F_AWADDR_HADDR0(13) => VCC_net_1, F_AWADDR_HADDR0(12) => 
        VCC_net_1, F_AWADDR_HADDR0(11) => VCC_net_1, 
        F_AWADDR_HADDR0(10) => VCC_net_1, F_AWADDR_HADDR0(9) => 
        VCC_net_1, F_AWADDR_HADDR0(8) => VCC_net_1, 
        F_AWADDR_HADDR0(7) => VCC_net_1, F_AWADDR_HADDR0(6) => 
        VCC_net_1, F_AWADDR_HADDR0(5) => VCC_net_1, 
        F_AWADDR_HADDR0(4) => VCC_net_1, F_AWADDR_HADDR0(3) => 
        VCC_net_1, F_AWADDR_HADDR0(2) => VCC_net_1, 
        F_AWADDR_HADDR0(1) => VCC_net_1, F_AWADDR_HADDR0(0) => 
        VCC_net_1, F_AWBURST_HTRANS0(1) => GND_net_1, 
        F_AWBURST_HTRANS0(0) => GND_net_1, F_AWID_HSEL0(3) => 
        GND_net_1, F_AWID_HSEL0(2) => GND_net_1, F_AWID_HSEL0(1)
         => GND_net_1, F_AWID_HSEL0(0) => GND_net_1, 
        F_AWLEN_HBURST0(3) => GND_net_1, F_AWLEN_HBURST0(2) => 
        GND_net_1, F_AWLEN_HBURST0(1) => GND_net_1, 
        F_AWLEN_HBURST0(0) => GND_net_1, F_AWLOCK_HMASTLOCK0(1)
         => GND_net_1, F_AWLOCK_HMASTLOCK0(0) => GND_net_1, 
        F_AWSIZE_HSIZE0(1) => GND_net_1, F_AWSIZE_HSIZE0(0) => 
        GND_net_1, F_AWVALID_HWRITE0 => GND_net_1, F_BREADY => 
        GND_net_1, F_RMW_AXI => GND_net_1, F_RREADY => GND_net_1, 
        F_WDATA_HWDATA01(63) => VCC_net_1, F_WDATA_HWDATA01(62)
         => VCC_net_1, F_WDATA_HWDATA01(61) => VCC_net_1, 
        F_WDATA_HWDATA01(60) => VCC_net_1, F_WDATA_HWDATA01(59)
         => VCC_net_1, F_WDATA_HWDATA01(58) => VCC_net_1, 
        F_WDATA_HWDATA01(57) => VCC_net_1, F_WDATA_HWDATA01(56)
         => VCC_net_1, F_WDATA_HWDATA01(55) => VCC_net_1, 
        F_WDATA_HWDATA01(54) => VCC_net_1, F_WDATA_HWDATA01(53)
         => VCC_net_1, F_WDATA_HWDATA01(52) => VCC_net_1, 
        F_WDATA_HWDATA01(51) => VCC_net_1, F_WDATA_HWDATA01(50)
         => VCC_net_1, F_WDATA_HWDATA01(49) => VCC_net_1, 
        F_WDATA_HWDATA01(48) => VCC_net_1, F_WDATA_HWDATA01(47)
         => VCC_net_1, F_WDATA_HWDATA01(46) => VCC_net_1, 
        F_WDATA_HWDATA01(45) => VCC_net_1, F_WDATA_HWDATA01(44)
         => VCC_net_1, F_WDATA_HWDATA01(43) => VCC_net_1, 
        F_WDATA_HWDATA01(42) => VCC_net_1, F_WDATA_HWDATA01(41)
         => VCC_net_1, F_WDATA_HWDATA01(40) => VCC_net_1, 
        F_WDATA_HWDATA01(39) => VCC_net_1, F_WDATA_HWDATA01(38)
         => VCC_net_1, F_WDATA_HWDATA01(37) => VCC_net_1, 
        F_WDATA_HWDATA01(36) => VCC_net_1, F_WDATA_HWDATA01(35)
         => VCC_net_1, F_WDATA_HWDATA01(34) => VCC_net_1, 
        F_WDATA_HWDATA01(33) => VCC_net_1, F_WDATA_HWDATA01(32)
         => VCC_net_1, F_WDATA_HWDATA01(31) => VCC_net_1, 
        F_WDATA_HWDATA01(30) => VCC_net_1, F_WDATA_HWDATA01(29)
         => VCC_net_1, F_WDATA_HWDATA01(28) => VCC_net_1, 
        F_WDATA_HWDATA01(27) => VCC_net_1, F_WDATA_HWDATA01(26)
         => VCC_net_1, F_WDATA_HWDATA01(25) => VCC_net_1, 
        F_WDATA_HWDATA01(24) => VCC_net_1, F_WDATA_HWDATA01(23)
         => VCC_net_1, F_WDATA_HWDATA01(22) => VCC_net_1, 
        F_WDATA_HWDATA01(21) => VCC_net_1, F_WDATA_HWDATA01(20)
         => VCC_net_1, F_WDATA_HWDATA01(19) => VCC_net_1, 
        F_WDATA_HWDATA01(18) => VCC_net_1, F_WDATA_HWDATA01(17)
         => VCC_net_1, F_WDATA_HWDATA01(16) => VCC_net_1, 
        F_WDATA_HWDATA01(15) => VCC_net_1, F_WDATA_HWDATA01(14)
         => VCC_net_1, F_WDATA_HWDATA01(13) => VCC_net_1, 
        F_WDATA_HWDATA01(12) => VCC_net_1, F_WDATA_HWDATA01(11)
         => VCC_net_1, F_WDATA_HWDATA01(10) => VCC_net_1, 
        F_WDATA_HWDATA01(9) => VCC_net_1, F_WDATA_HWDATA01(8) => 
        VCC_net_1, F_WDATA_HWDATA01(7) => VCC_net_1, 
        F_WDATA_HWDATA01(6) => VCC_net_1, F_WDATA_HWDATA01(5) => 
        VCC_net_1, F_WDATA_HWDATA01(4) => VCC_net_1, 
        F_WDATA_HWDATA01(3) => VCC_net_1, F_WDATA_HWDATA01(2) => 
        VCC_net_1, F_WDATA_HWDATA01(1) => VCC_net_1, 
        F_WDATA_HWDATA01(0) => VCC_net_1, F_WID_HREADY01(3) => 
        GND_net_1, F_WID_HREADY01(2) => GND_net_1, 
        F_WID_HREADY01(1) => GND_net_1, F_WID_HREADY01(0) => 
        GND_net_1, F_WLAST => GND_net_1, F_WSTRB(7) => GND_net_1, 
        F_WSTRB(6) => GND_net_1, F_WSTRB(5) => GND_net_1, 
        F_WSTRB(4) => GND_net_1, F_WSTRB(3) => GND_net_1, 
        F_WSTRB(2) => GND_net_1, F_WSTRB(1) => GND_net_1, 
        F_WSTRB(0) => GND_net_1, F_WVALID => GND_net_1, 
        FPGA_MDDR_ARESET_N => VCC_net_1, MDDR_FABRIC_PADDR(10)
         => CORECONFIGP_0_MDDR_APBmslave_PADDR(10), 
        MDDR_FABRIC_PADDR(9) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(9), 
        MDDR_FABRIC_PADDR(8) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(8), 
        MDDR_FABRIC_PADDR(7) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(7), 
        MDDR_FABRIC_PADDR(6) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(6), 
        MDDR_FABRIC_PADDR(5) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(5), 
        MDDR_FABRIC_PADDR(4) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(4), 
        MDDR_FABRIC_PADDR(3) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(3), 
        MDDR_FABRIC_PADDR(2) => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(2), 
        MDDR_FABRIC_PENABLE => 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE, MDDR_FABRIC_PSEL
         => CORECONFIGP_0_MDDR_APBmslave_PSELx, 
        MDDR_FABRIC_PWDATA(15) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(15), 
        MDDR_FABRIC_PWDATA(14) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(14), 
        MDDR_FABRIC_PWDATA(13) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(13), 
        MDDR_FABRIC_PWDATA(12) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(12), 
        MDDR_FABRIC_PWDATA(11) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(11), 
        MDDR_FABRIC_PWDATA(10) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(10), 
        MDDR_FABRIC_PWDATA(9) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(9), 
        MDDR_FABRIC_PWDATA(8) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(8), 
        MDDR_FABRIC_PWDATA(7) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(7), 
        MDDR_FABRIC_PWDATA(6) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(6), 
        MDDR_FABRIC_PWDATA(5) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(5), 
        MDDR_FABRIC_PWDATA(4) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(4), 
        MDDR_FABRIC_PWDATA(3) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(3), 
        MDDR_FABRIC_PWDATA(2) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(2), 
        MDDR_FABRIC_PWDATA(1) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(1), 
        MDDR_FABRIC_PWDATA(0) => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(0), 
        MDDR_FABRIC_PWRITE => CORECONFIGP_0_MDDR_APBmslave_PWRITE, 
        PRESET_N => \CORECONFIGP_0_APB_S_PRESET_N\, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_IN => GPIO_GPIO_3_BI_PAD_Y, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN => GPIO_GPIO_4_BI_PAD_Y, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_IN => GND_net_1, DM_IN(2)
         => GND_net_1, DM_IN(1) => MDDR_DM_RDQS_1_PAD_Y, DM_IN(0)
         => MDDR_DM_RDQS_0_PAD_Y, DRAM_DQ_IN(17) => GND_net_1, 
        DRAM_DQ_IN(16) => GND_net_1, DRAM_DQ_IN(15) => 
        MDDR_DQ_15_PAD_Y, DRAM_DQ_IN(14) => MDDR_DQ_14_PAD_Y, 
        DRAM_DQ_IN(13) => MDDR_DQ_13_PAD_Y, DRAM_DQ_IN(12) => 
        MDDR_DQ_12_PAD_Y, DRAM_DQ_IN(11) => MDDR_DQ_11_PAD_Y, 
        DRAM_DQ_IN(10) => MDDR_DQ_10_PAD_Y, DRAM_DQ_IN(9) => 
        MDDR_DQ_9_PAD_Y, DRAM_DQ_IN(8) => MDDR_DQ_8_PAD_Y, 
        DRAM_DQ_IN(7) => MDDR_DQ_7_PAD_Y, DRAM_DQ_IN(6) => 
        MDDR_DQ_6_PAD_Y, DRAM_DQ_IN(5) => MDDR_DQ_5_PAD_Y, 
        DRAM_DQ_IN(4) => MDDR_DQ_4_PAD_Y, DRAM_DQ_IN(3) => 
        MDDR_DQ_3_PAD_Y, DRAM_DQ_IN(2) => MDDR_DQ_2_PAD_Y, 
        DRAM_DQ_IN(1) => MDDR_DQ_1_PAD_Y, DRAM_DQ_IN(0) => 
        MDDR_DQ_0_PAD_Y, DRAM_DQS_IN(2) => GND_net_1, 
        DRAM_DQS_IN(1) => MDDR_DQS_1_PAD_Y, DRAM_DQS_IN(0) => 
        MDDR_DQS_0_PAD_Y, DRAM_FIFO_WE_IN(1) => GND_net_1, 
        DRAM_FIFO_WE_IN(0) => MDDR_DQS_TMATCH_0_IN_PAD_Y, 
        I2C0_SCL_USBC_DATA1_MGPIO31B_IN => GND_net_1, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_IN => GND_net_1, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_IN => I2C_1_SCL_PAD_Y, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_IN => I2C_1_SDA_PAD_Y, 
        MGPIO0B_IN => GPIO_GPIO_0_BI_PAD_Y, MGPIO10B_IN => 
        GND_net_1, MGPIO1B_IN => GND_net_1, MGPIO25A_IN => 
        GPIO_GPIO_25_BI_PAD_Y, MGPIO26A_IN => 
        GPIO_GPIO_26_BI_PAD_Y, MGPIO27A_IN => GND_net_1, 
        MGPIO28A_IN => GND_net_1, MGPIO29A_IN => GND_net_1, 
        MGPIO2B_IN => GND_net_1, MGPIO30A_IN => GND_net_1, 
        MGPIO31A_IN => GPIO_GPIO_31_BI_PAD_Y, MGPIO3B_IN => 
        GND_net_1, MGPIO4B_IN => GND_net_1, MGPIO5B_IN => 
        GND_net_1, MGPIO6B_IN => GND_net_1, MGPIO7B_IN => 
        GND_net_1, MGPIO8B_IN => GND_net_1, MGPIO9B_IN => 
        GND_net_1, MMUART0_CTS_USBC_DATA7_MGPIO19B_IN => 
        GND_net_1, MMUART0_DCD_MGPIO22B_IN => GND_net_1, 
        MMUART0_DSR_MGPIO20B_IN => GND_net_1, 
        MMUART0_DTR_USBC_DATA6_MGPIO18B_IN => GND_net_1, 
        MMUART0_RI_MGPIO21B_IN => GND_net_1, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_IN => GND_net_1, 
        MMUART0_RXD_USBC_STP_MGPIO28B_IN => GND_net_1, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_IN => GND_net_1, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_IN => GND_net_1, 
        MMUART1_CTS_MGPIO13B_IN => GND_net_1, 
        MMUART1_DCD_MGPIO16B_IN => GPIO_GPIO_16_BI_PAD_Y, 
        MMUART1_DSR_MGPIO14B_IN => GPIO_GPIO_14_BI_PAD_Y, 
        MMUART1_DTR_MGPIO12B_IN => GPIO_GPIO_12_BI_PAD_Y, 
        MMUART1_RI_MGPIO15B_IN => GPIO_GPIO_15_BI_PAD_Y, 
        MMUART1_RTS_MGPIO11B_IN => GND_net_1, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_IN => MMUART_1_RXD_PAD_Y, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_IN => GND_net_1, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_IN => GND_net_1, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN => GND_net_1, 
        RGMII_MDC_RMII_MDC_IN => GND_net_1, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN => GND_net_1, 
        RGMII_RX_CLK_IN => GND_net_1, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN => GND_net_1, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN => GND_net_1, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN => GND_net_1, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN => GND_net_1, 
        RGMII_RXD3_USBB_DATA4_IN => GND_net_1, RGMII_TX_CLK_IN
         => GND_net_1, RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN => 
        GND_net_1, RGMII_TXD0_RMII_TXD0_USBB_DIR_IN => GND_net_1, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_IN => GND_net_1, 
        RGMII_TXD2_USBB_DATA5_IN => GND_net_1, 
        RGMII_TXD3_USBB_DATA6_IN => GND_net_1, 
        SPI0_SCK_USBA_XCLK_IN => SPI_0_CLK_PAD_Y, 
        SPI0_SDI_USBA_DIR_MGPIO5A_IN => SPI_0_DI_PAD_Y, 
        SPI0_SDO_USBA_STP_MGPIO6A_IN => GND_net_1, 
        SPI0_SS0_USBA_NXT_MGPIO7A_IN => SPI_0_SS0_PAD_Y, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_IN => GND_net_1, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_IN => GND_net_1, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_IN => GND_net_1, 
        SPI0_SS4_MGPIO19A_IN => GND_net_1, SPI0_SS5_MGPIO20A_IN
         => GND_net_1, SPI0_SS6_MGPIO21A_IN => GND_net_1, 
        SPI0_SS7_MGPIO22A_IN => GND_net_1, SPI1_SCK_IN => 
        GND_net_1, SPI1_SDI_MGPIO11A_IN => GND_net_1, 
        SPI1_SDO_MGPIO12A_IN => GND_net_1, SPI1_SS0_MGPIO13A_IN
         => GND_net_1, SPI1_SS1_MGPIO14A_IN => GND_net_1, 
        SPI1_SS2_MGPIO15A_IN => GND_net_1, SPI1_SS3_MGPIO16A_IN
         => GND_net_1, SPI1_SS4_MGPIO17A_IN => 
        GPIO_GPIO_17_BI_PAD_Y, SPI1_SS5_MGPIO18A_IN => 
        GPIO_GPIO_18_BI_PAD_Y, SPI1_SS6_MGPIO23A_IN => GND_net_1, 
        SPI1_SS7_MGPIO24A_IN => GND_net_1, USBC_XCLK_IN => 
        GND_net_1, USBD_DATA0_IN => GND_net_1, USBD_DATA1_IN => 
        GND_net_1, USBD_DATA2_IN => GND_net_1, USBD_DATA3_IN => 
        GND_net_1, USBD_DATA4_IN => GND_net_1, USBD_DATA5_IN => 
        GND_net_1, USBD_DATA6_IN => GND_net_1, 
        USBD_DATA7_MGPIO23B_IN => GND_net_1, USBD_DIR_IN => 
        GND_net_1, USBD_NXT_IN => GND_net_1, USBD_STP_IN => 
        GND_net_1, USBD_XCLK_IN => GND_net_1, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT => 
        MSS_ADLIB_INST_CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT => 
        MSS_ADLIB_INST_CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT => OPEN, DRAM_ADDR(15)
         => \DRAM_ADDR_net_0[15]\, DRAM_ADDR(14) => 
        \DRAM_ADDR_net_0[14]\, DRAM_ADDR(13) => 
        \DRAM_ADDR_net_0[13]\, DRAM_ADDR(12) => 
        \DRAM_ADDR_net_0[12]\, DRAM_ADDR(11) => 
        \DRAM_ADDR_net_0[11]\, DRAM_ADDR(10) => 
        \DRAM_ADDR_net_0[10]\, DRAM_ADDR(9) => 
        \DRAM_ADDR_net_0[9]\, DRAM_ADDR(8) => 
        \DRAM_ADDR_net_0[8]\, DRAM_ADDR(7) => 
        \DRAM_ADDR_net_0[7]\, DRAM_ADDR(6) => 
        \DRAM_ADDR_net_0[6]\, DRAM_ADDR(5) => 
        \DRAM_ADDR_net_0[5]\, DRAM_ADDR(4) => 
        \DRAM_ADDR_net_0[4]\, DRAM_ADDR(3) => 
        \DRAM_ADDR_net_0[3]\, DRAM_ADDR(2) => 
        \DRAM_ADDR_net_0[2]\, DRAM_ADDR(1) => 
        \DRAM_ADDR_net_0[1]\, DRAM_ADDR(0) => 
        \DRAM_ADDR_net_0[0]\, DRAM_BA(2) => \DRAM_BA_net_0[2]\, 
        DRAM_BA(1) => \DRAM_BA_net_0[1]\, DRAM_BA(0) => 
        \DRAM_BA_net_0[0]\, DRAM_CASN => MSS_ADLIB_INST_DRAM_CASN, 
        DRAM_CKE => MSS_ADLIB_INST_DRAM_CKE, DRAM_CLK => 
        MSS_ADLIB_INST_DRAM_CLK, DRAM_CSN => 
        MSS_ADLIB_INST_DRAM_CSN, DRAM_DM_RDQS_OUT(2) => nc22, 
        DRAM_DM_RDQS_OUT(1) => \DRAM_DM_RDQS_OUT_net_0[1]\, 
        DRAM_DM_RDQS_OUT(0) => \DRAM_DM_RDQS_OUT_net_0[0]\, 
        DRAM_DQ_OUT(17) => nc210, DRAM_DQ_OUT(16) => nc185, 
        DRAM_DQ_OUT(15) => \DRAM_DQ_OUT_net_0[15]\, 
        DRAM_DQ_OUT(14) => \DRAM_DQ_OUT_net_0[14]\, 
        DRAM_DQ_OUT(13) => \DRAM_DQ_OUT_net_0[13]\, 
        DRAM_DQ_OUT(12) => \DRAM_DQ_OUT_net_0[12]\, 
        DRAM_DQ_OUT(11) => \DRAM_DQ_OUT_net_0[11]\, 
        DRAM_DQ_OUT(10) => \DRAM_DQ_OUT_net_0[10]\, 
        DRAM_DQ_OUT(9) => \DRAM_DQ_OUT_net_0[9]\, DRAM_DQ_OUT(8)
         => \DRAM_DQ_OUT_net_0[8]\, DRAM_DQ_OUT(7) => 
        \DRAM_DQ_OUT_net_0[7]\, DRAM_DQ_OUT(6) => 
        \DRAM_DQ_OUT_net_0[6]\, DRAM_DQ_OUT(5) => 
        \DRAM_DQ_OUT_net_0[5]\, DRAM_DQ_OUT(4) => 
        \DRAM_DQ_OUT_net_0[4]\, DRAM_DQ_OUT(3) => 
        \DRAM_DQ_OUT_net_0[3]\, DRAM_DQ_OUT(2) => 
        \DRAM_DQ_OUT_net_0[2]\, DRAM_DQ_OUT(1) => 
        \DRAM_DQ_OUT_net_0[1]\, DRAM_DQ_OUT(0) => 
        \DRAM_DQ_OUT_net_0[0]\, DRAM_DQS_OUT(2) => nc143, 
        DRAM_DQS_OUT(1) => \DRAM_DQS_OUT_net_0[1]\, 
        DRAM_DQS_OUT(0) => \DRAM_DQS_OUT_net_0[0]\, 
        DRAM_FIFO_WE_OUT(1) => nc77, DRAM_FIFO_WE_OUT(0) => 
        \DRAM_FIFO_WE_OUT_net_0[0]\, DRAM_ODT => 
        MSS_ADLIB_INST_DRAM_ODT, DRAM_RASN => 
        MSS_ADLIB_INST_DRAM_RASN, DRAM_RSTN => 
        MSS_ADLIB_INST_DRAM_RSTN, DRAM_WEN => 
        MSS_ADLIB_INST_DRAM_WEN, I2C0_SCL_USBC_DATA1_MGPIO31B_OUT
         => OPEN, I2C0_SDA_USBC_DATA0_MGPIO30B_OUT => OPEN, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_OUT => 
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OUT, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_OUT => 
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OUT, 
        MGPIO0B_OUT => MSS_ADLIB_INST_MGPIO0B_OUT, MGPIO10B_OUT
         => OPEN, MGPIO1B_OUT => OPEN, MGPIO25A_OUT => 
        MSS_ADLIB_INST_MGPIO25A_OUT, MGPIO26A_OUT => 
        MSS_ADLIB_INST_MGPIO26A_OUT, MGPIO27A_OUT => OPEN, 
        MGPIO28A_OUT => OPEN, MGPIO29A_OUT => OPEN, MGPIO2B_OUT
         => OPEN, MGPIO30A_OUT => OPEN, MGPIO31A_OUT => 
        MSS_ADLIB_INST_MGPIO31A_OUT, MGPIO3B_OUT => OPEN, 
        MGPIO4B_OUT => OPEN, MGPIO5B_OUT => OPEN, MGPIO6B_OUT => 
        OPEN, MGPIO7B_OUT => OPEN, MGPIO8B_OUT => OPEN, 
        MGPIO9B_OUT => OPEN, MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT
         => OPEN, MMUART0_DCD_MGPIO22B_OUT => OPEN, 
        MMUART0_DSR_MGPIO20B_OUT => OPEN, 
        MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT => OPEN, 
        MMUART0_RI_MGPIO21B_OUT => OPEN, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT => OPEN, 
        MMUART0_RXD_USBC_STP_MGPIO28B_OUT => OPEN, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OUT => OPEN, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_OUT => OPEN, 
        MMUART1_CTS_MGPIO13B_OUT => OPEN, 
        MMUART1_DCD_MGPIO16B_OUT => 
        MSS_ADLIB_INST_MMUART1_DCD_MGPIO16B_OUT, 
        MMUART1_DSR_MGPIO14B_OUT => 
        MSS_ADLIB_INST_MMUART1_DSR_MGPIO14B_OUT, 
        MMUART1_DTR_MGPIO12B_OUT => 
        MSS_ADLIB_INST_MMUART1_DTR_MGPIO12B_OUT, 
        MMUART1_RI_MGPIO15B_OUT => 
        MSS_ADLIB_INST_MMUART1_RI_MGPIO15B_OUT, 
        MMUART1_RTS_MGPIO11B_OUT => OPEN, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT => OPEN, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT => OPEN, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT => 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT => OPEN, 
        RGMII_MDC_RMII_MDC_OUT => OPEN, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT => OPEN, 
        RGMII_RX_CLK_OUT => OPEN, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT => OPEN, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT => OPEN, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT => OPEN, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT => OPEN, 
        RGMII_RXD3_USBB_DATA4_OUT => OPEN, RGMII_TX_CLK_OUT => 
        OPEN, RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT => OPEN, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT => OPEN, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_OUT => OPEN, 
        RGMII_TXD2_USBB_DATA5_OUT => OPEN, 
        RGMII_TXD3_USBB_DATA6_OUT => OPEN, SPI0_SCK_USBA_XCLK_OUT
         => MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT, 
        SPI0_SDI_USBA_DIR_MGPIO5A_OUT => OPEN, 
        SPI0_SDO_USBA_STP_MGPIO6A_OUT => 
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT, 
        SPI0_SS0_USBA_NXT_MGPIO7A_OUT => 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OUT => 
        MSS_ADLIB_INST_SPI0_SS1_USBA_DATA5_MGPIO8A_OUT, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OUT => OPEN, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OUT => OPEN, 
        SPI0_SS4_MGPIO19A_OUT => OPEN, SPI0_SS5_MGPIO20A_OUT => 
        MSS_ADLIB_INST_SPI0_SS5_MGPIO20A_OUT, 
        SPI0_SS6_MGPIO21A_OUT => OPEN, SPI0_SS7_MGPIO22A_OUT => 
        OPEN, SPI1_SCK_OUT => OPEN, SPI1_SDI_MGPIO11A_OUT => OPEN, 
        SPI1_SDO_MGPIO12A_OUT => OPEN, SPI1_SS0_MGPIO13A_OUT => 
        OPEN, SPI1_SS1_MGPIO14A_OUT => OPEN, 
        SPI1_SS2_MGPIO15A_OUT => OPEN, SPI1_SS3_MGPIO16A_OUT => 
        OPEN, SPI1_SS4_MGPIO17A_OUT => 
        MSS_ADLIB_INST_SPI1_SS4_MGPIO17A_OUT, 
        SPI1_SS5_MGPIO18A_OUT => 
        MSS_ADLIB_INST_SPI1_SS5_MGPIO18A_OUT, 
        SPI1_SS6_MGPIO23A_OUT => OPEN, SPI1_SS7_MGPIO24A_OUT => 
        OPEN, USBC_XCLK_OUT => OPEN, USBD_DATA0_OUT => OPEN, 
        USBD_DATA1_OUT => OPEN, USBD_DATA2_OUT => OPEN, 
        USBD_DATA3_OUT => OPEN, USBD_DATA4_OUT => OPEN, 
        USBD_DATA5_OUT => OPEN, USBD_DATA6_OUT => OPEN, 
        USBD_DATA7_MGPIO23B_OUT => OPEN, USBD_DIR_OUT => OPEN, 
        USBD_NXT_OUT => OPEN, USBD_STP_OUT => OPEN, USBD_XCLK_OUT
         => OPEN, CAN_RXBUS_USBA_DATA1_MGPIO3A_OE => 
        MSS_ADLIB_INST_CAN_RXBUS_USBA_DATA1_MGPIO3A_OE, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE => 
        MSS_ADLIB_INST_CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OE => OPEN, DM_OE(2) => nc6, 
        DM_OE(1) => \DM_OE_net_0[1]\, DM_OE(0) => 
        \DM_OE_net_0[0]\, DRAM_DQ_OE(17) => nc109, DRAM_DQ_OE(16)
         => nc87, DRAM_DQ_OE(15) => \DRAM_DQ_OE_net_0[15]\, 
        DRAM_DQ_OE(14) => \DRAM_DQ_OE_net_0[14]\, DRAM_DQ_OE(13)
         => \DRAM_DQ_OE_net_0[13]\, DRAM_DQ_OE(12) => 
        \DRAM_DQ_OE_net_0[12]\, DRAM_DQ_OE(11) => 
        \DRAM_DQ_OE_net_0[11]\, DRAM_DQ_OE(10) => 
        \DRAM_DQ_OE_net_0[10]\, DRAM_DQ_OE(9) => 
        \DRAM_DQ_OE_net_0[9]\, DRAM_DQ_OE(8) => 
        \DRAM_DQ_OE_net_0[8]\, DRAM_DQ_OE(7) => 
        \DRAM_DQ_OE_net_0[7]\, DRAM_DQ_OE(6) => 
        \DRAM_DQ_OE_net_0[6]\, DRAM_DQ_OE(5) => 
        \DRAM_DQ_OE_net_0[5]\, DRAM_DQ_OE(4) => 
        \DRAM_DQ_OE_net_0[4]\, DRAM_DQ_OE(3) => 
        \DRAM_DQ_OE_net_0[3]\, DRAM_DQ_OE(2) => 
        \DRAM_DQ_OE_net_0[2]\, DRAM_DQ_OE(1) => 
        \DRAM_DQ_OE_net_0[1]\, DRAM_DQ_OE(0) => 
        \DRAM_DQ_OE_net_0[0]\, DRAM_DQS_OE(2) => nc123, 
        DRAM_DQS_OE(1) => \DRAM_DQS_OE_net_0[1]\, DRAM_DQS_OE(0)
         => \DRAM_DQS_OE_net_0[0]\, 
        I2C0_SCL_USBC_DATA1_MGPIO31B_OE => OPEN, 
        I2C0_SDA_USBC_DATA0_MGPIO30B_OE => OPEN, 
        I2C1_SCL_USBA_DATA4_MGPIO1A_OE => 
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OE, 
        I2C1_SDA_USBA_DATA3_MGPIO0A_OE => 
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OE, MGPIO0B_OE
         => MSS_ADLIB_INST_MGPIO0B_OE, MGPIO10B_OE => OPEN, 
        MGPIO1B_OE => OPEN, MGPIO25A_OE => 
        MSS_ADLIB_INST_MGPIO25A_OE, MGPIO26A_OE => 
        MSS_ADLIB_INST_MGPIO26A_OE, MGPIO27A_OE => OPEN, 
        MGPIO28A_OE => OPEN, MGPIO29A_OE => OPEN, MGPIO2B_OE => 
        OPEN, MGPIO30A_OE => OPEN, MGPIO31A_OE => 
        MSS_ADLIB_INST_MGPIO31A_OE, MGPIO3B_OE => OPEN, 
        MGPIO4B_OE => OPEN, MGPIO5B_OE => OPEN, MGPIO6B_OE => 
        OPEN, MGPIO7B_OE => OPEN, MGPIO8B_OE => OPEN, MGPIO9B_OE
         => OPEN, MMUART0_CTS_USBC_DATA7_MGPIO19B_OE => OPEN, 
        MMUART0_DCD_MGPIO22B_OE => OPEN, MMUART0_DSR_MGPIO20B_OE
         => OPEN, MMUART0_DTR_USBC_DATA6_MGPIO18B_OE => OPEN, 
        MMUART0_RI_MGPIO21B_OE => OPEN, 
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OE => OPEN, 
        MMUART0_RXD_USBC_STP_MGPIO28B_OE => OPEN, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OE => OPEN, 
        MMUART0_TXD_USBC_DIR_MGPIO27B_OE => OPEN, 
        MMUART1_CTS_MGPIO13B_OE => OPEN, MMUART1_DCD_MGPIO16B_OE
         => MSS_ADLIB_INST_MMUART1_DCD_MGPIO16B_OE, 
        MMUART1_DSR_MGPIO14B_OE => 
        MSS_ADLIB_INST_MMUART1_DSR_MGPIO14B_OE, 
        MMUART1_DTR_MGPIO12B_OE => 
        MSS_ADLIB_INST_MMUART1_DTR_MGPIO12B_OE, 
        MMUART1_RI_MGPIO15B_OE => 
        MSS_ADLIB_INST_MMUART1_RI_MGPIO15B_OE, 
        MMUART1_RTS_MGPIO11B_OE => OPEN, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OE => OPEN, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OE => OPEN, 
        MMUART1_TXD_USBC_DATA2_MGPIO24B_OE => 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE => OPEN, 
        RGMII_MDC_RMII_MDC_OE => OPEN, 
        RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE => OPEN, 
        RGMII_RX_CLK_OE => OPEN, 
        RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE => OPEN, 
        RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE => OPEN, 
        RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE => OPEN, 
        RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE => OPEN, 
        RGMII_RXD3_USBB_DATA4_OE => OPEN, RGMII_TX_CLK_OE => OPEN, 
        RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE => OPEN, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OE => OPEN, 
        RGMII_TXD1_RMII_TXD1_USBB_STP_OE => OPEN, 
        RGMII_TXD2_USBB_DATA5_OE => OPEN, 
        RGMII_TXD3_USBB_DATA6_OE => OPEN, SPI0_SCK_USBA_XCLK_OE
         => MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE, 
        SPI0_SDI_USBA_DIR_MGPIO5A_OE => OPEN, 
        SPI0_SDO_USBA_STP_MGPIO6A_OE => 
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE, 
        SPI0_SS0_USBA_NXT_MGPIO7A_OE => 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OE => 
        MSS_ADLIB_INST_SPI0_SS1_USBA_DATA5_MGPIO8A_OE, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OE => OPEN, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OE => OPEN, 
        SPI0_SS4_MGPIO19A_OE => OPEN, SPI0_SS5_MGPIO20A_OE => 
        OPEN, SPI0_SS6_MGPIO21A_OE => OPEN, SPI0_SS7_MGPIO22A_OE
         => OPEN, SPI1_SCK_OE => OPEN, SPI1_SDI_MGPIO11A_OE => 
        OPEN, SPI1_SDO_MGPIO12A_OE => OPEN, SPI1_SS0_MGPIO13A_OE
         => OPEN, SPI1_SS1_MGPIO14A_OE => OPEN, 
        SPI1_SS2_MGPIO15A_OE => OPEN, SPI1_SS3_MGPIO16A_OE => 
        OPEN, SPI1_SS4_MGPIO17A_OE => 
        MSS_ADLIB_INST_SPI1_SS4_MGPIO17A_OE, SPI1_SS5_MGPIO18A_OE
         => MSS_ADLIB_INST_SPI1_SS5_MGPIO18A_OE, 
        SPI1_SS6_MGPIO23A_OE => OPEN, SPI1_SS7_MGPIO24A_OE => 
        OPEN, USBC_XCLK_OE => OPEN, USBD_DATA0_OE => OPEN, 
        USBD_DATA1_OE => OPEN, USBD_DATA2_OE => OPEN, 
        USBD_DATA3_OE => OPEN, USBD_DATA4_OE => OPEN, 
        USBD_DATA5_OE => OPEN, USBD_DATA6_OE => OPEN, 
        USBD_DATA7_MGPIO23B_OE => OPEN, USBD_DIR_OE => OPEN, 
        USBD_NXT_OE => OPEN, USBD_STP_OE => OPEN, USBD_XCLK_OE
         => OPEN);
    
    MDDR_RAS_N_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => MSS_ADLIB_INST_DRAM_RASN, PAD => MDDR_RAS_N);
    
    SPI_0_CLK_PAD : BIBUF
      port map(PAD => SPI_0_CLK, D => 
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT, E => 
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE, Y => 
        SPI_0_CLK_PAD_Y);
    
    MDDR_DQ_4_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(4), D => \DRAM_DQ_OUT_net_0[4]\, E
         => \DRAM_DQ_OE_net_0[4]\, Y => MDDR_DQ_4_PAD_Y);
    
    GPIO_GPIO_18_BI_PAD : BIBUF
      port map(PAD => GPIO_18_BI, D => 
        MSS_ADLIB_INST_SPI1_SS5_MGPIO18A_OUT, E => 
        MSS_ADLIB_INST_SPI1_SS5_MGPIO18A_OE, Y => 
        GPIO_GPIO_18_BI_PAD_Y);
    
    GPIO_GPIO_16_BI_PAD : BIBUF
      port map(PAD => GPIO_16_BI, D => 
        MSS_ADLIB_INST_MMUART1_DCD_MGPIO16B_OUT, E => 
        MSS_ADLIB_INST_MMUART1_DCD_MGPIO16B_OE, Y => 
        GPIO_GPIO_16_BI_PAD_Y);
    
    MDDR_ADDR_10_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[10]\, PAD => MDDR_ADDR(10));
    
    MDDR_DQS_TMATCH_0_IN_PAD : INBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQS_TMATCH_0_IN, Y => 
        MDDR_DQS_TMATCH_0_IN_PAD_Y);
    
    MDDR_CS_N_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => MSS_ADLIB_INST_DRAM_CSN, PAD => MDDR_CS_N);
    
    MDDR_ADDR_4_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[4]\, PAD => MDDR_ADDR(4));
    
    SPI_0_SS0_PAD : BIBUF
      port map(PAD => SPI_0_SS0, D => 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT, E => 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE, Y => 
        SPI_0_SS0_PAD_Y);
    
    MDDR_DQ_7_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(7), D => \DRAM_DQ_OUT_net_0[7]\, E
         => \DRAM_DQ_OE_net_0[7]\, Y => MDDR_DQ_7_PAD_Y);
    
    MDDR_WE_N_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => MSS_ADLIB_INST_DRAM_WEN, PAD => MDDR_WE_N);
    
    MDDR_ADDR_8_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[8]\, PAD => MDDR_ADDR(8));
    
    GPIO_GPIO_3_BI_PAD : BIBUF
      port map(PAD => GPIO_3_BI, D => 
        MSS_ADLIB_INST_CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT, E => 
        MSS_ADLIB_INST_CAN_RXBUS_USBA_DATA1_MGPIO3A_OE, Y => 
        GPIO_GPIO_3_BI_PAD_Y);
    
    MDDR_ADDR_15_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[15]\, PAD => MDDR_ADDR(15));
    
    MDDR_ADDR_0_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[0]\, PAD => MDDR_ADDR(0));
    
    MDDR_ADDR_1_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[1]\, PAD => MDDR_ADDR(1));
    
    GPIO_GPIO_20_OUT_PAD : OUTBUF
      port map(D => MSS_ADLIB_INST_SPI0_SS5_MGPIO20A_OUT, PAD => 
        GPIO_20_OUT);
    
    SPI_0_SS1_PAD : TRIBUFF
      port map(D => 
        MSS_ADLIB_INST_SPI0_SS1_USBA_DATA5_MGPIO8A_OUT, E => 
        MSS_ADLIB_INST_SPI0_SS1_USBA_DATA5_MGPIO8A_OE, PAD => 
        SPI_0_SS1);
    
    FIC_2_APB_M_PCLK_inferred_clock_RNIPG5 : CLKINT
      port map(A => FIC_2_APB_M_PCLK, Y => 
        \CORECONFIGP_0_APB_S_PCLK\);
    
    MDDR_DQ_13_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(13), D => \DRAM_DQ_OUT_net_0[13]\, 
        E => \DRAM_DQ_OE_net_0[13]\, Y => MDDR_DQ_13_PAD_Y);
    
    MDDR_ADDR_3_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_ADDR_net_0[3]\, PAD => MDDR_ADDR(3));
    
    MMUART_1_RXD_PAD : INBUF
      port map(PAD => MMUART_1_RXD, Y => MMUART_1_RXD_PAD_Y);
    
    MDDR_BA_0_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_BA_net_0[0]\, PAD => MDDR_BA(0));
    
    GPIO_GPIO_26_BI_PAD : BIBUF
      port map(PAD => GPIO_26_BI, D => 
        MSS_ADLIB_INST_MGPIO26A_OUT, E => 
        MSS_ADLIB_INST_MGPIO26A_OE, Y => GPIO_GPIO_26_BI_PAD_Y);
    
    MDDR_DQ_6_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(6), D => \DRAM_DQ_OUT_net_0[6]\, E
         => \DRAM_DQ_OE_net_0[6]\, Y => MDDR_DQ_6_PAD_Y);
    
    MDDR_CLK_PAD : OUTBUF_DIFF
      generic map(IOSTD => "LPDDRI")

      port map(D => MSS_ADLIB_INST_DRAM_CLK, PADP => MDDR_CLK, 
        PADN => MDDR_CLK_N);
    
    MDDR_DQ_14_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(14), D => \DRAM_DQ_OUT_net_0[14]\, 
        E => \DRAM_DQ_OE_net_0[14]\, Y => MDDR_DQ_14_PAD_Y);
    
    GPIO_GPIO_15_BI_PAD : BIBUF
      port map(PAD => GPIO_15_BI, D => 
        MSS_ADLIB_INST_MMUART1_RI_MGPIO15B_OUT, E => 
        MSS_ADLIB_INST_MMUART1_RI_MGPIO15B_OE, Y => 
        GPIO_GPIO_15_BI_PAD_Y);
    
    MDDR_DQS_TMATCH_0_OUT_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_FIFO_WE_OUT_net_0[0]\, PAD => 
        MDDR_DQS_TMATCH_0_OUT);
    
    MDDR_BA_1_PAD : OUTBUF
      generic map(IOSTD => "LVCMOS18")

      port map(D => \DRAM_BA_net_0[1]\, PAD => MDDR_BA(1));
    
    MDDR_DQ_5_PAD : BIBUF
      generic map(IOSTD => "LVCMOS18")

      port map(PAD => MDDR_DQ(5), D => \DRAM_DQ_OUT_net_0[5]\, E
         => \DRAM_DQ_OE_net_0[5]\, Y => MDDR_DQ_5_PAD_Y);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreResetP is

    port( CORECONFIGP_0_CONFIG2_DONE              : in    std_logic;
          CORECONFIGP_0_CONFIG1_DONE              : in    std_logic;
          CORECONFIGP_0_APB_S_PRESET_N            : in    std_logic;
          m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F : in    std_logic;
          m2s010_som_sb_0_POWER_ON_RESET_N        : in    std_logic;
          INIT_DONE                               : out   std_logic;
          FABOSC_0_RCOSC_25_50MHZ_O2F             : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz               : in    std_logic
        );

end CoreResetP;

architecture DEF_ARCH of CoreResetP is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \sm0_areset_n_rcosc\, sm0_areset_n_rcosc_0, 
        \sm0_areset_n_clk_base\, sm0_areset_n_clk_base_0, 
        \count_ddr[0]_net_1\, \count_ddr_s[0]\, \mss_ready_state\, 
        VCC_net_1, \POWER_ON_RESET_N_clk_base\, 
        \RESET_N_M2F_clk_base\, GND_net_1, \ddr_settled\, 
        \un14_count_ddr\, \count_ddr_enable\, 
        next_count_ddr_enable_0_sqmuxa, 
        \un1_next_ddr_ready_0_sqmuxa\, \mss_ready_select\, 
        \un6_fic_2_apb_m_preset_n_clk_base\, \sm0_state[0]_net_1\, 
        \sm0_state[6]_net_1\, \sm0_state[5]_net_1\, 
        \sm0_state[4]_net_1\, \sm0_state_ns[2]_net_1\, 
        \sm0_state[3]_net_1\, \sm0_state_ns[3]_net_1\, 
        \sm0_state[2]_net_1\, \sm0_state_ns[4]_net_1\, 
        \sm0_state[1]_net_1\, \sm0_state_ns[5]_net_1\, 
        \sm0_state_ns_a3[6]_net_1\, \MSS_HPMS_READY_int\, 
        \MSS_HPMS_READY_int_3\, sm0_areset_n_rcosc_q1, 
        sm0_areset_n_i_i, \release_sdif0_core_q1\, 
        \release_sdif0_core\, \POWER_ON_RESET_N_q1\, 
        \RESET_N_M2F_q1\, \FIC_2_APB_M_PRESET_N_q1\, 
        \sdif3_spll_lock_q1\, \count_ddr_enable_rcosc\, 
        \count_ddr_enable_q1\, \ddr_settled_clk_base\, 
        \ddr_settled_q1\, \release_sdif0_core_clk_base\, 
        \FIC_2_APB_M_PRESET_N_clk_base\, \sm0_areset_n_q1\, 
        \CONFIG1_DONE_clk_base\, \CONFIG1_DONE_q1\, 
        \CONFIG2_DONE_clk_base\, \CONFIG2_DONE_q1\, 
        \sdif3_spll_lock_q2\, \count_ddr[1]_net_1\, 
        \count_ddr_s[1]\, \count_ddr[2]_net_1\, \count_ddr_s[2]\, 
        \count_ddr[3]_net_1\, \count_ddr_s[3]\, 
        \count_ddr[4]_net_1\, \count_ddr_s[4]\, 
        \count_ddr[5]_net_1\, \count_ddr_s[5]\, 
        \count_ddr[6]_net_1\, \count_ddr_s[6]\, 
        \count_ddr[7]_net_1\, \count_ddr_s[7]\, 
        \count_ddr[8]_net_1\, \count_ddr_s[8]\, 
        \count_ddr[9]_net_1\, \count_ddr_s[9]\, 
        \count_ddr[10]_net_1\, \count_ddr_s[10]\, 
        \count_ddr[11]_net_1\, \count_ddr_s[11]\, 
        \count_ddr[12]_net_1\, \count_ddr_s[12]\, 
        \count_ddr[13]_net_1\, \count_ddr_s[13]_net_1\, 
        count_ddr_s_915_FCO, \count_ddr_cry[1]_net_1\, 
        \count_ddr_cry[2]_net_1\, \count_ddr_cry[3]_net_1\, 
        \count_ddr_cry[4]_net_1\, \count_ddr_cry[5]_net_1\, 
        \count_ddr_cry[6]_net_1\, \count_ddr_cry[7]_net_1\, 
        \count_ddr_cry[8]_net_1\, \count_ddr_cry[9]_net_1\, 
        \count_ddr_cry[10]_net_1\, \count_ddr_cry[11]_net_1\, 
        \count_ddr_cry[12]_net_1\, \un14_count_ddr_6\, 
        \un8_ddr_settled_clk_base\, \un14_count_ddr_9\, 
        \un14_count_ddr_8\, \un14_count_ddr_7\ : std_logic;

begin 


    un14_count_ddr : CFG4
      generic map(INIT => x"8000")

      port map(A => \un14_count_ddr_7\, B => \un14_count_ddr_6\, 
        C => \un14_count_ddr_8\, D => \un14_count_ddr_9\, Y => 
        \un14_count_ddr\);
    
    \sm0_state_ns[4]\ : CFG4
      generic map(INIT => x"FF70")

      port map(A => \release_sdif0_core_clk_base\, B => 
        \ddr_settled_clk_base\, C => \sm0_state[2]_net_1\, D => 
        next_count_ddr_enable_0_sqmuxa, Y => 
        \sm0_state_ns[4]_net_1\);
    
    sm0_areset_n_rcosc : SLE
      port map(D => sm0_areset_n_rcosc_q1, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => VCC_net_1, ALn => 
        sm0_areset_n_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        sm0_areset_n_rcosc_0);
    
    \count_ddr[3]\ : SLE
      port map(D => \count_ddr_s[3]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[3]_net_1\);
    
    sm0_areset_n_q1 : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => sm0_areset_n_i_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sm0_areset_n_q1\);
    
    MSS_HPMS_READY_int_RNINOKG : CFG2
      generic map(INIT => x"8")

      port map(A => \MSS_HPMS_READY_int\, B => 
        m2s010_som_sb_0_POWER_ON_RESET_N, Y => sm0_areset_n_i_i);
    
    count_ddr_enable_q1 : SLE
      port map(D => \count_ddr_enable\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => VCC_net_1, ALn => 
        \sm0_areset_n_rcosc\, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \count_ddr_enable_q1\);
    
    \sm0_state[6]\ : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => \sm0_areset_n_clk_base\, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sm0_state[6]_net_1\);
    
    \sm0_state[2]\ : SLE
      port map(D => \sm0_state_ns[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sm0_state[2]_net_1\);
    
    FIC_2_APB_M_PRESET_N_clk_base : SLE
      port map(D => \FIC_2_APB_M_PRESET_N_q1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \FIC_2_APB_M_PRESET_N_clk_base\);
    
    \count_ddr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[3]_net_1\, S => \count_ddr_s[4]\, Y => 
        OPEN, FCO => \count_ddr_cry[4]_net_1\);
    
    un8_ddr_settled_clk_base : CFG2
      generic map(INIT => x"8")

      port map(A => \ddr_settled_clk_base\, B => 
        \release_sdif0_core_clk_base\, Y => 
        \un8_ddr_settled_clk_base\);
    
    INIT_DONE_int : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \sm0_state[0]_net_1\, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        INIT_DONE);
    
    \count_ddr[9]\ : SLE
      port map(D => \count_ddr_s[9]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[9]_net_1\);
    
    MSS_HPMS_READY_int : SLE
      port map(D => \MSS_HPMS_READY_int_3\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \POWER_ON_RESET_N_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \MSS_HPMS_READY_int\);
    
    count_ddr_enable_rcosc : SLE
      port map(D => \count_ddr_enable_q1\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => VCC_net_1, ALn => 
        \sm0_areset_n_rcosc\, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \count_ddr_enable_rcosc\);
    
    sm0_areset_n_clk_base_RNIEFM9 : CLKINT
      port map(A => sm0_areset_n_clk_base_0, Y => 
        \sm0_areset_n_clk_base\);
    
    \count_ddr[7]\ : SLE
      port map(D => \count_ddr_s[7]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[7]_net_1\);
    
    \sm0_state_ns_a3[6]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \CONFIG2_DONE_clk_base\, B => 
        \sm0_state[1]_net_1\, Y => \sm0_state_ns_a3[6]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sm0_state[4]\ : SLE
      port map(D => \sm0_state_ns[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sm0_state[4]_net_1\);
    
    MSS_HPMS_READY_int_3 : CFG3
      generic map(INIT => x"E0")

      port map(A => \RESET_N_M2F_clk_base\, B => 
        \mss_ready_select\, C => \FIC_2_APB_M_PRESET_N_clk_base\, 
        Y => \MSS_HPMS_READY_int_3\);
    
    count_ddr_enable : SLE
      port map(D => next_count_ddr_enable_0_sqmuxa, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        \un1_next_ddr_ready_0_sqmuxa\, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \count_ddr_enable\);
    
    \count_ddr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[9]_net_1\, S => \count_ddr_s[10]\, Y => 
        OPEN, FCO => \count_ddr_cry[10]_net_1\);
    
    \sm0_state[5]\ : SLE
      port map(D => \sm0_state[6]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sm0_state[5]_net_1\);
    
    \count_ddr_cry[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[10]_net_1\, S => \count_ddr_s[11]\, Y => 
        OPEN, FCO => \count_ddr_cry[11]_net_1\);
    
    \count_ddr[8]\ : SLE
      port map(D => \count_ddr_s[8]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[8]_net_1\);
    
    \sm0_state_ns[2]\ : CFG3
      generic map(INIT => x"AE")

      port map(A => \sm0_state[5]_net_1\, B => 
        \sm0_state[4]_net_1\, C => \CONFIG1_DONE_clk_base\, Y => 
        \sm0_state_ns[2]_net_1\);
    
    sm0_areset_n_clk_base : SLE
      port map(D => \sm0_areset_n_q1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        sm0_areset_n_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        sm0_areset_n_clk_base_0);
    
    \count_ddr_cry[12]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[12]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[11]_net_1\, S => \count_ddr_s[12]\, Y => 
        OPEN, FCO => \count_ddr_cry[12]_net_1\);
    
    mss_ready_state : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \RESET_N_M2F_clk_base\, ALn => 
        \POWER_ON_RESET_N_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mss_ready_state\);
    
    \sm0_state[1]\ : SLE
      port map(D => \sm0_state_ns[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sm0_state[1]_net_1\);
    
    next_count_ddr_enable_0_sqmuxa_0_a3 : CFG2
      generic map(INIT => x"8")

      port map(A => \sdif3_spll_lock_q2\, B => 
        \sm0_state[3]_net_1\, Y => next_count_ddr_enable_0_sqmuxa);
    
    count_ddr_s_915 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => count_ddr_s_915_FCO);
    
    ddr_settled_clk_base : SLE
      port map(D => \ddr_settled_q1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ddr_settled_clk_base\);
    
    FIC_2_APB_M_PRESET_N_q1 : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \FIC_2_APB_M_PRESET_N_q1\);
    
    un14_count_ddr_7 : CFG4
      generic map(INIT => x"8000")

      port map(A => \count_ddr[10]_net_1\, B => 
        \count_ddr[9]_net_1\, C => \count_ddr[8]_net_1\, D => 
        \count_ddr[4]_net_1\, Y => \un14_count_ddr_7\);
    
    \count_ddr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[7]_net_1\, S => \count_ddr_s[8]\, Y => 
        OPEN, FCO => \count_ddr_cry[8]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \count_ddr_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \count_ddr[0]_net_1\, Y => \count_ddr_s[0]\);
    
    POWER_ON_RESET_N_clk_base : SLE
      port map(D => \POWER_ON_RESET_N_q1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        m2s010_som_sb_0_POWER_ON_RESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \POWER_ON_RESET_N_clk_base\);
    
    \count_ddr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => count_ddr_s_915_FCO, S
         => \count_ddr_s[1]\, Y => OPEN, FCO => 
        \count_ddr_cry[1]_net_1\);
    
    RESET_N_M2F_q1 : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => 
        m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \RESET_N_M2F_q1\);
    
    release_sdif0_core_q1 : SLE
      port map(D => \release_sdif0_core\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \release_sdif0_core_q1\);
    
    \count_ddr[10]\ : SLE
      port map(D => \count_ddr_s[10]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[10]_net_1\);
    
    \count_ddr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[5]_net_1\, S => \count_ddr_s[6]\, Y => 
        OPEN, FCO => \count_ddr_cry[6]_net_1\);
    
    \count_ddr_s[13]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[13]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[12]_net_1\, S => \count_ddr_s[13]_net_1\, 
        Y => OPEN, FCO => OPEN);
    
    \count_ddr[5]\ : SLE
      port map(D => \count_ddr_s[5]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[5]_net_1\);
    
    \count_ddr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[2]_net_1\, S => \count_ddr_s[3]\, Y => 
        OPEN, FCO => \count_ddr_cry[3]_net_1\);
    
    \count_ddr[2]\ : SLE
      port map(D => \count_ddr_s[2]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[2]_net_1\);
    
    sdif0_areset_n_rcosc_q1 : SLE
      port map(D => VCC_net_1, CLK => FABOSC_0_RCOSC_25_50MHZ_O2F, 
        EN => VCC_net_1, ALn => sm0_areset_n_i_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => sm0_areset_n_rcosc_q1);
    
    \count_ddr[1]\ : SLE
      port map(D => \count_ddr_s[1]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[1]_net_1\);
    
    \sm0_state[0]\ : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \sm0_state_ns_a3[6]_net_1\, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sm0_state[0]_net_1\);
    
    un14_count_ddr_8 : CFG4
      generic map(INIT => x"0001")

      port map(A => \count_ddr[7]_net_1\, B => 
        \count_ddr[6]_net_1\, C => \count_ddr[5]_net_1\, D => 
        \count_ddr[3]_net_1\, Y => \un14_count_ddr_8\);
    
    \count_ddr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[1]_net_1\, S => \count_ddr_s[2]\, Y => 
        OPEN, FCO => \count_ddr_cry[2]_net_1\);
    
    \count_ddr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[4]_net_1\, S => \count_ddr_s[5]\, Y => 
        OPEN, FCO => \count_ddr_cry[5]_net_1\);
    
    ddr_settled_q1 : SLE
      port map(D => \ddr_settled\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ddr_settled_q1\);
    
    \count_ddr[11]\ : SLE
      port map(D => \count_ddr_s[11]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[11]_net_1\);
    
    un14_count_ddr_9 : CFG4
      generic map(INIT => x"0001")

      port map(A => \count_ddr[12]_net_1\, B => 
        \count_ddr[11]_net_1\, C => \count_ddr[2]_net_1\, D => 
        \count_ddr[1]_net_1\, Y => \un14_count_ddr_9\);
    
    \sm0_state[3]\ : SLE
      port map(D => \sm0_state_ns[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sm0_state[3]_net_1\);
    
    \sm0_state_ns[3]\ : CFG4
      generic map(INIT => x"F222")

      port map(A => \sm0_state[3]_net_1\, B => 
        \sdif3_spll_lock_q2\, C => \sm0_state[4]_net_1\, D => 
        \CONFIG1_DONE_clk_base\, Y => \sm0_state_ns[3]_net_1\);
    
    \count_ddr[0]\ : SLE
      port map(D => \count_ddr_s[0]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[0]_net_1\);
    
    CONFIG2_DONE_q1 : SLE
      port map(D => CORECONFIGP_0_CONFIG2_DONE, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \CONFIG2_DONE_q1\);
    
    CONFIG2_DONE_clk_base : SLE
      port map(D => \CONFIG2_DONE_q1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \CONFIG2_DONE_clk_base\);
    
    CONFIG1_DONE_clk_base : SLE
      port map(D => \CONFIG1_DONE_q1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \CONFIG1_DONE_clk_base\);
    
    sm0_areset_n_rcosc_RNIKFSA : CLKINT
      port map(A => sm0_areset_n_rcosc_0, Y => 
        \sm0_areset_n_rcosc\);
    
    mss_ready_select : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \un6_fic_2_apb_m_preset_n_clk_base\, ALn => 
        \POWER_ON_RESET_N_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \mss_ready_select\);
    
    un6_fic_2_apb_m_preset_n_clk_base : CFG2
      generic map(INIT => x"8")

      port map(A => \FIC_2_APB_M_PRESET_N_clk_base\, B => 
        \mss_ready_state\, Y => 
        \un6_fic_2_apb_m_preset_n_clk_base\);
    
    \count_ddr[4]\ : SLE
      port map(D => \count_ddr_s[4]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[4]_net_1\);
    
    \count_ddr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[6]_net_1\, S => \count_ddr_s[7]\, Y => 
        OPEN, FCO => \count_ddr_cry[7]_net_1\);
    
    release_sdif0_core : SLE
      port map(D => VCC_net_1, CLK => FABOSC_0_RCOSC_25_50MHZ_O2F, 
        EN => VCC_net_1, ALn => \sm0_areset_n_rcosc\, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \release_sdif0_core\);
    
    POWER_ON_RESET_N_q1 : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => m2s010_som_sb_0_POWER_ON_RESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \POWER_ON_RESET_N_q1\);
    
    \count_ddr[12]\ : SLE
      port map(D => \count_ddr_s[12]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[12]_net_1\);
    
    ddr_settled : SLE
      port map(D => VCC_net_1, CLK => FABOSC_0_RCOSC_25_50MHZ_O2F, 
        EN => \un14_count_ddr\, ALn => \sm0_areset_n_rcosc\, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \ddr_settled\);
    
    \count_ddr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \count_ddr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \count_ddr_cry[8]_net_1\, S => \count_ddr_s[9]\, Y => 
        OPEN, FCO => \count_ddr_cry[9]_net_1\);
    
    \count_ddr[6]\ : SLE
      port map(D => \count_ddr_s[6]\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[6]_net_1\);
    
    CONFIG1_DONE_q1 : SLE
      port map(D => CORECONFIGP_0_CONFIG1_DONE, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \CONFIG1_DONE_q1\);
    
    un14_count_ddr_6 : CFG2
      generic map(INIT => x"4")

      port map(A => \count_ddr[0]_net_1\, B => 
        \count_ddr[13]_net_1\, Y => \un14_count_ddr_6\);
    
    sdif3_spll_lock_q1 : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => \sm0_areset_n_clk_base\, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \sdif3_spll_lock_q1\);
    
    release_sdif0_core_clk_base : SLE
      port map(D => \release_sdif0_core_q1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \release_sdif0_core_clk_base\);
    
    sdif3_spll_lock_q2 : SLE
      port map(D => \sdif3_spll_lock_q1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        \sm0_areset_n_clk_base\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sdif3_spll_lock_q2\);
    
    RESET_N_M2F_clk_base : SLE
      port map(D => \RESET_N_M2F_q1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \RESET_N_M2F_clk_base\);
    
    un1_next_ddr_ready_0_sqmuxa : CFG4
      generic map(INIT => x"F888")

      port map(A => \sdif3_spll_lock_q2\, B => 
        \sm0_state[3]_net_1\, C => \ddr_settled_clk_base\, D => 
        \sm0_state[2]_net_1\, Y => \un1_next_ddr_ready_0_sqmuxa\);
    
    \count_ddr[13]\ : SLE
      port map(D => \count_ddr_s[13]_net_1\, CLK => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, EN => 
        \count_ddr_enable_rcosc\, ALn => \sm0_areset_n_rcosc\, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \count_ddr[13]_net_1\);
    
    \sm0_state_ns[5]\ : CFG4
      generic map(INIT => x"F444")

      port map(A => \CONFIG2_DONE_clk_base\, B => 
        \sm0_state[1]_net_1\, C => \un8_ddr_settled_clk_base\, D
         => \sm0_state[2]_net_1\, Y => \sm0_state_ns[5]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb_GPIO_6_IO is

    port( GPIO_6_PAD_0                      : inout std_logic := 'Z';
          GPIO_6_Y_0                        : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_6_M2F_OE : in    std_logic;
          m2s010_som_sb_MSS_0_GPIO_6_M2F    : in    std_logic
        );

end m2s010_som_sb_GPIO_6_IO;

architecture DEF_ARCH of m2s010_som_sb_GPIO_6_IO is 

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    U0_0 : BIBUF
      generic map(IOSTD => "LVCMOS33")

      port map(PAD => GPIO_6_PAD_0, D => 
        m2s010_som_sb_MSS_0_GPIO_6_M2F, E => 
        m2s010_som_sb_MSS_0_GPIO_6_M2F_OE, Y => GPIO_6_Y_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CoreConfigP is

    port( CORECONFIGP_0_MDDR_APBmslave_PRDATA              : in    std_logic_vector(15 downto 0);
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR   : in    std_logic_vector(15 downto 2);
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA  : out   std_logic_vector(17 downto 0);
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA  : in    std_logic_vector(16 downto 0);
          CORECONFIGP_0_MDDR_APBmslave_PADDR               : out   std_logic_vector(10 downto 2);
          CORECONFIGP_0_MDDR_APBmslave_PWDATA              : out   std_logic_vector(15 downto 0);
          CORECONFIGP_0_MDDR_APBmslave_PSLVERR             : in    std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx   : in    std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE : in    std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PREADY              : in    std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PSELx               : out   std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PENABLE             : out   std_logic;
          INIT_DONE                                        : in    std_logic;
          CORECONFIGP_0_APB_S_PCLK_i                       : in    std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE  : in    std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PWRITE              : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY  : out   std_logic;
          CORECONFIGP_0_CONFIG2_DONE                       : out   std_logic;
          CORECONFIGP_0_CONFIG1_DONE                       : out   std_logic;
          CORECONFIGP_0_APB_S_PCLK                         : in    std_logic;
          CORECONFIGP_0_APB_S_PRESET_N                     : in    std_logic
        );

end CoreConfigP;

architecture DEF_ARCH of CoreConfigP is 

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \state_d[2]\, GND_net_1, \paddr[12]_net_1\, 
        \paddr_60\, \paddr[13]_net_1\, \paddr_61\, 
        \paddr[15]_net_1\, \paddr_63\, 
        \CORECONFIGP_0_CONFIG1_DONE\, \un8_int_psel\, 
        \CORECONFIGP_0_CONFIG2_DONE\, \prdata[13]\, 
        \state[1]_net_1\, \prdata[14]\, \prdata[15]\, 
        \prdata[16]\, \int_prdata_5_sqmuxa\, 
        \soft_reset_reg[15]_net_1\, \un17_int_psel\, 
        \soft_reset_reg[16]_net_1\, \prdata[0]\, \prdata[1]\, 
        \prdata[2]\, \prdata[3]\, \prdata[4]\, \prdata[5]\, 
        \prdata[6]\, \prdata[7]\, \prdata[8]\, \prdata[9]\, 
        \prdata[10]\, \prdata[11]\, \prdata[12]\, 
        \soft_reset_reg[0]_net_1\, \soft_reset_reg[1]_net_1\, 
        \soft_reset_reg[2]_net_1\, \soft_reset_reg[3]_net_1\, 
        \soft_reset_reg[4]_net_1\, \soft_reset_reg[5]_net_1\, 
        \soft_reset_reg[6]_net_1\, \soft_reset_reg[7]_net_1\, 
        \soft_reset_reg[8]_net_1\, \soft_reset_reg[9]_net_1\, 
        \soft_reset_reg[10]_net_1\, \soft_reset_reg[11]_net_1\, 
        \soft_reset_reg[12]_net_1\, \soft_reset_reg[13]_net_1\, 
        \soft_reset_reg[14]_net_1\, 
        un1_next_FIC_2_APB_M_PREADY_0_sqmuxa, pslverr, 
        \state[0]_net_1\, \state_ns[0]\, \state_ns[1]\, \psel\, 
        \state_d_i[2]\, \INIT_DONE_q2\, \INIT_DONE_q1\, 
        \MDDR_PENABLE_0_1\, \un1_fic_2_apb_m_psel\, pready, 
        int_prdata_5_sqmuxa_1, \prdata_0_iv_1_0[16]\, 
        \prdata_0_iv_1[8]\, \soft_reset_reg_m_0[9]\, 
        \soft_reset_reg_m_0[13]\, \soft_reset_reg_m_0[12]\, 
        \soft_reset_reg_m_0[7]\, \soft_reset_reg_m_0[11]\, 
        \soft_reset_reg_m_0[2]\, \soft_reset_reg_m_0[4]\, 
        \soft_reset_reg_m_0[10]\, \prdata_0_iv_1[16]_net_1\, 
        N_486, \prdata_0_iv_0_N_2L1\, \prdata_m2_0_a3\, 
        \prdata_0_iv_0_N_3L3\, 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, 
        \paddr_RNI09N31[12]_net_1\, prdata_N_14, \prdata_m9_1\, 
        \int_prdata_5_sqmuxa_0\, \un6_int_psel_1\, N_471, N_468, 
        prdata_N_9_mux, \soft_reset_reg_m[15]\, 
        \soft_reset_reg_m[14]\, \soft_reset_reg_m[3]\, 
        \soft_reset_reg_m[6]\, \soft_reset_reg_m[0]\, 
        prdata_N_12_mux : std_logic;

begin 

    CORECONFIGP_0_MDDR_APBmslave_PSELx <= 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\;
    CORECONFIGP_0_CONFIG2_DONE <= \CORECONFIGP_0_CONFIG2_DONE\;
    CORECONFIGP_0_CONFIG1_DONE <= \CORECONFIGP_0_CONFIG1_DONE\;

    int_prdata_4_sqmuxa_s : CFG3
      generic map(INIT => x"2A")

      port map(A => N_471, B => \paddr[15]_net_1\, C => \psel\, Y
         => \prdata_0_iv_1[16]_net_1\);
    
    \state[0]\ : SLE
      port map(D => \state_ns[0]\, CLK => 
        CORECONFIGP_0_APB_S_PCLK, EN => VCC_net_1, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \state[0]_net_1\);
    
    psel_RNI30HQ1 : CFG3
      generic map(INIT => x"DF")

      port map(A => \paddr_RNI09N31[12]_net_1\, B => 
        CORECONFIGP_0_MDDR_APBmslave_PREADY, C => \psel\, Y => 
        pready);
    
    \FIC_2_APB_M_PRDATA_0[9]\ : SLE
      port map(D => \prdata[9]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(9));
    
    FIC_2_APB_M_PSLVERR_0_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => CORECONFIGP_0_MDDR_APBmslave_PSLVERR, B => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, Y => pslverr);
    
    \FIC_2_APB_M_PRDATA_0[5]\ : SLE
      port map(D => \prdata[5]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(5));
    
    \paddr[5]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(5), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(5));
    
    \FIC_2_APB_M_PRDATA_0[4]\ : SLE
      port map(D => \prdata[4]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(4));
    
    \paddr[2]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(2));
    
    \FIC_2_APB_M_PRDATA_0[13]\ : SLE
      port map(D => \prdata[13]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(13));
    
    \prdata_0_iv_RNO[15]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => int_prdata_5_sqmuxa_1, B => N_486, C => N_471, 
        D => \soft_reset_reg[15]_net_1\, Y => 
        \soft_reset_reg_m[15]\);
    
    FIC_2_APB_M_PREADY_0 : SLE
      port map(D => \state[1]_net_1\, CLK => 
        CORECONFIGP_0_APB_S_PCLK, EN => 
        un1_next_FIC_2_APB_M_PREADY_0_sqmuxa, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY);
    
    \control_reg_1[1]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(1), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un8_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \CORECONFIGP_0_CONFIG2_DONE\);
    
    \pwdata[8]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(8), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(8));
    
    \prdata_0_iv[11]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => \soft_reset_reg_m_0[11]\, B => 
        \prdata_0_iv_1[16]_net_1\, C => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, D => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(11), Y => 
        \prdata[11]\);
    
    prdata_m2_0_a2 : CFG4
      generic map(INIT => x"CDEF")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), C => 
        \CORECONFIGP_0_CONFIG1_DONE\, D => \INIT_DONE_q2\, Y => 
        prdata_N_9_mux);
    
    paddr_63 : CFG3
      generic map(INIT => x"D8")

      port map(A => \state_d[2]\, B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(15), C => 
        \paddr[15]_net_1\, Y => \paddr_63\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \FIC_2_APB_M_PRDATA_0[8]\ : SLE
      port map(D => \prdata[8]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(8));
    
    \prdata_0_iv_RNO[3]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => int_prdata_5_sqmuxa_1, B => N_486, C => N_471, 
        D => \soft_reset_reg[3]_net_1\, Y => 
        \soft_reset_reg_m[3]\);
    
    \pwdata[10]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(10), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(10));
    
    \pwdata[4]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(4), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(4));
    
    \soft_reset_reg[6]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(6), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[6]_net_1\);
    
    prdata_m2_0_a3 : CFG2
      generic map(INIT => x"4")

      port map(A => \paddr[15]_net_1\, B => \paddr[13]_net_1\, Y
         => \prdata_m2_0_a3\);
    
    \FIC_2_APB_M_PRDATA_0[6]\ : SLE
      port map(D => \prdata[6]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(6));
    
    \pwdata[7]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(7), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(7));
    
    \paddr[7]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(7), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(7));
    
    \pwdata[0]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(0), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(0));
    
    \FIC_2_APB_M_PRDATA_0[16]\ : SLE
      port map(D => \prdata[16]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(16));
    
    \pwdata[13]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(13), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(13));
    
    \soft_reset_reg[3]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(3), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[3]_net_1\);
    
    \soft_reset_reg[15]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(15), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[15]_net_1\);
    
    \prdata_0_iv_RNO[11]\ : CFG4
      generic map(INIT => x"F0B0")

      port map(A => \paddr[15]_net_1\, B => \psel\, C => 
        \soft_reset_reg[11]_net_1\, D => \paddr[13]_net_1\, Y => 
        \soft_reset_reg_m_0[11]\);
    
    \paddr[12]\ : SLE
      port map(D => \paddr_60\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => VCC_net_1, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \paddr[12]_net_1\);
    
    \FIC_2_APB_M_PRDATA_0[10]\ : SLE
      port map(D => \prdata[10]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(10));
    
    psel : SLE
      port map(D => \state_d_i[2]\, CLK => 
        CORECONFIGP_0_APB_S_PCLK_i, EN => VCC_net_1, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => \psel\);
    
    \soft_reset_reg[2]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(2), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[2]_net_1\);
    
    \FIC_2_APB_M_PRDATA_0[0]\ : SLE
      port map(D => \prdata[0]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(0));
    
    \paddr[13]\ : SLE
      port map(D => \paddr_61\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => VCC_net_1, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \paddr[13]_net_1\);
    
    prdata_0_iv_0_N_3L3 : CFG2
      generic map(INIT => x"2")

      port map(A => \psel\, B => \prdata_m2_0_a3\, Y => 
        \prdata_0_iv_0_N_3L3\);
    
    \FIC_2_APB_M_PRDATA_0[7]\ : SLE
      port map(D => \prdata[7]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(7));
    
    un11_int_psel : CFG3
      generic map(INIT => x"01")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), C => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), Y => 
        N_468);
    
    \soft_reset_reg[14]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(14), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[14]_net_1\);
    
    \prdata_0_iv[3]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => CORECONFIGP_0_MDDR_APBmslave_PRDATA(3), B => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, C => 
        \soft_reset_reg_m[3]\, Y => \prdata[3]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    un6_int_psel_1 : CFG3
      generic map(INIT => x"80")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE, B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE, C => 
        \paddr[13]_net_1\, Y => \un6_int_psel_1\);
    
    \FIC_2_APB_M_PRDATA_0[15]\ : SLE
      port map(D => \prdata[15]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(15));
    
    \prdata_0_iv_RNO[14]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => int_prdata_5_sqmuxa_1, B => N_486, C => N_471, 
        D => \soft_reset_reg[14]_net_1\, Y => 
        \soft_reset_reg_m[14]\);
    
    un8_int_psel : CFG4
      generic map(INIT => x"4000")

      port map(A => \paddr[15]_net_1\, B => N_468, C => \psel\, D
         => \un6_int_psel_1\, Y => \un8_int_psel\);
    
    \soft_reset_reg[8]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(8), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[8]_net_1\);
    
    \prdata_0_iv_RNO[10]\ : CFG4
      generic map(INIT => x"F0B0")

      port map(A => \paddr[15]_net_1\, B => \psel\, C => 
        \soft_reset_reg[10]_net_1\, D => \paddr[13]_net_1\, Y => 
        \soft_reset_reg_m_0[10]\);
    
    \prdata_0_iv[10]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => \soft_reset_reg_m_0[10]\, B => 
        \prdata_0_iv_1[16]_net_1\, C => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, D => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(10), Y => 
        \prdata[10]\);
    
    un20_int_psel : CFG3
      generic map(INIT => x"02")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), C => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), Y => 
        N_471);
    
    un1_next_FIC_2_APB_M_PREADY_0_sqmuxa_0 : CFG4
      generic map(INIT => x"ECA0")

      port map(A => \un1_fic_2_apb_m_psel\, B => \state[1]_net_1\, 
        C => \state_d[2]\, D => pready, Y => 
        un1_next_FIC_2_APB_M_PREADY_0_sqmuxa);
    
    \prdata_0_iv_RNO[6]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => int_prdata_5_sqmuxa_1, B => N_486, C => N_471, 
        D => \soft_reset_reg[6]_net_1\, Y => 
        \soft_reset_reg_m[6]\);
    
    \prdata_0_iv_RNO[7]\ : CFG4
      generic map(INIT => x"F0B0")

      port map(A => \paddr[15]_net_1\, B => \psel\, C => 
        \soft_reset_reg[7]_net_1\, D => \paddr[13]_net_1\, Y => 
        \soft_reset_reg_m_0[7]\);
    
    MDDR_PENABLE_0_1 : CFG4
      generic map(INIT => x"0100")

      port map(A => \paddr[12]_net_1\, B => \paddr[13]_net_1\, C
         => \paddr[15]_net_1\, D => \state[1]_net_1\, Y => 
        \MDDR_PENABLE_0_1\);
    
    \FIC_2_APB_M_PRDATA_0[11]\ : SLE
      port map(D => \prdata[11]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(11));
    
    prdata_m6_e : CFG4
      generic map(INIT => x"135F")

      port map(A => N_468, B => N_471, C => 
        \CORECONFIGP_0_CONFIG2_DONE\, D => 
        \soft_reset_reg[1]_net_1\, Y => prdata_N_14);
    
    \soft_reset_reg[0]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(0), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[0]_net_1\);
    
    \prdata_0_iv_0[5]\ : CFG4
      generic map(INIT => x"F444")

      port map(A => \prdata_0_iv_0_N_3L3\, B => 
        \prdata_0_iv_0_N_2L1\, C => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(5), D => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, Y => \prdata[5]\);
    
    \pwdata[1]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(1), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(1));
    
    prdata_m9 : CFG4
      generic map(INIT => x"0595")

      port map(A => prdata_N_14, B => \prdata_m9_1\, C => \psel\, 
        D => \paddr[15]_net_1\, Y => \prdata[1]\);
    
    prdata_0_iv_0_N_2L1 : CFG4
      generic map(INIT => x"0A40")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), B => 
        \soft_reset_reg[5]_net_1\, C => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), Y => 
        \prdata_0_iv_0_N_2L1\);
    
    \prdata_0_iv_RNO[4]\ : CFG4
      generic map(INIT => x"F0B0")

      port map(A => \paddr[15]_net_1\, B => \psel\, C => 
        \soft_reset_reg[4]_net_1\, D => \paddr[13]_net_1\, Y => 
        \soft_reset_reg_m_0[4]\);
    
    un1_fic_2_apb_m_psel : CFG2
      generic map(INIT => x"4")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE, B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx, Y => 
        \un1_fic_2_apb_m_psel\);
    
    \prdata_0_iv_1[16]\ : CFG4
      generic map(INIT => x"BFFF")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), C => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), D => 
        int_prdata_5_sqmuxa_1, Y => \prdata_0_iv_1_0[16]\);
    
    prdata_m6 : CFG4
      generic map(INIT => x"1011")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), B => 
        prdata_N_9_mux, C => \prdata_m2_0_a3\, D => \psel\, Y => 
        prdata_N_12_mux);
    
    \soft_reset_reg[1]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(1), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[1]_net_1\);
    
    \paddr[9]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(9), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(9));
    
    un1_next_FIC_2_APB_M_PREADY_0_sqmuxa_0_a3 : CFG2
      generic map(INIT => x"8")

      port map(A => \state_d[2]\, B => \un1_fic_2_apb_m_psel\, Y
         => \state_ns[0]\);
    
    \prdata_0_iv[9]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => \soft_reset_reg_m_0[9]\, B => 
        \prdata_0_iv_1[16]_net_1\, C => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, D => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(9), Y => \prdata[9]\);
    
    \paddr[15]\ : SLE
      port map(D => \paddr_63\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => VCC_net_1, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \paddr[15]_net_1\);
    
    \prdata_0_iv_RNO[0]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => int_prdata_5_sqmuxa_1, B => N_486, C => N_471, 
        D => \soft_reset_reg[0]_net_1\, Y => 
        \soft_reset_reg_m[0]\);
    
    \prdata_0_iv[12]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => \soft_reset_reg_m_0[12]\, B => 
        \prdata_0_iv_1[16]_net_1\, C => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, D => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(12), Y => 
        \prdata[12]\);
    
    \FIC_2_APB_M_PRDATA_0[12]\ : SLE
      port map(D => \prdata[12]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(12));
    
    \control_reg_1[0]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(0), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un8_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \CORECONFIGP_0_CONFIG1_DONE\);
    
    \soft_reset_reg[5]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(5), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[5]_net_1\);
    
    \prdata_0_iv[14]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => CORECONFIGP_0_MDDR_APBmslave_PRDATA(14), B
         => \CORECONFIGP_0_MDDR_APBmslave_PSELx\, C => 
        \soft_reset_reg_m[14]\, Y => \prdata[14]\);
    
    \FIC_2_APB_M_PRDATA_0[14]\ : SLE
      port map(D => \prdata[14]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(14));
    
    psel_RNIPF3R : CFG2
      generic map(INIT => x"7")

      port map(A => \psel\, B => \paddr[15]_net_1\, Y => 
        int_prdata_5_sqmuxa_1);
    
    \paddr[3]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(3));
    
    INIT_DONE_q2 : SLE
      port map(D => \INIT_DONE_q1\, CLK => 
        CORECONFIGP_0_APB_S_PCLK, EN => VCC_net_1, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \INIT_DONE_q2\);
    
    \paddr_RNI09N31[12]\ : CFG3
      generic map(INIT => x"01")

      port map(A => \paddr[12]_net_1\, B => \paddr[13]_net_1\, C
         => \paddr[15]_net_1\, Y => \paddr_RNI09N31[12]_net_1\);
    
    state_s0_0_a2_i : CFG2
      generic map(INIT => x"E")

      port map(A => \state[1]_net_1\, B => \state[0]_net_1\, Y
         => \state_d_i[2]\);
    
    int_prdata_5_sqmuxa_0 : CFG2
      generic map(INIT => x"4")

      port map(A => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3), B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), Y => 
        \int_prdata_5_sqmuxa_0\);
    
    pwrite : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE, CLK => 
        CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWRITE);
    
    MDDR_PENABLE_0 : SLE
      port map(D => \MDDR_PENABLE_0_1\, CLK => 
        CORECONFIGP_0_APB_S_PCLK_i, EN => VCC_net_1, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE);
    
    \soft_reset_reg[10]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(10), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[10]_net_1\);
    
    \soft_reset_reg[4]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(4), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[4]_net_1\);
    
    \prdata_0_iv[13]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => \soft_reset_reg_m_0[13]\, B => 
        \prdata_0_iv_1[16]_net_1\, C => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, D => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(13), Y => 
        \prdata[13]\);
    
    \pwdata[6]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(6), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(6));
    
    \prdata_0_iv_RNO[8]\ : CFG4
      generic map(INIT => x"F0B0")

      port map(A => \paddr[15]_net_1\, B => \psel\, C => 
        \soft_reset_reg[8]_net_1\, D => \paddr[13]_net_1\, Y => 
        \prdata_0_iv_1[8]\);
    
    \prdata_0_iv[16]\ : CFG4
      generic map(INIT => x"00B3")

      port map(A => \prdata_0_iv_1[16]_net_1\, B => 
        \prdata_0_iv_1_0[16]\, C => \soft_reset_reg[16]_net_1\, D
         => N_486, Y => \prdata[16]\);
    
    \prdata_0_iv_RNO[12]\ : CFG4
      generic map(INIT => x"F0B0")

      port map(A => \paddr[15]_net_1\, B => \psel\, C => 
        \soft_reset_reg[12]_net_1\, D => \paddr[13]_net_1\, Y => 
        \soft_reset_reg_m_0[12]\);
    
    int_prdata_5_sqmuxa : CFG4
      generic map(INIT => x"0080")

      port map(A => \int_prdata_5_sqmuxa_0\, B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2), C => 
        int_prdata_5_sqmuxa_1, D => N_486, Y => 
        \int_prdata_5_sqmuxa\);
    
    int_sel_1_sqmuxa_1 : CFG3
      generic map(INIT => x"10")

      port map(A => \paddr[13]_net_1\, B => \paddr[15]_net_1\, C
         => \psel\, Y => N_486);
    
    \state_ns_0[1]\ : CFG3
      generic map(INIT => x"F2")

      port map(A => \state[1]_net_1\, B => pready, C => 
        \state[0]_net_1\, Y => \state_ns[1]\);
    
    \pwdata[11]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(11), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(11));
    
    \paddr[6]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(6), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(6));
    
    FIC_2_APB_M_PSLVERR_0 : SLE
      port map(D => pslverr, CLK => CORECONFIGP_0_APB_S_PCLK, EN
         => \state[1]_net_1\, ALn => CORECONFIGP_0_APB_S_PRESET_N, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR);
    
    \pwdata[12]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(12), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(12));
    
    \prdata_0_iv[0]\ : CFG4
      generic map(INIT => x"FEFA")

      port map(A => \soft_reset_reg_m[0]\, B => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(0), C => 
        prdata_N_12_mux, D => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, Y => \prdata[0]\);
    
    \paddr[4]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(4));
    
    \pwdata[9]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(9), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(9));
    
    \prdata_0_iv[15]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => CORECONFIGP_0_MDDR_APBmslave_PRDATA(15), B
         => \CORECONFIGP_0_MDDR_APBmslave_PSELx\, C => 
        \soft_reset_reg_m[15]\, Y => \prdata[15]\);
    
    prdata_m9_1 : CFG4
      generic map(INIT => x"1203")

      port map(A => \paddr[12]_net_1\, B => \paddr[13]_net_1\, C
         => prdata_N_14, D => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(1), Y => 
        \prdata_m9_1\);
    
    \prdata_0_iv[7]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => \soft_reset_reg_m_0[7]\, B => 
        \prdata_0_iv_1[16]_net_1\, C => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, D => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(7), Y => \prdata[7]\);
    
    \state[1]\ : SLE
      port map(D => \state_ns[1]\, CLK => 
        CORECONFIGP_0_APB_S_PCLK, EN => VCC_net_1, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \state[1]_net_1\);
    
    \soft_reset_reg[13]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(13), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[13]_net_1\);
    
    \FIC_2_APB_M_PRDATA_0[17]\ : SLE
      port map(D => \int_prdata_5_sqmuxa\, CLK => 
        CORECONFIGP_0_APB_S_PCLK, EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(17));
    
    \prdata_0_iv_RNO[2]\ : CFG4
      generic map(INIT => x"F0B0")

      port map(A => \paddr[15]_net_1\, B => \psel\, C => 
        \soft_reset_reg[2]_net_1\, D => \paddr[13]_net_1\, Y => 
        \soft_reset_reg_m_0[2]\);
    
    \pwdata[15]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(15), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(15));
    
    \pwdata[5]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(5), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(5));
    
    INIT_DONE_q1 : SLE
      port map(D => INIT_DONE, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => VCC_net_1, ALn => CORECONFIGP_0_APB_S_PRESET_N, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \INIT_DONE_q1\);
    
    state_s0_0_a2 : CFG2
      generic map(INIT => x"1")

      port map(A => \state[1]_net_1\, B => \state[0]_net_1\, Y
         => \state_d[2]\);
    
    \prdata_0_iv[6]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => CORECONFIGP_0_MDDR_APBmslave_PRDATA(6), B => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, C => 
        \soft_reset_reg_m[6]\, Y => \prdata[6]\);
    
    \prdata_0_iv[2]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => \soft_reset_reg_m_0[2]\, B => 
        \prdata_0_iv_1[16]_net_1\, C => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, D => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(2), Y => \prdata[2]\);
    
    un17_int_psel : CFG4
      generic map(INIT => x"4000")

      port map(A => \paddr[15]_net_1\, B => N_471, C => \psel\, D
         => \un6_int_psel_1\, Y => \un17_int_psel\);
    
    \prdata_0_iv[8]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => \prdata_0_iv_1[8]\, B => 
        \prdata_0_iv_1[16]_net_1\, C => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, D => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(8), Y => \prdata[8]\);
    
    \prdata_0_iv[4]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => \soft_reset_reg_m_0[4]\, B => 
        \prdata_0_iv_1[16]_net_1\, C => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\, D => 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(4), Y => \prdata[4]\);
    
    \paddr[10]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(10), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(10));
    
    paddr_61 : CFG3
      generic map(INIT => x"D8")

      port map(A => \state_d[2]\, B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(13), C => 
        \paddr[13]_net_1\, Y => \paddr_61\);
    
    \soft_reset_reg[9]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(9), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[9]_net_1\);
    
    \soft_reset_reg[11]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(11), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[11]_net_1\);
    
    \pwdata[2]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(2), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(2));
    
    \soft_reset_reg[16]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(16), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[16]_net_1\);
    
    \FIC_2_APB_M_PRDATA_0[2]\ : SLE
      port map(D => \prdata[2]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(2));
    
    \pwdata[14]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(14), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(14));
    
    \pwdata[3]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(3), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(3));
    
    \prdata_0_iv_RNO[9]\ : CFG4
      generic map(INIT => x"F0B0")

      port map(A => \paddr[15]_net_1\, B => \psel\, C => 
        \soft_reset_reg[9]_net_1\, D => \paddr[13]_net_1\, Y => 
        \soft_reset_reg_m_0[9]\);
    
    \FIC_2_APB_M_PRDATA_0[3]\ : SLE
      port map(D => \prdata[3]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(3));
    
    \paddr[8]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(8), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \state_d[2]\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(8));
    
    \FIC_2_APB_M_PRDATA_0[1]\ : SLE
      port map(D => \prdata[1]\, CLK => CORECONFIGP_0_APB_S_PCLK, 
        EN => \state[1]_net_1\, ALn => 
        CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(1));
    
    \prdata_0_iv_RNO[13]\ : CFG4
      generic map(INIT => x"F0B0")

      port map(A => \paddr[15]_net_1\, B => \psel\, C => 
        \soft_reset_reg[13]_net_1\, D => \paddr[13]_net_1\, Y => 
        \soft_reset_reg_m_0[13]\);
    
    \soft_reset_reg[7]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(7), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[7]_net_1\);
    
    \soft_reset_reg[12]\ : SLE
      port map(D => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(12), CLK
         => CORECONFIGP_0_APB_S_PCLK, EN => \un17_int_psel\, ALn
         => CORECONFIGP_0_APB_S_PRESET_N, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \soft_reset_reg[12]_net_1\);
    
    \paddr_RNI2KTI1[12]\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \paddr[12]_net_1\, B => \paddr[13]_net_1\, C
         => \paddr[15]_net_1\, D => \psel\, Y => 
        \CORECONFIGP_0_MDDR_APBmslave_PSELx\);
    
    paddr_60 : CFG3
      generic map(INIT => x"D8")

      port map(A => \state_d[2]\, B => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(12), C => 
        \paddr[12]_net_1\, Y => \paddr_60\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb_CCC_0_FCCC is

    port( m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC : in    std_logic;
          FAB_CCC_LOCK                              : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz                 : out   std_logic
        );

end m2s010_som_sb_CCC_0_FCCC;

architecture DEF_ARCH of m2s010_som_sb_CCC_0_FCCC is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CCC

            generic (INIT:std_logic_vector(209 downto 0) := "00" & x"0000000000000000000000000000000000000000000000000000"; 
        VCOFREQUENCY:real := 0.0);

    port( Y0              : out   std_logic;
          Y1              : out   std_logic;
          Y2              : out   std_logic;
          Y3              : out   std_logic;
          PRDATA          : out   std_logic_vector(7 downto 0);
          LOCK            : out   std_logic;
          BUSY            : out   std_logic;
          CLK0            : in    std_logic := 'U';
          CLK1            : in    std_logic := 'U';
          CLK2            : in    std_logic := 'U';
          CLK3            : in    std_logic := 'U';
          NGMUX0_SEL      : in    std_logic := 'U';
          NGMUX1_SEL      : in    std_logic := 'U';
          NGMUX2_SEL      : in    std_logic := 'U';
          NGMUX3_SEL      : in    std_logic := 'U';
          NGMUX0_HOLD_N   : in    std_logic := 'U';
          NGMUX1_HOLD_N   : in    std_logic := 'U';
          NGMUX2_HOLD_N   : in    std_logic := 'U';
          NGMUX3_HOLD_N   : in    std_logic := 'U';
          NGMUX0_ARST_N   : in    std_logic := 'U';
          NGMUX1_ARST_N   : in    std_logic := 'U';
          NGMUX2_ARST_N   : in    std_logic := 'U';
          NGMUX3_ARST_N   : in    std_logic := 'U';
          PLL_BYPASS_N    : in    std_logic := 'U';
          PLL_ARST_N      : in    std_logic := 'U';
          PLL_POWERDOWN_N : in    std_logic := 'U';
          GPD0_ARST_N     : in    std_logic := 'U';
          GPD1_ARST_N     : in    std_logic := 'U';
          GPD2_ARST_N     : in    std_logic := 'U';
          GPD3_ARST_N     : in    std_logic := 'U';
          PRESET_N        : in    std_logic := 'U';
          PCLK            : in    std_logic := 'U';
          PSEL            : in    std_logic := 'U';
          PENABLE         : in    std_logic := 'U';
          PWRITE          : in    std_logic := 'U';
          PADDR           : in    std_logic_vector(7 downto 2) := (others => 'U');
          PWDATA          : in    std_logic_vector(7 downto 0) := (others => 'U');
          CLK0_PAD        : in    std_logic := 'U';
          CLK1_PAD        : in    std_logic := 'U';
          CLK2_PAD        : in    std_logic := 'U';
          CLK3_PAD        : in    std_logic := 'U';
          GL0             : out   std_logic;
          GL1             : out   std_logic;
          GL2             : out   std_logic;
          GL3             : out   std_logic;
          RCOSC_25_50MHZ  : in    std_logic := 'U';
          RCOSC_1MHZ      : in    std_logic := 'U';
          XTLOSC          : in    std_logic := 'U'
        );
  end component;

    signal GL0_net, VCC_net_1, GND_net_1 : std_logic;
    signal nc8, nc7, nc6, nc2, nc5, nc4, nc3, nc1 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    GL0_INST : CLKINT
      port map(A => GL0_net, Y => m2s010_som_sb_0_CCC_71MHz);
    
    CCC_INST : CCC

              generic map(INIT => "00" & x"000007F88000044D64000318C6318C1F18C61E40404040404613",
         VCOFREQUENCY => 568.0)

      port map(Y0 => OPEN, Y1 => OPEN, Y2 => OPEN, Y3 => OPEN, 
        PRDATA(7) => nc8, PRDATA(6) => nc7, PRDATA(5) => nc6, 
        PRDATA(4) => nc2, PRDATA(3) => nc5, PRDATA(2) => nc4, 
        PRDATA(1) => nc3, PRDATA(0) => nc1, LOCK => FAB_CCC_LOCK, 
        BUSY => OPEN, CLK0 => VCC_net_1, CLK1 => VCC_net_1, CLK2
         => VCC_net_1, CLK3 => VCC_net_1, NGMUX0_SEL => GND_net_1, 
        NGMUX1_SEL => GND_net_1, NGMUX2_SEL => GND_net_1, 
        NGMUX3_SEL => GND_net_1, NGMUX0_HOLD_N => VCC_net_1, 
        NGMUX1_HOLD_N => VCC_net_1, NGMUX2_HOLD_N => VCC_net_1, 
        NGMUX3_HOLD_N => VCC_net_1, NGMUX0_ARST_N => VCC_net_1, 
        NGMUX1_ARST_N => VCC_net_1, NGMUX2_ARST_N => VCC_net_1, 
        NGMUX3_ARST_N => VCC_net_1, PLL_BYPASS_N => VCC_net_1, 
        PLL_ARST_N => VCC_net_1, PLL_POWERDOWN_N => VCC_net_1, 
        GPD0_ARST_N => VCC_net_1, GPD1_ARST_N => VCC_net_1, 
        GPD2_ARST_N => VCC_net_1, GPD3_ARST_N => VCC_net_1, 
        PRESET_N => GND_net_1, PCLK => VCC_net_1, PSEL => 
        VCC_net_1, PENABLE => VCC_net_1, PWRITE => VCC_net_1, 
        PADDR(7) => VCC_net_1, PADDR(6) => VCC_net_1, PADDR(5)
         => VCC_net_1, PADDR(4) => VCC_net_1, PADDR(3) => 
        VCC_net_1, PADDR(2) => VCC_net_1, PWDATA(7) => VCC_net_1, 
        PWDATA(6) => VCC_net_1, PWDATA(5) => VCC_net_1, PWDATA(4)
         => VCC_net_1, PWDATA(3) => VCC_net_1, PWDATA(2) => 
        VCC_net_1, PWDATA(1) => VCC_net_1, PWDATA(0) => VCC_net_1, 
        CLK0_PAD => GND_net_1, CLK1_PAD => GND_net_1, CLK2_PAD
         => GND_net_1, CLK3_PAD => GND_net_1, GL0 => GL0_net, GL1
         => OPEN, GL2 => OPEN, GL3 => OPEN, RCOSC_25_50MHZ => 
        GND_net_1, RCOSC_1MHZ => GND_net_1, XTLOSC => 
        m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb_OTH_SPI_1_SS0_IO is

    port( SPI_1_SS0_OTH_0                      : inout std_logic := 'Z';
          OTH_SPI_1_SS0_Y_0                    : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE : in    std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F    : in    std_logic
        );

end m2s010_som_sb_OTH_SPI_1_SS0_IO;

architecture DEF_ARCH of m2s010_som_sb_OTH_SPI_1_SS0_IO is 

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    U0_0 : BIBUF
      port map(PAD => SPI_1_SS0_OTH_0, D => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F, E => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE, Y => 
        OTH_SPI_1_SS0_Y_0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb_FABOSC_0_OSC is

    port( XTL                                       : in    std_logic;
          m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC : out   std_logic;
          FABOSC_0_RCOSC_25_50MHZ_O2F               : out   std_logic
        );

end m2s010_som_sb_FABOSC_0_OSC;

architecture DEF_ARCH of m2s010_som_sb_FABOSC_0_OSC is 

  component RCOSC_25_50MHZ_FAB
    port( A      : in    std_logic := 'U';
          CLKOUT : out   std_logic
        );
  end component;

  component RCOSC_25_50MHZ
    generic (FREQUENCY:real := 50.0);

    port( CLKOUT : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component XTLOSC
    generic (MODE:std_logic_vector(1 downto 0) := "11"; 
        FREQUENCY:real := 20.0);

    port( XTL    : in    std_logic := 'U';
          CLKOUT : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal N_RCOSC_25_50MHZ_CLKINT, N_RCOSC_25_50MHZ_CLKOUT, 
        GND_net_1, VCC_net_1 : std_logic;

begin 


    I_RCOSC_25_50MHZ_FAB : RCOSC_25_50MHZ_FAB
      port map(A => N_RCOSC_25_50MHZ_CLKOUT, CLKOUT => 
        N_RCOSC_25_50MHZ_CLKINT);
    
    I_RCOSC_25_50MHZ : RCOSC_25_50MHZ
      generic map(FREQUENCY => 50.0)

      port map(CLKOUT => N_RCOSC_25_50MHZ_CLKOUT);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    I_XTLOSC : XTLOSC
      generic map(MODE => "11", FREQUENCY => 20.0)

      port map(XTL => XTL, CLKOUT => 
        m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC);
    
    I_RCOSC_25_50MHZ_FAB_CLKINT : CLKINT
      port map(A => N_RCOSC_25_50MHZ_CLKINT, Y => 
        FABOSC_0_RCOSC_25_50MHZ_O2F);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som_sb is

    port( MDDR_DQS                                  : inout std_logic_vector(1 downto 0) := (others => 'Z');
          MDDR_DQ                                   : inout std_logic_vector(15 downto 0) := (others => 'Z');
          MDDR_DM_RDQS                              : inout std_logic_vector(1 downto 0) := (others => 'Z');
          MDDR_BA                                   : out   std_logic_vector(2 downto 0);
          MDDR_ADDR                                 : out   std_logic_vector(15 downto 0);
          CoreAPB3_0_APBmslave0_PADDR               : out   std_logic_vector(7 downto 0);
          m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR    : out   std_logic_vector(15 downto 12);
          CoreAPB3_0_APBmslave0_PWDATA              : out   std_logic_vector(7 downto 0);
          MAC_MII_TXD_c                             : out   std_logic_vector(3 downto 0);
          CoreAPB3_0_APBmslave0_PRDATA_m            : in    std_logic_vector(7 downto 0);
          Y_net_0                                   : in    std_logic_vector(3 downto 0);
          MAC_MII_RXD_c                             : in    std_logic_vector(3 downto 0);
          SPI_1_SS0_OTH_0                           : inout std_logic := 'Z';
          DEBOUNCE_OUT_net_0_0                      : in    std_logic;
          GPIO_7_PADI_0                             : inout std_logic := 'Z';
          GPIO_6_PAD_0                              : inout std_logic := 'Z';
          GPIO_1_BI_0                               : inout std_logic := 'Z';
          SPI_1_SS0_CAM_0                           : inout std_logic := 'Z';
          SPI_1_CLK_0                               : inout std_logic := 'Z';
          SPI_0_SS1                                 : out   std_logic;
          SPI_0_SS0                                 : inout std_logic := 'Z';
          SPI_0_DO                                  : out   std_logic;
          SPI_0_DI                                  : in    std_logic;
          SPI_0_CLK                                 : inout std_logic := 'Z';
          MMUART_1_TXD                              : out   std_logic;
          MMUART_1_RXD                              : in    std_logic;
          MDDR_WE_N                                 : out   std_logic;
          MDDR_RESET_N                              : out   std_logic;
          MDDR_RAS_N                                : out   std_logic;
          MDDR_ODT                                  : out   std_logic;
          MDDR_DQS_TMATCH_0_OUT                     : out   std_logic;
          MDDR_DQS_TMATCH_0_IN                      : in    std_logic;
          MDDR_CS_N                                 : out   std_logic;
          MDDR_CKE                                  : out   std_logic;
          MDDR_CAS_N                                : out   std_logic;
          I2C_1_SDA                                 : inout std_logic := 'Z';
          I2C_1_SCL                                 : inout std_logic := 'Z';
          GPIO_31_BI                                : inout std_logic := 'Z';
          GPIO_26_BI                                : inout std_logic := 'Z';
          GPIO_25_BI                                : inout std_logic := 'Z';
          GPIO_20_OUT                               : out   std_logic;
          GPIO_18_BI                                : inout std_logic := 'Z';
          GPIO_17_BI                                : inout std_logic := 'Z';
          GPIO_16_BI                                : inout std_logic := 'Z';
          GPIO_15_BI                                : inout std_logic := 'Z';
          GPIO_14_BI                                : inout std_logic := 'Z';
          GPIO_12_BI                                : inout std_logic := 'Z';
          GPIO_4_BI                                 : inout std_logic := 'Z';
          GPIO_3_BI                                 : inout std_logic := 'Z';
          GPIO_0_BI                                 : inout std_logic := 'Z';
          CoreAPB3_0_APBmslave0_PENABLE             : out   std_logic;
          m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx    : out   std_logic;
          CoreAPB3_0_APBmslave0_PWRITE              : out   std_logic;
          MAC_MII_MDC_c                             : out   std_logic;
          GPIO_22_M2F_c                             : out   std_logic;
          GPIO_21_M2F_c                             : out   std_logic;
          m2s010_som_sb_0_GPIO_28_SW_RESET          : out   std_logic;
          MMUART_0_TXD_M2F_c                        : out   std_logic;
          GPIO_24_M2F_c                             : out   std_logic;
          GPIO_5_M2F_c                              : out   std_logic;
          GPIO_8_M2F_c                              : out   std_logic;
          GPIO_11_M2F_c                             : out   std_logic;
          MAC_MII_TX_EN_c                           : out   std_logic;
          MAC_MII_COL_c                             : in    std_logic;
          MAC_MII_CRS_c                             : in    std_logic;
          CommsFPGA_top_0_INT                       : in    std_logic;
          CoreAPB3_0_APBmslave0_PREADY_i_m_i        : in    std_logic;
          DEBOUNCE_OUT_1_c                          : in    std_logic;
          DEBOUNCE_OUT_2_c                          : in    std_logic;
          MMUART_0_RXD_F2M_c                        : in    std_logic;
          MAC_MII_RX_CLK_c                          : in    std_logic;
          MAC_MII_RX_DV_c                           : in    std_logic;
          MAC_MII_RX_ER_c                           : in    std_logic;
          MAC_MII_TX_CLK_c                          : in    std_logic;
          MDDR_CLK_N                                : out   std_logic;
          MDDR_CLK                                  : out   std_logic;
          XTL                                       : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz                 : out   std_logic;
          m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC : inout std_logic := 'Z';
          SPI_1_DI_CAM_c                            : in    std_logic;
          SPI_1_DI_OTH_c                            : in    std_logic;
          CommsFPGA_top_0_CAMERA_NODE               : in    std_logic;
          DEVRST_N                                  : in    std_logic;
          m2s010_som_sb_0_POWER_ON_RESET_N          : out   std_logic;
          MAC_MII_MDIO                              : inout std_logic := 'Z';
          SPI_1_DO_CAM_c                            : inout std_logic := 'Z';
          SPI_1_DO_OTH                              : out   std_logic
        );

end m2s010_som_sb;

architecture DEF_ARCH of m2s010_som_sb is 

  component m2s010_som_sb_GPIO_1_IO
    port( GPIO_1_BI_0                       : inout   std_logic;
          GPIO_1_in_0                       : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_1_M2F_OE : in    std_logic := 'U';
          GPIO_1_M2F                        : in    std_logic := 'U'
        );
  end component;

  component m2s010_som_sb_CAM_SPI_1_CLK_IO
    port( CAM_SPI_1_CLK_Y_0                    : out   std_logic;
          SPI_1_CLK_0                          : inout   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE : in    std_logic := 'U';
          m2s010_som_sb_MSS_0_SPI_1_CLK_M2F    : in    std_logic := 'U'
        );
  end component;

  component m2s010_som_sb_GPIO_7_IO
    port( GPIO_7_PADI_0                     : inout   std_logic;
          GPIO_7_Y_0                        : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_7_M2F_OE : in    std_logic := 'U';
          m2s010_som_sb_MSS_0_GPIO_7_M2F    : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component m2s010_som_sb_CAM_SPI_1_SS0_IO
    port( SPI_1_SS0_CAM_0                      : inout   std_logic;
          CAM_SPI_1_SS0_Y_0                    : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE : in    std_logic := 'U';
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F    : in    std_logic := 'U'
        );
  end component;

  component m2s010_som_sb_MSS
    port( CORECONFIGP_0_MDDR_APBmslave_PWDATA              : in    std_logic_vector(15 downto 0) := (others => 'U');
          CORECONFIGP_0_MDDR_APBmslave_PADDR               : in    std_logic_vector(10 downto 2) := (others => 'U');
          MAC_MII_RXD_c                                    : in    std_logic_vector(3 downto 0) := (others => 'U');
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA  : in    std_logic_vector(17 downto 0) := (others => 'U');
          Y_net_0                                          : in    std_logic_vector(3 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PRDATA_m                   : in    std_logic_vector(7 downto 0) := (others => 'U');
          CORECONFIGP_0_MDDR_APBmslave_PRDATA              : out   std_logic_vector(15 downto 0);
          MAC_MII_TXD_c                                    : out   std_logic_vector(3 downto 0);
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA  : out   std_logic_vector(16 downto 0);
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR   : out   std_logic_vector(15 downto 2);
          CoreAPB3_0_APBmslave0_PWDATA                     : out   std_logic_vector(7 downto 0);
          m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR           : out   std_logic_vector(15 downto 12);
          CoreAPB3_0_APBmslave0_PADDR                      : out   std_logic_vector(7 downto 0);
          MDDR_ADDR                                        : out   std_logic_vector(15 downto 0);
          MDDR_BA                                          : out   std_logic_vector(2 downto 0);
          MDDR_DM_RDQS                                     : inout   std_logic_vector(1 downto 0);
          MDDR_DQ                                          : inout   std_logic_vector(15 downto 0);
          MDDR_DQS                                         : inout   std_logic_vector(1 downto 0);
          CAM_SPI_1_CLK_Y_0                                : in    std_logic := 'U';
          GPIO_7_Y_0                                       : in    std_logic := 'U';
          GPIO_6_Y_0                                       : in    std_logic := 'U';
          DEBOUNCE_OUT_net_0_0                             : in    std_logic := 'U';
          GPIO_1_in_0                                      : in    std_logic := 'U';
          MDDR_CLK                                         : out   std_logic;
          MDDR_CLK_N                                       : out   std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PWRITE              : in    std_logic := 'U';
          CORECONFIGP_0_MDDR_APBmslave_PSELx               : in    std_logic := 'U';
          CORECONFIGP_0_MDDR_APBmslave_PENABLE             : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz                        : in    std_logic := 'U';
          MAC_MII_TX_CLK_c                                 : in    std_logic := 'U';
          SPI_1_SS0_MX_Y                                   : in    std_logic := 'U';
          SPI_1_DI                                         : in    std_logic := 'U';
          MAC_MII_RX_ER_c                                  : in    std_logic := 'U';
          MAC_MII_RX_DV_c                                  : in    std_logic := 'U';
          MAC_MII_RX_CLK_c                                 : in    std_logic := 'U';
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR : in    std_logic := 'U';
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY  : in    std_logic := 'U';
          MMUART_0_RXD_F2M_c                               : in    std_logic := 'U';
          DEBOUNCE_OUT_2_c                                 : in    std_logic := 'U';
          DEBOUNCE_OUT_1_c                                 : in    std_logic := 'U';
          BIBUF_0_Y                                        : in    std_logic := 'U';
          FAB_CCC_LOCK                                     : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PREADY_i_m_i               : in    std_logic := 'U';
          CommsFPGA_top_0_INT                              : in    std_logic := 'U';
          MAC_MII_CRS_c                                    : in    std_logic := 'U';
          MAC_MII_COL_c                                    : in    std_logic := 'U';
          CORECONFIGP_0_MDDR_APBmslave_PSLVERR             : out   std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PREADY              : out   std_logic;
          MAC_MII_TX_EN_c                                  : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE             : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F                : out   std_logic;
          SPI_1_DO_CAM_c                                   : out   std_logic;
          GPIO_11_M2F_c                                    : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_CLK_M2F                : out   std_logic;
          GPIO_8_M2F_c                                     : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_7_M2F                   : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_7_M2F_OE                : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_6_M2F                   : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_6_M2F_OE                : out   std_logic;
          GPIO_5_M2F_c                                     : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE  : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx   : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE : out   std_logic;
          GPIO_24_M2F_c                                    : out   std_logic;
          MMUART_0_TXD_M2F_c                               : out   std_logic;
          m2s010_som_sb_0_GPIO_28_SW_RESET                 : out   std_logic;
          GPIO_21_M2F_c                                    : out   std_logic;
          GPIO_22_M2F_c                                    : out   std_logic;
          m2s010_som_sb_MSS_0_MAC_MII_MDO                  : out   std_logic;
          m2s010_som_sb_MSS_0_MAC_MII_MDO_EN               : out   std_logic;
          MAC_MII_MDC_c                                    : out   std_logic;
          GPIO_1_M2F                                       : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_1_M2F_OE                : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F          : out   std_logic;
          CoreAPB3_0_APBmslave0_PWRITE                     : out   std_logic;
          m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx           : out   std_logic;
          CoreAPB3_0_APBmslave0_PENABLE                    : out   std_logic;
          GPIO_0_BI                                        : inout   std_logic;
          GPIO_3_BI                                        : inout   std_logic;
          GPIO_4_BI                                        : inout   std_logic;
          GPIO_12_BI                                       : inout   std_logic;
          GPIO_14_BI                                       : inout   std_logic;
          GPIO_15_BI                                       : inout   std_logic;
          GPIO_16_BI                                       : inout   std_logic;
          GPIO_17_BI                                       : inout   std_logic;
          GPIO_18_BI                                       : inout   std_logic;
          GPIO_20_OUT                                      : out   std_logic;
          GPIO_25_BI                                       : inout   std_logic;
          GPIO_26_BI                                       : inout   std_logic;
          GPIO_31_BI                                       : inout   std_logic;
          I2C_1_SCL                                        : inout   std_logic;
          I2C_1_SDA                                        : inout   std_logic;
          MDDR_CAS_N                                       : out   std_logic;
          MDDR_CKE                                         : out   std_logic;
          MDDR_CS_N                                        : out   std_logic;
          MDDR_DQS_TMATCH_0_IN                             : in    std_logic := 'U';
          MDDR_DQS_TMATCH_0_OUT                            : out   std_logic;
          MDDR_ODT                                         : out   std_logic;
          MDDR_RAS_N                                       : out   std_logic;
          MDDR_RESET_N                                     : out   std_logic;
          MDDR_WE_N                                        : out   std_logic;
          MMUART_1_RXD                                     : in    std_logic := 'U';
          MMUART_1_TXD                                     : out   std_logic;
          SPI_0_CLK                                        : inout   std_logic;
          SPI_0_DI                                         : in    std_logic := 'U';
          SPI_0_DO                                         : out   std_logic;
          SPI_0_SS0                                        : inout   std_logic;
          SPI_0_SS1                                        : out   std_logic;
          CORECONFIGP_0_APB_S_PCLK_i                       : out   std_logic;
          CORECONFIGP_0_APB_S_PRESET_N                     : out   std_logic;
          CORECONFIGP_0_APB_S_PCLK                         : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CoreResetP
    port( CORECONFIGP_0_CONFIG2_DONE              : in    std_logic := 'U';
          CORECONFIGP_0_CONFIG1_DONE              : in    std_logic := 'U';
          CORECONFIGP_0_APB_S_PRESET_N            : in    std_logic := 'U';
          m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F : in    std_logic := 'U';
          m2s010_som_sb_0_POWER_ON_RESET_N        : in    std_logic := 'U';
          INIT_DONE                               : out   std_logic;
          FABOSC_0_RCOSC_25_50MHZ_O2F             : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz               : in    std_logic := 'U'
        );
  end component;

  component SYSRESET
    port( POWER_ON_RESET_N : out   std_logic;
          DEVRST_N         : in    std_logic := 'U'
        );
  end component;

  component BIBUF
    generic (IOSTD:string := "");

    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component OUTBUF
    generic (IOSTD:string := "");

    port( D   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component m2s010_som_sb_GPIO_6_IO
    port( GPIO_6_PAD_0                      : inout   std_logic;
          GPIO_6_Y_0                        : out   std_logic;
          m2s010_som_sb_MSS_0_GPIO_6_M2F_OE : in    std_logic := 'U';
          m2s010_som_sb_MSS_0_GPIO_6_M2F    : in    std_logic := 'U'
        );
  end component;

  component CoreConfigP
    port( CORECONFIGP_0_MDDR_APBmslave_PRDATA              : in    std_logic_vector(15 downto 0) := (others => 'U');
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR   : in    std_logic_vector(15 downto 2) := (others => 'U');
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA  : out   std_logic_vector(17 downto 0);
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA  : in    std_logic_vector(16 downto 0) := (others => 'U');
          CORECONFIGP_0_MDDR_APBmslave_PADDR               : out   std_logic_vector(10 downto 2);
          CORECONFIGP_0_MDDR_APBmslave_PWDATA              : out   std_logic_vector(15 downto 0);
          CORECONFIGP_0_MDDR_APBmslave_PSLVERR             : in    std_logic := 'U';
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx   : in    std_logic := 'U';
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE : in    std_logic := 'U';
          CORECONFIGP_0_MDDR_APBmslave_PREADY              : in    std_logic := 'U';
          CORECONFIGP_0_MDDR_APBmslave_PSELx               : out   std_logic;
          CORECONFIGP_0_MDDR_APBmslave_PENABLE             : out   std_logic;
          INIT_DONE                                        : in    std_logic := 'U';
          CORECONFIGP_0_APB_S_PCLK_i                       : in    std_logic := 'U';
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE  : in    std_logic := 'U';
          CORECONFIGP_0_MDDR_APBmslave_PWRITE              : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR : out   std_logic;
          m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY  : out   std_logic;
          CORECONFIGP_0_CONFIG2_DONE                       : out   std_logic;
          CORECONFIGP_0_CONFIG1_DONE                       : out   std_logic;
          CORECONFIGP_0_APB_S_PCLK                         : in    std_logic := 'U';
          CORECONFIGP_0_APB_S_PRESET_N                     : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component m2s010_som_sb_CCC_0_FCCC
    port( m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC : in    std_logic := 'U';
          FAB_CCC_LOCK                              : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz                 : out   std_logic
        );
  end component;

  component m2s010_som_sb_OTH_SPI_1_SS0_IO
    port( SPI_1_SS0_OTH_0                      : inout   std_logic;
          OTH_SPI_1_SS0_Y_0                    : out   std_logic;
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE : in    std_logic := 'U';
          m2s010_som_sb_MSS_0_SPI_1_SS0_M2F    : in    std_logic := 'U'
        );
  end component;

  component m2s010_som_sb_FABOSC_0_OSC
    port( XTL                                       : in    std_logic := 'U';
          m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC : out   std_logic;
          FABOSC_0_RCOSC_25_50MHZ_O2F               : out   std_logic
        );
  end component;

    signal BIBUF_0_Y, m2s010_som_sb_MSS_0_MAC_MII_MDO, 
        m2s010_som_sb_MSS_0_MAC_MII_MDO_EN, 
        \m2s010_som_sb_0_POWER_ON_RESET_N\, SPI_1_SS0_MX_Y, 
        \OTH_SPI_1_SS0_Y[0]\, \CAM_SPI_1_SS0_Y[0]\, SPI_1_DI, 
        \CAM_SPI_1_CLK_Y[0]\, 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE, 
        m2s010_som_sb_MSS_0_SPI_1_CLK_M2F, 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F, FAB_CCC_LOCK, 
        \m2s010_som_sb_0_CCC_71MHz\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[0]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[1]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[2]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[3]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[4]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[5]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[6]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[7]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[8]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[9]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[10]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[11]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[12]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[13]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[14]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[15]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[2]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[3]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[4]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[5]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[6]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[7]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[8]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[9]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[10]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[12]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[13]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[15]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[0]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[1]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[2]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[3]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[4]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[5]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[6]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[7]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[8]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[9]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[10]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[11]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[12]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[13]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[14]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[15]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[16]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[17]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[0]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[1]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[2]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[3]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[4]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[5]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[6]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[7]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[8]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[9]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[10]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[11]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[12]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[13]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[14]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[15]\, 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[16]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[2]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[3]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[4]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[5]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[6]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[7]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[8]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[9]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[10]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[0]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[1]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[2]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[3]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[4]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[5]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[6]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[7]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[8]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[9]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[10]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[11]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[12]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[13]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[14]\, 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[15]\, 
        CORECONFIGP_0_MDDR_APBmslave_PSLVERR, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE, 
        CORECONFIGP_0_MDDR_APBmslave_PREADY, 
        CORECONFIGP_0_MDDR_APBmslave_PSELx, 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE, INIT_DONE, 
        CORECONFIGP_0_APB_S_PCLK_i, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE, 
        CORECONFIGP_0_MDDR_APBmslave_PWRITE, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY, 
        CORECONFIGP_0_CONFIG2_DONE, CORECONFIGP_0_CONFIG1_DONE, 
        CORECONFIGP_0_APB_S_PCLK, CORECONFIGP_0_APB_S_PRESET_N, 
        m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        FABOSC_0_RCOSC_25_50MHZ_O2F, \GPIO_1_in[0]\, 
        m2s010_som_sb_MSS_0_GPIO_1_M2F_OE, GPIO_1_M2F, 
        \GPIO_6_Y[0]\, m2s010_som_sb_MSS_0_GPIO_6_M2F_OE, 
        m2s010_som_sb_MSS_0_GPIO_6_M2F, \GPIO_7_Y[0]\, 
        m2s010_som_sb_MSS_0_GPIO_7_M2F_OE, 
        m2s010_som_sb_MSS_0_GPIO_7_M2F, GND_net_1, VCC_net_1
         : std_logic;
    signal nc2, nc4, nc3, nc1 : std_logic;

    for all : m2s010_som_sb_GPIO_1_IO
	Use entity work.m2s010_som_sb_GPIO_1_IO(DEF_ARCH);
    for all : m2s010_som_sb_CAM_SPI_1_CLK_IO
	Use entity work.m2s010_som_sb_CAM_SPI_1_CLK_IO(DEF_ARCH);
    for all : m2s010_som_sb_GPIO_7_IO
	Use entity work.m2s010_som_sb_GPIO_7_IO(DEF_ARCH);
    for all : m2s010_som_sb_CAM_SPI_1_SS0_IO
	Use entity work.m2s010_som_sb_CAM_SPI_1_SS0_IO(DEF_ARCH);
    for all : m2s010_som_sb_MSS
	Use entity work.m2s010_som_sb_MSS(DEF_ARCH);
    for all : CoreResetP
	Use entity work.CoreResetP(DEF_ARCH);
    for all : m2s010_som_sb_GPIO_6_IO
	Use entity work.m2s010_som_sb_GPIO_6_IO(DEF_ARCH);
    for all : CoreConfigP
	Use entity work.CoreConfigP(DEF_ARCH);
    for all : m2s010_som_sb_CCC_0_FCCC
	Use entity work.m2s010_som_sb_CCC_0_FCCC(DEF_ARCH);
    for all : m2s010_som_sb_OTH_SPI_1_SS0_IO
	Use entity work.m2s010_som_sb_OTH_SPI_1_SS0_IO(DEF_ARCH);
    for all : m2s010_som_sb_FABOSC_0_OSC
	Use entity work.m2s010_som_sb_FABOSC_0_OSC(DEF_ARCH);
begin 

    m2s010_som_sb_0_CCC_71MHz <= \m2s010_som_sb_0_CCC_71MHz\;
    m2s010_som_sb_0_POWER_ON_RESET_N <= 
        \m2s010_som_sb_0_POWER_ON_RESET_N\;

    GPIO_1 : m2s010_som_sb_GPIO_1_IO
      port map(GPIO_1_BI_0 => GPIO_1_BI_0, GPIO_1_in_0 => 
        \GPIO_1_in[0]\, m2s010_som_sb_MSS_0_GPIO_1_M2F_OE => 
        m2s010_som_sb_MSS_0_GPIO_1_M2F_OE, GPIO_1_M2F => 
        GPIO_1_M2F);
    
    CAM_SPI_1_CLK : m2s010_som_sb_CAM_SPI_1_CLK_IO
      port map(CAM_SPI_1_CLK_Y_0 => \CAM_SPI_1_CLK_Y[0]\, 
        SPI_1_CLK_0 => SPI_1_CLK_0, 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE, 
        m2s010_som_sb_MSS_0_SPI_1_CLK_M2F => 
        m2s010_som_sb_MSS_0_SPI_1_CLK_M2F);
    
    GPIO_7 : m2s010_som_sb_GPIO_7_IO
      port map(GPIO_7_PADI_0 => GPIO_7_PADI_0, GPIO_7_Y_0 => 
        \GPIO_7_Y[0]\, m2s010_som_sb_MSS_0_GPIO_7_M2F_OE => 
        m2s010_som_sb_MSS_0_GPIO_7_M2F_OE, 
        m2s010_som_sb_MSS_0_GPIO_7_M2F => 
        m2s010_som_sb_MSS_0_GPIO_7_M2F);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    CAM_SPI_1_SS0 : m2s010_som_sb_CAM_SPI_1_SS0_IO
      port map(SPI_1_SS0_CAM_0 => SPI_1_SS0_CAM_0, 
        CAM_SPI_1_SS0_Y_0 => \CAM_SPI_1_SS0_Y[0]\, 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE, 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F);
    
    m2s010_som_sb_MSS_0 : m2s010_som_sb_MSS
      port map(CORECONFIGP_0_MDDR_APBmslave_PWDATA(15) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[15]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(14) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[14]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(13) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[13]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(12) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[12]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(11) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[11]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(10) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[10]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(9) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[9]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(8) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[8]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(7) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[7]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(6) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[6]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(5) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[5]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(4) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[4]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(3) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[3]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(2) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[2]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(1) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[1]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(0) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[0]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(10) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[10]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(9) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[9]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(8) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[8]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(7) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[7]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(6) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[6]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(5) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[5]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(4) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[4]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(3) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[3]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(2) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[2]\, MAC_MII_RXD_c(3)
         => MAC_MII_RXD_c(3), MAC_MII_RXD_c(2) => 
        MAC_MII_RXD_c(2), MAC_MII_RXD_c(1) => MAC_MII_RXD_c(1), 
        MAC_MII_RXD_c(0) => MAC_MII_RXD_c(0), 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(17) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[17]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(16) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[16]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(15) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[15]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(14) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[14]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(13) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[13]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(12) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[12]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(11) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[11]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(10) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[10]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(9) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[9]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(8) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[8]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(7) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[7]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(6) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[6]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(5) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[5]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(4) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[4]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(3) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[3]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(2) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[2]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(1) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[1]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(0) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[0]\, 
        Y_net_0(3) => Y_net_0(3), Y_net_0(2) => Y_net_0(2), 
        Y_net_0(1) => Y_net_0(1), Y_net_0(0) => Y_net_0(0), 
        CoreAPB3_0_APBmslave0_PRDATA_m(7) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(7), 
        CoreAPB3_0_APBmslave0_PRDATA_m(6) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(6), 
        CoreAPB3_0_APBmslave0_PRDATA_m(5) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(5), 
        CoreAPB3_0_APBmslave0_PRDATA_m(4) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(4), 
        CoreAPB3_0_APBmslave0_PRDATA_m(3) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(3), 
        CoreAPB3_0_APBmslave0_PRDATA_m(2) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(2), 
        CoreAPB3_0_APBmslave0_PRDATA_m(1) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(1), 
        CoreAPB3_0_APBmslave0_PRDATA_m(0) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(0), 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(15) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[15]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(14) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[14]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(13) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[13]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(12) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[12]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(11) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[11]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(10) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[10]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(9) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[9]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(8) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[8]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(7) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[7]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(6) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[6]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(5) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[5]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(4) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[4]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(3) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[3]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(2) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[2]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(1) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[1]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(0) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[0]\, 
        MAC_MII_TXD_c(3) => MAC_MII_TXD_c(3), MAC_MII_TXD_c(2)
         => MAC_MII_TXD_c(2), MAC_MII_TXD_c(1) => 
        MAC_MII_TXD_c(1), MAC_MII_TXD_c(0) => MAC_MII_TXD_c(0), 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(16) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[16]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(15) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[15]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(14) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[14]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(13) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[13]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(12) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[12]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(11) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[11]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(10) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[10]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(9) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[9]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(8) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[8]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(7) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[7]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(6) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[6]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(5) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[5]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(4) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[4]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(3) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[3]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(2) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[2]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(1) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[1]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(0) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[0]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(15) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[15]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(14) => nc2, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(13) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[13]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(12) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[12]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(11) => nc4, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(10) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[10]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(9) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[9]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(8) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[8]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(7) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[7]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(6) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[6]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(5) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[5]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[4]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[3]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[2]\, 
        CoreAPB3_0_APBmslave0_PWDATA(7) => 
        CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(15) => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(15), 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(14) => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(14), 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(13) => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(13), 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(12) => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(12), 
        CoreAPB3_0_APBmslave0_PADDR(7) => 
        CoreAPB3_0_APBmslave0_PADDR(7), 
        CoreAPB3_0_APBmslave0_PADDR(6) => 
        CoreAPB3_0_APBmslave0_PADDR(6), 
        CoreAPB3_0_APBmslave0_PADDR(5) => 
        CoreAPB3_0_APBmslave0_PADDR(5), 
        CoreAPB3_0_APBmslave0_PADDR(4) => 
        CoreAPB3_0_APBmslave0_PADDR(4), 
        CoreAPB3_0_APBmslave0_PADDR(3) => 
        CoreAPB3_0_APBmslave0_PADDR(3), 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        CoreAPB3_0_APBmslave0_PADDR(2), 
        CoreAPB3_0_APBmslave0_PADDR(1) => 
        CoreAPB3_0_APBmslave0_PADDR(1), 
        CoreAPB3_0_APBmslave0_PADDR(0) => 
        CoreAPB3_0_APBmslave0_PADDR(0), MDDR_ADDR(15) => 
        MDDR_ADDR(15), MDDR_ADDR(14) => MDDR_ADDR(14), 
        MDDR_ADDR(13) => MDDR_ADDR(13), MDDR_ADDR(12) => 
        MDDR_ADDR(12), MDDR_ADDR(11) => MDDR_ADDR(11), 
        MDDR_ADDR(10) => MDDR_ADDR(10), MDDR_ADDR(9) => 
        MDDR_ADDR(9), MDDR_ADDR(8) => MDDR_ADDR(8), MDDR_ADDR(7)
         => MDDR_ADDR(7), MDDR_ADDR(6) => MDDR_ADDR(6), 
        MDDR_ADDR(5) => MDDR_ADDR(5), MDDR_ADDR(4) => 
        MDDR_ADDR(4), MDDR_ADDR(3) => MDDR_ADDR(3), MDDR_ADDR(2)
         => MDDR_ADDR(2), MDDR_ADDR(1) => MDDR_ADDR(1), 
        MDDR_ADDR(0) => MDDR_ADDR(0), MDDR_BA(2) => MDDR_BA(2), 
        MDDR_BA(1) => MDDR_BA(1), MDDR_BA(0) => MDDR_BA(0), 
        MDDR_DM_RDQS(1) => MDDR_DM_RDQS(1), MDDR_DM_RDQS(0) => 
        MDDR_DM_RDQS(0), MDDR_DQ(15) => MDDR_DQ(15), MDDR_DQ(14)
         => MDDR_DQ(14), MDDR_DQ(13) => MDDR_DQ(13), MDDR_DQ(12)
         => MDDR_DQ(12), MDDR_DQ(11) => MDDR_DQ(11), MDDR_DQ(10)
         => MDDR_DQ(10), MDDR_DQ(9) => MDDR_DQ(9), MDDR_DQ(8) => 
        MDDR_DQ(8), MDDR_DQ(7) => MDDR_DQ(7), MDDR_DQ(6) => 
        MDDR_DQ(6), MDDR_DQ(5) => MDDR_DQ(5), MDDR_DQ(4) => 
        MDDR_DQ(4), MDDR_DQ(3) => MDDR_DQ(3), MDDR_DQ(2) => 
        MDDR_DQ(2), MDDR_DQ(1) => MDDR_DQ(1), MDDR_DQ(0) => 
        MDDR_DQ(0), MDDR_DQS(1) => MDDR_DQS(1), MDDR_DQS(0) => 
        MDDR_DQS(0), CAM_SPI_1_CLK_Y_0 => \CAM_SPI_1_CLK_Y[0]\, 
        GPIO_7_Y_0 => \GPIO_7_Y[0]\, GPIO_6_Y_0 => \GPIO_6_Y[0]\, 
        DEBOUNCE_OUT_net_0_0 => DEBOUNCE_OUT_net_0_0, GPIO_1_in_0
         => \GPIO_1_in[0]\, MDDR_CLK => MDDR_CLK, MDDR_CLK_N => 
        MDDR_CLK_N, CORECONFIGP_0_MDDR_APBmslave_PWRITE => 
        CORECONFIGP_0_MDDR_APBmslave_PWRITE, 
        CORECONFIGP_0_MDDR_APBmslave_PSELx => 
        CORECONFIGP_0_MDDR_APBmslave_PSELx, 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE => 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE, 
        m2s010_som_sb_0_CCC_71MHz => \m2s010_som_sb_0_CCC_71MHz\, 
        MAC_MII_TX_CLK_c => MAC_MII_TX_CLK_c, SPI_1_SS0_MX_Y => 
        SPI_1_SS0_MX_Y, SPI_1_DI => SPI_1_DI, MAC_MII_RX_ER_c => 
        MAC_MII_RX_ER_c, MAC_MII_RX_DV_c => MAC_MII_RX_DV_c, 
        MAC_MII_RX_CLK_c => MAC_MII_RX_CLK_c, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY, 
        MMUART_0_RXD_F2M_c => MMUART_0_RXD_F2M_c, 
        DEBOUNCE_OUT_2_c => DEBOUNCE_OUT_2_c, DEBOUNCE_OUT_1_c
         => DEBOUNCE_OUT_1_c, BIBUF_0_Y => BIBUF_0_Y, 
        FAB_CCC_LOCK => FAB_CCC_LOCK, 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i => 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i, CommsFPGA_top_0_INT
         => CommsFPGA_top_0_INT, MAC_MII_CRS_c => MAC_MII_CRS_c, 
        MAC_MII_COL_c => MAC_MII_COL_c, 
        CORECONFIGP_0_MDDR_APBmslave_PSLVERR => 
        CORECONFIGP_0_MDDR_APBmslave_PSLVERR, 
        CORECONFIGP_0_MDDR_APBmslave_PREADY => 
        CORECONFIGP_0_MDDR_APBmslave_PREADY, MAC_MII_TX_EN_c => 
        MAC_MII_TX_EN_c, m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE, 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F, SPI_1_DO_CAM_c => 
        SPI_1_DO_CAM_c, GPIO_11_M2F_c => GPIO_11_M2F_c, 
        m2s010_som_sb_MSS_0_SPI_1_CLK_M2F => 
        m2s010_som_sb_MSS_0_SPI_1_CLK_M2F, GPIO_8_M2F_c => 
        GPIO_8_M2F_c, m2s010_som_sb_MSS_0_GPIO_7_M2F => 
        m2s010_som_sb_MSS_0_GPIO_7_M2F, 
        m2s010_som_sb_MSS_0_GPIO_7_M2F_OE => 
        m2s010_som_sb_MSS_0_GPIO_7_M2F_OE, 
        m2s010_som_sb_MSS_0_GPIO_6_M2F => 
        m2s010_som_sb_MSS_0_GPIO_6_M2F, 
        m2s010_som_sb_MSS_0_GPIO_6_M2F_OE => 
        m2s010_som_sb_MSS_0_GPIO_6_M2F_OE, GPIO_5_M2F_c => 
        GPIO_5_M2F_c, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE, 
        GPIO_24_M2F_c => GPIO_24_M2F_c, MMUART_0_TXD_M2F_c => 
        MMUART_0_TXD_M2F_c, m2s010_som_sb_0_GPIO_28_SW_RESET => 
        m2s010_som_sb_0_GPIO_28_SW_RESET, GPIO_21_M2F_c => 
        GPIO_21_M2F_c, GPIO_22_M2F_c => GPIO_22_M2F_c, 
        m2s010_som_sb_MSS_0_MAC_MII_MDO => 
        m2s010_som_sb_MSS_0_MAC_MII_MDO, 
        m2s010_som_sb_MSS_0_MAC_MII_MDO_EN => 
        m2s010_som_sb_MSS_0_MAC_MII_MDO_EN, MAC_MII_MDC_c => 
        MAC_MII_MDC_c, GPIO_1_M2F => GPIO_1_M2F, 
        m2s010_som_sb_MSS_0_GPIO_1_M2F_OE => 
        m2s010_som_sb_MSS_0_GPIO_1_M2F_OE, 
        m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F => 
        m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        CoreAPB3_0_APBmslave0_PWRITE => 
        CoreAPB3_0_APBmslave0_PWRITE, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx, 
        CoreAPB3_0_APBmslave0_PENABLE => 
        CoreAPB3_0_APBmslave0_PENABLE, GPIO_0_BI => GPIO_0_BI, 
        GPIO_3_BI => GPIO_3_BI, GPIO_4_BI => GPIO_4_BI, 
        GPIO_12_BI => GPIO_12_BI, GPIO_14_BI => GPIO_14_BI, 
        GPIO_15_BI => GPIO_15_BI, GPIO_16_BI => GPIO_16_BI, 
        GPIO_17_BI => GPIO_17_BI, GPIO_18_BI => GPIO_18_BI, 
        GPIO_20_OUT => GPIO_20_OUT, GPIO_25_BI => GPIO_25_BI, 
        GPIO_26_BI => GPIO_26_BI, GPIO_31_BI => GPIO_31_BI, 
        I2C_1_SCL => I2C_1_SCL, I2C_1_SDA => I2C_1_SDA, 
        MDDR_CAS_N => MDDR_CAS_N, MDDR_CKE => MDDR_CKE, MDDR_CS_N
         => MDDR_CS_N, MDDR_DQS_TMATCH_0_IN => 
        MDDR_DQS_TMATCH_0_IN, MDDR_DQS_TMATCH_0_OUT => 
        MDDR_DQS_TMATCH_0_OUT, MDDR_ODT => MDDR_ODT, MDDR_RAS_N
         => MDDR_RAS_N, MDDR_RESET_N => MDDR_RESET_N, MDDR_WE_N
         => MDDR_WE_N, MMUART_1_RXD => MMUART_1_RXD, MMUART_1_TXD
         => MMUART_1_TXD, SPI_0_CLK => SPI_0_CLK, SPI_0_DI => 
        SPI_0_DI, SPI_0_DO => SPI_0_DO, SPI_0_SS0 => SPI_0_SS0, 
        SPI_0_SS1 => SPI_0_SS1, CORECONFIGP_0_APB_S_PCLK_i => 
        CORECONFIGP_0_APB_S_PCLK_i, CORECONFIGP_0_APB_S_PRESET_N
         => CORECONFIGP_0_APB_S_PRESET_N, 
        CORECONFIGP_0_APB_S_PCLK => CORECONFIGP_0_APB_S_PCLK);
    
    SPI_1_SS0_MX : MX2
      port map(A => \OTH_SPI_1_SS0_Y[0]\, B => 
        \CAM_SPI_1_SS0_Y[0]\, S => CommsFPGA_top_0_CAMERA_NODE, Y
         => SPI_1_SS0_MX_Y);
    
    CORERESETP_0 : CoreResetP
      port map(CORECONFIGP_0_CONFIG2_DONE => 
        CORECONFIGP_0_CONFIG2_DONE, CORECONFIGP_0_CONFIG1_DONE
         => CORECONFIGP_0_CONFIG1_DONE, 
        CORECONFIGP_0_APB_S_PRESET_N => 
        CORECONFIGP_0_APB_S_PRESET_N, 
        m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F => 
        m2s010_som_sb_MSS_TMP_0_MSS_RESET_N_M2F, 
        m2s010_som_sb_0_POWER_ON_RESET_N => 
        \m2s010_som_sb_0_POWER_ON_RESET_N\, INIT_DONE => 
        INIT_DONE, FABOSC_0_RCOSC_25_50MHZ_O2F => 
        FABOSC_0_RCOSC_25_50MHZ_O2F, m2s010_som_sb_0_CCC_71MHz
         => \m2s010_som_sb_0_CCC_71MHz\);
    
    SYSRESET_POR : SYSRESET
      port map(POWER_ON_RESET_N => 
        \m2s010_som_sb_0_POWER_ON_RESET_N\, DEVRST_N => DEVRST_N);
    
    BIBUF_0 : BIBUF
      port map(PAD => MAC_MII_MDIO, D => 
        m2s010_som_sb_MSS_0_MAC_MII_MDO, E => 
        m2s010_som_sb_MSS_0_MAC_MII_MDO_EN, Y => BIBUF_0_Y);
    
    SPI_1_D0_OUT : OUTBUF
      port map(D => SPI_1_DO_CAM_c, PAD => SPI_1_DO_OTH);
    
    GPIO_6 : m2s010_som_sb_GPIO_6_IO
      port map(GPIO_6_PAD_0 => GPIO_6_PAD_0, GPIO_6_Y_0 => 
        \GPIO_6_Y[0]\, m2s010_som_sb_MSS_0_GPIO_6_M2F_OE => 
        m2s010_som_sb_MSS_0_GPIO_6_M2F_OE, 
        m2s010_som_sb_MSS_0_GPIO_6_M2F => 
        m2s010_som_sb_MSS_0_GPIO_6_M2F);
    
    CORECONFIGP_0 : CoreConfigP
      port map(CORECONFIGP_0_MDDR_APBmslave_PRDATA(15) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[15]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(14) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[14]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(13) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[13]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(12) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[12]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(11) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[11]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(10) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[10]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(9) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[9]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(8) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[8]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(7) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[7]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(6) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[6]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(5) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[5]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(4) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[4]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(3) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[3]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(2) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[2]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(1) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[1]\, 
        CORECONFIGP_0_MDDR_APBmslave_PRDATA(0) => 
        \CORECONFIGP_0_MDDR_APBmslave_PRDATA[0]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(15) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[15]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(14) => nc3, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(13) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[13]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(12) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[12]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(11) => nc1, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(10) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[10]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(9) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[9]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(8) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[8]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(7) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[7]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(6) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[6]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(5) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[5]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(4) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[4]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(3) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[3]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR(2) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PADDR[2]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(17) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[17]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(16) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[16]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(15) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[15]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(14) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[14]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(13) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[13]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(12) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[12]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(11) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[11]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(10) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[10]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(9) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[9]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(8) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[8]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(7) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[7]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(6) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[6]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(5) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[5]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(4) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[4]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(3) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[3]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(2) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[2]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(1) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[1]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA(0) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PRDATA[0]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(16) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[16]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(15) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[15]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(14) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[14]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(13) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[13]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(12) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[12]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(11) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[11]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(10) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[10]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(9) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[9]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(8) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[8]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(7) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[7]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(6) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[6]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(5) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[5]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(4) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[4]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(3) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[3]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(2) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[2]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(1) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[1]\, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA(0) => 
        \m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWDATA[0]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(10) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[10]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(9) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[9]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(8) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[8]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(7) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[7]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(6) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[6]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(5) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[5]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(4) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[4]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(3) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[3]\, 
        CORECONFIGP_0_MDDR_APBmslave_PADDR(2) => 
        \CORECONFIGP_0_MDDR_APBmslave_PADDR[2]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(15) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[15]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(14) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[14]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(13) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[13]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(12) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[12]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(11) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[11]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(10) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[10]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(9) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[9]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(8) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[8]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(7) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[7]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(6) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[6]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(5) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[5]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(4) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[4]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(3) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[3]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(2) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[2]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(1) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[1]\, 
        CORECONFIGP_0_MDDR_APBmslave_PWDATA(0) => 
        \CORECONFIGP_0_MDDR_APBmslave_PWDATA[0]\, 
        CORECONFIGP_0_MDDR_APBmslave_PSLVERR => 
        CORECONFIGP_0_MDDR_APBmslave_PSLVERR, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSELx, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PENABLE, 
        CORECONFIGP_0_MDDR_APBmslave_PREADY => 
        CORECONFIGP_0_MDDR_APBmslave_PREADY, 
        CORECONFIGP_0_MDDR_APBmslave_PSELx => 
        CORECONFIGP_0_MDDR_APBmslave_PSELx, 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE => 
        CORECONFIGP_0_MDDR_APBmslave_PENABLE, INIT_DONE => 
        INIT_DONE, CORECONFIGP_0_APB_S_PCLK_i => 
        CORECONFIGP_0_APB_S_PCLK_i, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PWRITE, 
        CORECONFIGP_0_MDDR_APBmslave_PWRITE => 
        CORECONFIGP_0_MDDR_APBmslave_PWRITE, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PSLVERR, 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY => 
        m2s010_som_sb_MSS_TMP_0_FIC_2_APB_MASTER_PREADY, 
        CORECONFIGP_0_CONFIG2_DONE => CORECONFIGP_0_CONFIG2_DONE, 
        CORECONFIGP_0_CONFIG1_DONE => CORECONFIGP_0_CONFIG1_DONE, 
        CORECONFIGP_0_APB_S_PCLK => CORECONFIGP_0_APB_S_PCLK, 
        CORECONFIGP_0_APB_S_PRESET_N => 
        CORECONFIGP_0_APB_S_PRESET_N);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    CCC_0 : m2s010_som_sb_CCC_0_FCCC
      port map(m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC => 
        m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC, FAB_CCC_LOCK
         => FAB_CCC_LOCK, m2s010_som_sb_0_CCC_71MHz => 
        \m2s010_som_sb_0_CCC_71MHz\);
    
    SPI_1_DI_MX : MX2
      port map(A => SPI_1_DI_OTH_c, B => SPI_1_DI_CAM_c, S => 
        CommsFPGA_top_0_CAMERA_NODE, Y => SPI_1_DI);
    
    OTH_SPI_1_SS0 : m2s010_som_sb_OTH_SPI_1_SS0_IO
      port map(SPI_1_SS0_OTH_0 => SPI_1_SS0_OTH_0, 
        OTH_SPI_1_SS0_Y_0 => \OTH_SPI_1_SS0_Y[0]\, 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F_OE, 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F => 
        m2s010_som_sb_MSS_0_SPI_1_SS0_M2F);
    
    FABOSC_0 : m2s010_som_sb_FABOSC_0_OSC
      port map(XTL => XTL, 
        m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC => 
        m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC, 
        FABOSC_0_RCOSC_25_50MHZ_O2F => 
        FABOSC_0_RCOSC_25_50MHZ_O2F);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity Debounce_1 is

    port( DEBOUNCE_IN_c_0  : in    std_logic;
          RESET            : in    std_logic;
          DEBOUNCE_OUT_2_c : out   std_logic;
          RESET_set        : in    std_logic;
          BIT_CLK          : in    std_logic
        );

end Debounce_1;

architecture DEF_ARCH of Debounce_1 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \debounce_cntr[1]_net_1\, VCC_net_1, 
        un2_debounce_in_i, un3_debounce_cntr_1_cry_1_S_1, 
        GND_net_1, \debounce_cntr[2]_net_1\, 
        un3_debounce_cntr_1_cry_2_S_1, \debounce_cntr[3]_net_1\, 
        un3_debounce_cntr_1_cry_3_S_1, \debounce_cntrrs[4]\, 
        un3_debounce_in_rs_1, \debounce_cntr[4]\, 
        un3_debounce_in_i, un3_debounce_cntr_1_cry_4_S_1, 
        \debounce_cntrrs[6]\, \debounce_cntr[6]\, 
        un3_debounce_cntr_1_cry_6_S_1, \debounce_cntr[5]\, 
        un3_debounce_cntr_1_cry_5_S_1, \debounce_cntr[7]\, 
        un3_debounce_cntr_1_cry_7_S_1, \debounce_cntrrs[8]\, 
        \debounce_cntr[8]_net_1\, un3_debounce_cntr_1_cry_8_S_1, 
        \debounce_cntrrs[9]\, \debounce_cntr[9]_net_1\, 
        un3_debounce_cntr_1_cry_9_S_1, \debounce_cntr[10]_net_1\, 
        un3_debounce_cntr_1_cry_10_S_1, \debounce_cntr[11]_net_1\, 
        un3_debounce_cntr_1_cry_11_S_1, \debounce_cntr[12]_net_1\, 
        un3_debounce_cntr_1_cry_12_S_1, \debounce_cntr[13]_net_1\, 
        un3_debounce_cntr_1_cry_13_S_1, \debounce_cntrrs[14]\, 
        \debounce_cntr[14]_net_1\, un3_debounce_cntr_1_cry_14_S_1, 
        \debounce_cntrrs[15]\, \debounce_cntr[15]_net_1\, 
        un3_debounce_cntr_1_s_15_S_1, \debounce_cntr[0]_net_1\, 
        \debounce_cntr_4[0]_net_1\, DEBOUNCE_OUT_2_crs, 
        un1_debounce_cntr, un3_debounce_cntr_1_s_1_919_FCO, 
        \un3_debounce_cntr_1_cry_1\, \un3_debounce_cntr_1_cry_2\, 
        \un3_debounce_cntr_1_cry_3\, \un3_debounce_cntr_1_cry_4\, 
        \un3_debounce_cntr_1_cry_5\, \un3_debounce_cntr_1_cry_6\, 
        \un3_debounce_cntr_1_cry_7\, \un3_debounce_cntr_1_cry_8\, 
        \un3_debounce_cntr_1_cry_9\, \un3_debounce_cntr_1_cry_10\, 
        \un3_debounce_cntr_1_cry_11\, 
        \un3_debounce_cntr_1_cry_12\, 
        \un3_debounce_cntr_1_cry_13\, 
        \un3_debounce_cntr_1_cry_14\, un1_debounce_cntr_11, 
        un1_debounce_cntr_10, un1_debounce_cntr_9, 
        un1_debounce_cntr_8 : std_logic;

begin 


    \debounce_cntr_0_0[0]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_5_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[5]\);
    
    un3_debounce_cntr_1_cry_9 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[9]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_8\, S => 
        un3_debounce_cntr_1_cry_9_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_9\);
    
    \debounce_cntr[12]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_12_S_1, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => un2_debounce_in_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[12]_net_1\);
    
    \debounce_cntr_RNICP4M[9]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \debounce_cntrrs[9]\, B => 
        un3_debounce_in_rs_1, C => RESET_set, Y => 
        \debounce_cntr[9]_net_1\);
    
    un3_debounce_cntr_1_s_1_919 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[0]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => 
        OPEN, Y => OPEN, FCO => un3_debounce_cntr_1_s_1_919_FCO);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_8\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \debounce_cntr[2]_net_1\, B => 
        \debounce_cntr[1]_net_1\, C => \debounce_cntr[15]_net_1\, 
        D => \debounce_cntr[14]_net_1\, Y => un1_debounce_cntr_8);
    
    \DEBOUNCE_PROC.un3_debounce_in_rs\ : SLE
      port map(D => VCC_net_1, CLK => RESET, EN => VCC_net_1, ALn
         => un3_debounce_in_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => VCC_net_1, Q => 
        un3_debounce_in_rs_1);
    
    \debounce_cntr[15]\ : SLE
      port map(D => un3_debounce_cntr_1_s_15_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[15]\);
    
    un3_debounce_cntr_1_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_4\, S => 
        un3_debounce_cntr_1_cry_5_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_5\);
    
    un3_debounce_cntr_1_cry_2 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[2]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_1\, S => 
        un3_debounce_cntr_1_cry_2_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_2\);
    
    \debounce_cntr[3]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_3_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[3]_net_1\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_9\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \debounce_cntr[9]_net_1\, B => 
        \debounce_cntr[8]_net_1\, C => \debounce_cntr[6]\, D => 
        \debounce_cntr[4]\, Y => un1_debounce_cntr_9);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_10\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \debounce_cntr[13]_net_1\, B => 
        \debounce_cntr[12]_net_1\, C => \debounce_cntr[11]_net_1\, 
        D => \debounce_cntr[10]_net_1\, Y => un1_debounce_cntr_10);
    
    \debounce_cntr_0_RNIIE8T[0]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \debounce_cntrrs[4]\, B => 
        un3_debounce_in_rs_1, C => RESET_set, Y => 
        \debounce_cntr[4]\);
    
    debounce_out : SLE
      port map(D => un1_debounce_cntr, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => un3_debounce_in_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => DEBOUNCE_OUT_2_crs);
    
    \debounce_cntr[10]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_10_S_1, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => un2_debounce_in_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[10]_net_1\);
    
    \debounce_cntr_RNIOP221[14]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \debounce_cntrrs[14]\, B => 
        un3_debounce_in_rs_1, C => RESET_set, Y => 
        \debounce_cntr[14]_net_1\);
    
    un3_debounce_cntr_1_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_3\, S => 
        un3_debounce_cntr_1_cry_4_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_4\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \debounce_cntr[13]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_13_S_1, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => un2_debounce_in_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[13]_net_1\);
    
    un3_debounce_cntr_1_cry_14 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[14]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_13\, S => 
        un3_debounce_cntr_1_cry_14_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_14\);
    
    \debounce_cntr_0_0[1]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_7_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[7]\);
    
    un3_debounce_cntr_1_cry_13 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[13]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_12\, S => 
        un3_debounce_cntr_1_cry_13_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_13\);
    
    \debounce_cntr[9]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_9_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[9]\);
    
    un3_debounce_cntr_1_cry_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_6\, S => 
        un3_debounce_cntr_1_cry_7_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_7\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \DEBOUNCE_PROC.un2_debounce_in\ : CFG2
      generic map(INIT => x"2")

      port map(A => DEBOUNCE_IN_c_0, B => RESET, Y => 
        un2_debounce_in_i);
    
    \debounce_cntr[1]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_1_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[1]_net_1\);
    
    debounce_out_RNISK1S : CFG3
      generic map(INIT => x"F8")

      port map(A => un3_debounce_in_rs_1, B => RESET_set, C => 
        DEBOUNCE_OUT_2_crs, Y => DEBOUNCE_OUT_2_c);
    
    \debounce_cntr_0[0]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_4_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[4]\);
    
    \debounce_cntr[14]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_14_S_1, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => un3_debounce_in_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[14]\);
    
    un3_debounce_cntr_1_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_5\, S => 
        un3_debounce_cntr_1_cry_6_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_6\);
    
    \debounce_cntr_0_RNIJF8T[1]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \debounce_cntrrs[6]\, B => 
        un3_debounce_in_rs_1, C => RESET_set, Y => 
        \debounce_cntr[6]\);
    
    un3_debounce_cntr_1_cry_11 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[11]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_10\, S => 
        un3_debounce_cntr_1_cry_11_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_11\);
    
    \debounce_cntr_RNIBO4M[8]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \debounce_cntrrs[8]\, B => 
        un3_debounce_in_rs_1, C => RESET_set, Y => 
        \debounce_cntr[8]_net_1\);
    
    \debounce_cntr_RNIPQ221[15]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \debounce_cntrrs[15]\, B => 
        un3_debounce_in_rs_1, C => RESET_set, Y => 
        \debounce_cntr[15]_net_1\);
    
    \debounce_cntr_4[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => un1_debounce_cntr, B => 
        \debounce_cntr[0]_net_1\, Y => \debounce_cntr_4[0]_net_1\);
    
    \debounce_cntr[8]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_8_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[8]\);
    
    \debounce_cntr[0]\ : SLE
      port map(D => \debounce_cntr_4[0]_net_1\, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[0]_net_1\);
    
    \debounce_cntr_0[1]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_6_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[6]\);
    
    un3_debounce_cntr_1_cry_8 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[8]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_7\, S => 
        un3_debounce_cntr_1_cry_8_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_8\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr\ : CFG4
      generic map(INIT => x"8000")

      port map(A => un1_debounce_cntr_11, B => 
        un1_debounce_cntr_10, C => un1_debounce_cntr_8, D => 
        un1_debounce_cntr_9, Y => un1_debounce_cntr);
    
    un3_debounce_cntr_1_cry_12 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[12]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_11\, S => 
        un3_debounce_cntr_1_cry_12_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_12\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_11\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \debounce_cntr[7]\, B => \debounce_cntr[5]\, 
        C => \debounce_cntr[3]_net_1\, D => 
        \debounce_cntr[0]_net_1\, Y => un1_debounce_cntr_11);
    
    un3_debounce_cntr_1_s_15 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[15]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_14\, S => 
        un3_debounce_cntr_1_s_15_S_1, Y => OPEN, FCO => OPEN);
    
    un3_debounce_cntr_1_cry_10 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[10]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_9\, S => 
        un3_debounce_cntr_1_cry_10_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_10\);
    
    \debounce_cntr[2]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_2_S_1, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[2]_net_1\);
    
    \debounce_cntr[11]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_11_S_1, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => un2_debounce_in_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[11]_net_1\);
    
    un3_debounce_cntr_1_cry_1 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[1]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        un3_debounce_cntr_1_s_1_919_FCO, S => 
        un3_debounce_cntr_1_cry_1_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_1\);
    
    un3_debounce_cntr_1_cry_3 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[3]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_2\, S => 
        un3_debounce_cntr_1_cry_3_S_1, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_3\);
    
    \DEBOUNCE_PROC.un3_debounce_in\ : CFG2
      generic map(INIT => x"E")

      port map(A => DEBOUNCE_IN_c_0, B => RESET, Y => 
        un3_debounce_in_i);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity Debounce_0 is

    port( DEBOUNCE_IN_c_0  : in    std_logic;
          RESET            : in    std_logic;
          DEBOUNCE_OUT_1_c : out   std_logic;
          RESET_set        : in    std_logic;
          BIT_CLK          : in    std_logic
        );

end Debounce_0;

architecture DEF_ARCH of Debounce_0 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \debounce_cntr[1]_net_1\, VCC_net_1, 
        un2_debounce_in_i, un3_debounce_cntr_1_cry_1_S_0, 
        GND_net_1, \debounce_cntr[2]_net_1\, 
        un3_debounce_cntr_1_cry_2_S_0, \debounce_cntr[3]_net_1\, 
        un3_debounce_cntr_1_cry_3_S_0, \debounce_cntrrs[4]\, 
        un3_debounce_in_rs_0, \debounce_cntr[4]\, 
        un3_debounce_in_i, un3_debounce_cntr_1_cry_4_S_0, 
        \debounce_cntrrs[6]\, \debounce_cntr[6]\, 
        un3_debounce_cntr_1_cry_6_S_0, \debounce_cntr[5]\, 
        un3_debounce_cntr_1_cry_5_S_0, \debounce_cntr[7]\, 
        un3_debounce_cntr_1_cry_7_S_0, \debounce_cntrrs[8]\, 
        \debounce_cntr[8]_net_1\, un3_debounce_cntr_1_cry_8_S_0, 
        \debounce_cntrrs[9]\, \debounce_cntr[9]_net_1\, 
        un3_debounce_cntr_1_cry_9_S_0, \debounce_cntr[10]_net_1\, 
        un3_debounce_cntr_1_cry_10_S_0, \debounce_cntr[11]_net_1\, 
        un3_debounce_cntr_1_cry_11_S_0, \debounce_cntr[12]_net_1\, 
        un3_debounce_cntr_1_cry_12_S_0, \debounce_cntr[13]_net_1\, 
        un3_debounce_cntr_1_cry_13_S_0, \debounce_cntrrs[14]\, 
        \debounce_cntr[14]_net_1\, un3_debounce_cntr_1_cry_14_S_0, 
        \debounce_cntrrs[15]\, \debounce_cntr[15]_net_1\, 
        un3_debounce_cntr_1_s_15_S_0, \debounce_cntr[0]_net_1\, 
        \debounce_cntr_4[0]_net_1\, DEBOUNCE_OUT_1_crs, 
        un1_debounce_cntr, un3_debounce_cntr_1_s_1_918_FCO, 
        \un3_debounce_cntr_1_cry_1\, \un3_debounce_cntr_1_cry_2\, 
        \un3_debounce_cntr_1_cry_3\, \un3_debounce_cntr_1_cry_4\, 
        \un3_debounce_cntr_1_cry_5\, \un3_debounce_cntr_1_cry_6\, 
        \un3_debounce_cntr_1_cry_7\, \un3_debounce_cntr_1_cry_8\, 
        \un3_debounce_cntr_1_cry_9\, \un3_debounce_cntr_1_cry_10\, 
        \un3_debounce_cntr_1_cry_11\, 
        \un3_debounce_cntr_1_cry_12\, 
        \un3_debounce_cntr_1_cry_13\, 
        \un3_debounce_cntr_1_cry_14\, un1_debounce_cntr_11, 
        un1_debounce_cntr_10, un1_debounce_cntr_9, 
        un1_debounce_cntr_8 : std_logic;

begin 


    \debounce_cntr_0_0[0]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_5_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[5]\);
    
    un3_debounce_cntr_1_cry_9 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[9]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_8\, S => 
        un3_debounce_cntr_1_cry_9_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_9\);
    
    \debounce_cntr_0_RNIHHJ21[1]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => RESET_set, B => \debounce_cntrrs[6]\, C => 
        un3_debounce_in_rs_0, Y => \debounce_cntr[6]\);
    
    \debounce_cntr[12]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_12_S_0, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => un2_debounce_in_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[12]_net_1\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_8\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \debounce_cntr[2]_net_1\, B => 
        \debounce_cntr[1]_net_1\, C => \debounce_cntr[15]_net_1\, 
        D => \debounce_cntr[14]_net_1\, Y => un1_debounce_cntr_8);
    
    \DEBOUNCE_PROC.un3_debounce_in_rs\ : SLE
      port map(D => VCC_net_1, CLK => RESET, EN => VCC_net_1, ALn
         => un3_debounce_in_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => VCC_net_1, Q => 
        un3_debounce_in_rs_0);
    
    \debounce_cntr[15]\ : SLE
      port map(D => un3_debounce_cntr_1_s_15_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[15]\);
    
    un3_debounce_cntr_1_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_4\, S => 
        un3_debounce_cntr_1_cry_5_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_5\);
    
    un3_debounce_cntr_1_cry_2 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[2]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_1\, S => 
        un3_debounce_cntr_1_cry_2_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_2\);
    
    \debounce_cntr[3]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_3_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[3]_net_1\);
    
    un3_debounce_cntr_1_s_1_918 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[0]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => 
        OPEN, Y => OPEN, FCO => un3_debounce_cntr_1_s_1_918_FCO);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_9\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \debounce_cntr[9]_net_1\, B => 
        \debounce_cntr[8]_net_1\, C => \debounce_cntr[6]\, D => 
        \debounce_cntr[4]\, Y => un1_debounce_cntr_9);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_10\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \debounce_cntr[13]_net_1\, B => 
        \debounce_cntr[12]_net_1\, C => \debounce_cntr[11]_net_1\, 
        D => \debounce_cntr[10]_net_1\, Y => un1_debounce_cntr_10);
    
    debounce_out : SLE
      port map(D => un1_debounce_cntr, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => un3_debounce_in_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => DEBOUNCE_OUT_1_crs);
    
    \debounce_cntr[10]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_10_S_0, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => un2_debounce_in_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[10]_net_1\);
    
    un3_debounce_cntr_1_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_3\, S => 
        un3_debounce_cntr_1_cry_4_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_4\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \debounce_cntr[13]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_13_S_0, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => un2_debounce_in_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[13]_net_1\);
    
    un3_debounce_cntr_1_cry_14 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[14]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_13\, S => 
        un3_debounce_cntr_1_cry_14_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_14\);
    
    \debounce_cntr_0_0[1]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_7_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[7]\);
    
    un3_debounce_cntr_1_cry_13 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[13]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_12\, S => 
        un3_debounce_cntr_1_cry_13_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_13\);
    
    \debounce_cntr[9]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_9_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[9]\);
    
    un3_debounce_cntr_1_cry_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_6\, S => 
        un3_debounce_cntr_1_cry_7_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_7\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \DEBOUNCE_PROC.un2_debounce_in\ : CFG2
      generic map(INIT => x"2")

      port map(A => DEBOUNCE_IN_c_0, B => RESET, Y => 
        un2_debounce_in_i);
    
    \debounce_cntr[1]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_1_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[1]_net_1\);
    
    \debounce_cntr_0[0]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_4_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[4]\);
    
    \debounce_cntr_RNI9SS01[8]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => RESET_set, B => \debounce_cntrrs[8]\, C => 
        un3_debounce_in_rs_0, Y => \debounce_cntr[8]_net_1\);
    
    \debounce_cntr[14]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_14_S_0, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => un3_debounce_in_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[14]\);
    
    un3_debounce_cntr_1_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_5\, S => 
        un3_debounce_cntr_1_cry_6_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_6\);
    
    un3_debounce_cntr_1_cry_11 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[11]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_10\, S => 
        un3_debounce_cntr_1_cry_11_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_11\);
    
    \debounce_cntr_4[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => un1_debounce_cntr, B => 
        \debounce_cntr[0]_net_1\, Y => \debounce_cntr_4[0]_net_1\);
    
    \debounce_cntr_RNINT451[15]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => RESET_set, B => \debounce_cntrrs[15]\, C => 
        un3_debounce_in_rs_0, Y => \debounce_cntr[15]_net_1\);
    
    \debounce_cntr[8]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_8_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[8]\);
    
    \debounce_cntr[0]\ : SLE
      port map(D => \debounce_cntr_4[0]_net_1\, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[0]_net_1\);
    
    \debounce_cntr_0[1]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_6_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[6]\);
    
    un3_debounce_cntr_1_cry_8 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[8]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_7\, S => 
        un3_debounce_cntr_1_cry_8_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_8\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr\ : CFG4
      generic map(INIT => x"8000")

      port map(A => un1_debounce_cntr_11, B => 
        un1_debounce_cntr_10, C => un1_debounce_cntr_8, D => 
        un1_debounce_cntr_9, Y => un1_debounce_cntr);
    
    un3_debounce_cntr_1_cry_12 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[12]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_11\, S => 
        un3_debounce_cntr_1_cry_12_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_12\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_11\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \debounce_cntr[7]\, B => \debounce_cntr[5]\, 
        C => \debounce_cntr[3]_net_1\, D => 
        \debounce_cntr[0]_net_1\, Y => un1_debounce_cntr_11);
    
    un3_debounce_cntr_1_s_15 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[15]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_14\, S => 
        un3_debounce_cntr_1_s_15_S_0, Y => OPEN, FCO => OPEN);
    
    un3_debounce_cntr_1_cry_10 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[10]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_9\, S => 
        un3_debounce_cntr_1_cry_10_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_10\);
    
    \debounce_cntr_RNIMS451[14]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => RESET_set, B => \debounce_cntrrs[14]\, C => 
        un3_debounce_in_rs_0, Y => \debounce_cntr[14]_net_1\);
    
    \debounce_cntr_0_RNIGGJ21[0]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => RESET_set, B => \debounce_cntrrs[4]\, C => 
        un3_debounce_in_rs_0, Y => \debounce_cntr[4]\);
    
    debounce_out_RNIQS7T : CFG3
      generic map(INIT => x"EA")

      port map(A => DEBOUNCE_OUT_1_crs, B => un3_debounce_in_rs_0, 
        C => RESET_set, Y => DEBOUNCE_OUT_1_c);
    
    \debounce_cntr[2]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_2_S_0, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[2]_net_1\);
    
    \debounce_cntr[11]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_11_S_0, CLK => 
        BIT_CLK, EN => VCC_net_1, ALn => un2_debounce_in_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[11]_net_1\);
    
    \debounce_cntr_RNIATS01[9]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => RESET_set, B => \debounce_cntrrs[9]\, C => 
        un3_debounce_in_rs_0, Y => \debounce_cntr[9]_net_1\);
    
    un3_debounce_cntr_1_cry_1 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[1]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        un3_debounce_cntr_1_s_1_918_FCO, S => 
        un3_debounce_cntr_1_cry_1_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_1\);
    
    un3_debounce_cntr_1_cry_3 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[3]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_2\, S => 
        un3_debounce_cntr_1_cry_3_S_0, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_3\);
    
    \DEBOUNCE_PROC.un3_debounce_in\ : CFG2
      generic map(INIT => x"E")

      port map(A => DEBOUNCE_IN_c_0, B => RESET, Y => 
        un3_debounce_in_i);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity Debounce is

    port( DEBOUNCE_IN_c_0      : in    std_logic;
          DEBOUNCE_OUT_net_0_0 : out   std_logic;
          RESET                : in    std_logic;
          RESET_set            : in    std_logic;
          BIT_CLK              : in    std_logic
        );

end Debounce;

architecture DEF_ARCH of Debounce is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \debounce_cntr[1]_net_1\, VCC_net_1, 
        un2_debounce_in_i, un3_debounce_cntr_1_cry_1_S, GND_net_1, 
        \debounce_cntr[2]_net_1\, un3_debounce_cntr_1_cry_2_S, 
        \debounce_cntr[3]_net_1\, un3_debounce_cntr_1_cry_3_S, 
        \debounce_cntrrs[4]\, un3_debounce_in_rs, 
        \debounce_cntr[4]\, un3_debounce_in_i, 
        un3_debounce_cntr_1_cry_4_S, \debounce_cntrrs[6]\, 
        \debounce_cntr[6]\, un3_debounce_cntr_1_cry_6_S, 
        \debounce_cntr[5]\, un3_debounce_cntr_1_cry_5_S, 
        \debounce_cntr[7]\, un3_debounce_cntr_1_cry_7_S, 
        \debounce_cntrrs[8]\, \debounce_cntr[8]_net_1\, 
        un3_debounce_cntr_1_cry_8_S, \debounce_cntrrs[9]\, 
        \debounce_cntr[9]_net_1\, un3_debounce_cntr_1_cry_9_S, 
        \debounce_cntr[10]_net_1\, un3_debounce_cntr_1_cry_10_S, 
        \debounce_cntr[11]_net_1\, un3_debounce_cntr_1_cry_11_S, 
        \debounce_cntr[12]_net_1\, un3_debounce_cntr_1_cry_12_S, 
        \debounce_cntr[13]_net_1\, un3_debounce_cntr_1_cry_13_S, 
        \debounce_cntrrs[14]\, \debounce_cntr[14]_net_1\, 
        un3_debounce_cntr_1_cry_14_S, \debounce_cntrrs[15]\, 
        \debounce_cntr[15]_net_1\, un3_debounce_cntr_1_s_15_S, 
        \debounce_cntr[0]_net_1\, \debounce_cntr_4[0]_net_1\, 
        \DEBOUNCE_OUT_net_0rs[0]\, un1_debounce_cntr, 
        un3_debounce_cntr_1_s_1_917_FCO, 
        \un3_debounce_cntr_1_cry_1\, \un3_debounce_cntr_1_cry_2\, 
        \un3_debounce_cntr_1_cry_3\, \un3_debounce_cntr_1_cry_4\, 
        \un3_debounce_cntr_1_cry_5\, \un3_debounce_cntr_1_cry_6\, 
        \un3_debounce_cntr_1_cry_7\, \un3_debounce_cntr_1_cry_8\, 
        \un3_debounce_cntr_1_cry_9\, \un3_debounce_cntr_1_cry_10\, 
        \un3_debounce_cntr_1_cry_11\, 
        \un3_debounce_cntr_1_cry_12\, 
        \un3_debounce_cntr_1_cry_13\, 
        \un3_debounce_cntr_1_cry_14\, un1_debounce_cntr_11, 
        un1_debounce_cntr_10, un1_debounce_cntr_9, 
        un1_debounce_cntr_8 : std_logic;

begin 


    \debounce_cntr_0_0[0]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_5_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[5]\);
    
    un3_debounce_cntr_1_cry_9 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[9]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_8\, S => 
        un3_debounce_cntr_1_cry_9_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_9\);
    
    \debounce_cntr[12]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_12_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[12]_net_1\);
    
    un3_debounce_cntr_1_s_1_917 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[0]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => 
        OPEN, Y => OPEN, FCO => un3_debounce_cntr_1_s_1_917_FCO);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_8\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \debounce_cntr[2]_net_1\, B => 
        \debounce_cntr[1]_net_1\, C => \debounce_cntr[15]_net_1\, 
        D => \debounce_cntr[14]_net_1\, Y => un1_debounce_cntr_8);
    
    \DEBOUNCE_PROC.un3_debounce_in_rs\ : SLE
      port map(D => VCC_net_1, CLK => RESET, EN => VCC_net_1, ALn
         => un3_debounce_in_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => VCC_net_1, Q => 
        un3_debounce_in_rs);
    
    \debounce_cntr[15]\ : SLE
      port map(D => un3_debounce_cntr_1_s_15_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[15]\);
    
    un3_debounce_cntr_1_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_4\, S => 
        un3_debounce_cntr_1_cry_5_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_5\);
    
    un3_debounce_cntr_1_cry_2 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[2]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_1\, S => 
        un3_debounce_cntr_1_cry_2_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_2\);
    
    \debounce_cntr[3]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_3_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[3]_net_1\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_9\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \debounce_cntr[9]_net_1\, B => 
        \debounce_cntr[8]_net_1\, C => \debounce_cntr[6]\, D => 
        \debounce_cntr[4]\, Y => un1_debounce_cntr_9);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_10\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \debounce_cntr[13]_net_1\, B => 
        \debounce_cntr[12]_net_1\, C => \debounce_cntr[11]_net_1\, 
        D => \debounce_cntr[10]_net_1\, Y => un1_debounce_cntr_10);
    
    debounce_out : SLE
      port map(D => un1_debounce_cntr, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => un3_debounce_in_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \DEBOUNCE_OUT_net_0rs[0]\);
    
    \debounce_cntr[10]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_10_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[10]_net_1\);
    
    \debounce_cntr_RNI70LR[8]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => RESET_set, B => \debounce_cntrrs[8]\, C => 
        un3_debounce_in_rs, Y => \debounce_cntr[8]_net_1\);
    
    un3_debounce_cntr_1_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_3\, S => 
        un3_debounce_cntr_1_cry_4_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_4\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \debounce_cntr[13]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_13_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[13]_net_1\);
    
    un3_debounce_cntr_1_cry_14 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[14]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_13\, S => 
        un3_debounce_cntr_1_cry_14_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_14\);
    
    \debounce_cntr_0_0[1]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_7_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[7]\);
    
    \debounce_cntr_0_RNIFJUN[1]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => RESET_set, B => \debounce_cntrrs[6]\, C => 
        un3_debounce_in_rs, Y => \debounce_cntr[6]\);
    
    un3_debounce_cntr_1_cry_13 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[13]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_12\, S => 
        un3_debounce_cntr_1_cry_13_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_13\);
    
    \debounce_cntr[9]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_9_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[9]\);
    
    un3_debounce_cntr_1_cry_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_6\, S => 
        un3_debounce_cntr_1_cry_7_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_7\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \DEBOUNCE_PROC.un2_debounce_in\ : CFG2
      generic map(INIT => x"2")

      port map(A => DEBOUNCE_IN_c_0, B => RESET, Y => 
        un2_debounce_in_i);
    
    \debounce_cntr[1]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_1_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[1]_net_1\);
    
    \debounce_cntr_0[0]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_4_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[4]\);
    
    \debounce_cntr[14]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_14_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[14]\);
    
    un3_debounce_cntr_1_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_5\, S => 
        un3_debounce_cntr_1_cry_6_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_6\);
    
    un3_debounce_cntr_1_cry_11 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[11]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_10\, S => 
        un3_debounce_cntr_1_cry_11_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_11\);
    
    \debounce_cntr_4[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => un1_debounce_cntr, B => 
        \debounce_cntr[0]_net_1\, Y => \debounce_cntr_4[0]_net_1\);
    
    \debounce_cntr[8]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_8_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[8]\);
    
    \debounce_cntr[0]\ : SLE
      port map(D => \debounce_cntr_4[0]_net_1\, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[0]_net_1\);
    
    \debounce_cntr_0[1]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_6_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un3_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntrrs[6]\);
    
    \debounce_cntr_RNIKV6O[14]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => RESET_set, B => \debounce_cntrrs[14]\, C => 
        un3_debounce_in_rs, Y => \debounce_cntr[14]_net_1\);
    
    \debounce_cntr_RNI81LR[9]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => RESET_set, B => \debounce_cntrrs[9]\, C => 
        un3_debounce_in_rs, Y => \debounce_cntr[9]_net_1\);
    
    un3_debounce_cntr_1_cry_8 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[8]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_7\, S => 
        un3_debounce_cntr_1_cry_8_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_8\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr\ : CFG4
      generic map(INIT => x"8000")

      port map(A => un1_debounce_cntr_11, B => 
        un1_debounce_cntr_10, C => un1_debounce_cntr_8, D => 
        un1_debounce_cntr_9, Y => un1_debounce_cntr);
    
    un3_debounce_cntr_1_cry_12 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[12]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_11\, S => 
        un3_debounce_cntr_1_cry_12_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_12\);
    
    \DEBOUNCE_PROC.un1_debounce_cntr_11\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \debounce_cntr[7]\, B => \debounce_cntr[5]\, 
        C => \debounce_cntr[3]_net_1\, D => 
        \debounce_cntr[0]_net_1\, Y => un1_debounce_cntr_11);
    
    un3_debounce_cntr_1_s_15 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[15]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_14\, S => 
        un3_debounce_cntr_1_s_15_S, Y => OPEN, FCO => OPEN);
    
    un3_debounce_cntr_1_cry_10 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[10]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_9\, S => 
        un3_debounce_cntr_1_cry_10_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_10\);
    
    \debounce_cntr_0_RNIEIUN[0]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => RESET_set, B => \debounce_cntrrs[4]\, C => 
        un3_debounce_in_rs, Y => \debounce_cntr[4]\);
    
    \debounce_cntr[2]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_2_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[2]_net_1\);
    
    \debounce_cntr[11]\ : SLE
      port map(D => un3_debounce_cntr_1_cry_11_S, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => un2_debounce_in_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \debounce_cntr[11]_net_1\);
    
    debounce_out_RNIO4EU : CFG3
      generic map(INIT => x"EA")

      port map(A => \DEBOUNCE_OUT_net_0rs[0]\, B => 
        un3_debounce_in_rs, C => RESET_set, Y => 
        DEBOUNCE_OUT_net_0_0);
    
    un3_debounce_cntr_1_cry_1 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[1]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        un3_debounce_cntr_1_s_1_917_FCO, S => 
        un3_debounce_cntr_1_cry_1_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_1\);
    
    \debounce_cntr_RNIL07O[15]\ : CFG3
      generic map(INIT => x"EC")

      port map(A => RESET_set, B => \debounce_cntrrs[15]\, C => 
        un3_debounce_in_rs, Y => \debounce_cntr[15]_net_1\);
    
    un3_debounce_cntr_1_cry_3 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \debounce_cntr[3]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un3_debounce_cntr_1_cry_2\, S => 
        un3_debounce_cntr_1_cry_3_S, Y => OPEN, FCO => 
        \un3_debounce_cntr_1_cry_3\);
    
    \DEBOUNCE_PROC.un3_debounce_in\ : CFG2
      generic map(INIT => x"E")

      port map(A => DEBOUNCE_IN_c_0, B => RESET, Y => 
        un3_debounce_in_i);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity TriDebounce is

    port( DEBOUNCE_IN_c        : in    std_logic_vector(2 downto 0);
          DEBOUNCE_OUT_net_0_0 : out   std_logic;
          DEBOUNCE_OUT_2_c     : out   std_logic;
          DEBOUNCE_OUT_1_c     : out   std_logic;
          BIT_CLK              : in    std_logic;
          RESET_set            : in    std_logic;
          RESET                : in    std_logic
        );

end TriDebounce;

architecture DEF_ARCH of TriDebounce is 

  component Debounce_1
    port( DEBOUNCE_IN_c_0  : in    std_logic := 'U';
          RESET            : in    std_logic := 'U';
          DEBOUNCE_OUT_2_c : out   std_logic;
          RESET_set        : in    std_logic := 'U';
          BIT_CLK          : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component Debounce_0
    port( DEBOUNCE_IN_c_0  : in    std_logic := 'U';
          RESET            : in    std_logic := 'U';
          DEBOUNCE_OUT_1_c : out   std_logic;
          RESET_set        : in    std_logic := 'U';
          BIT_CLK          : in    std_logic := 'U'
        );
  end component;

  component Debounce
    port( DEBOUNCE_IN_c_0      : in    std_logic := 'U';
          DEBOUNCE_OUT_net_0_0 : out   std_logic;
          RESET                : in    std_logic := 'U';
          RESET_set            : in    std_logic := 'U';
          BIT_CLK              : in    std_logic := 'U'
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : Debounce_1
	Use entity work.Debounce_1(DEF_ARCH);
    for all : Debounce_0
	Use entity work.Debounce_0(DEF_ARCH);
    for all : Debounce
	Use entity work.Debounce(DEF_ARCH);
begin 


    DEBOUNCE_2_INST : Debounce_1
      port map(DEBOUNCE_IN_c_0 => DEBOUNCE_IN_c(2), RESET => 
        RESET, DEBOUNCE_OUT_2_c => DEBOUNCE_OUT_2_c, RESET_set
         => RESET_set, BIT_CLK => BIT_CLK);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    DEBOUNCE_1_INST : Debounce_0
      port map(DEBOUNCE_IN_c_0 => DEBOUNCE_IN_c(1), RESET => 
        RESET, DEBOUNCE_OUT_1_c => DEBOUNCE_OUT_1_c, RESET_set
         => RESET_set, BIT_CLK => BIT_CLK);
    
    DEBOUNCE_0_INST : Debounce
      port map(DEBOUNCE_IN_c_0 => DEBOUNCE_IN_c(0), 
        DEBOUNCE_OUT_net_0_0 => DEBOUNCE_OUT_net_0_0, RESET => 
        RESET, RESET_set => RESET_set, BIT_CLK => BIT_CLK);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CRC16_Generator_0 is

    port( TX_FIFO_DOUT   : in    std_logic_vector(7 downto 0);
          tx_crc_data    : out   std_logic_vector(15 downto 0);
          tx_crc_gen     : in    std_logic;
          byte_clk_en    : in    std_logic;
          BIT_CLK        : in    std_logic;
          tx_crc_reset_i : in    std_logic
        );

end CRC16_Generator_0;

architecture DEF_ARCH of CRC16_Generator_0 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \tx_crc_data[13]\, GND_net_1, \tx_crc_data[5]\, 
        \lfsr_q_0_sqmuxa\, VCC_net_1, \tx_crc_data[14]\, 
        \tx_crc_data[6]\, \tx_crc_data[15]\, \lfsr_c[15]\, 
        \tx_crc_data[0]\, \lfsr_c[0]\, \tx_crc_data[1]\, 
        \lfsr_c[1]\, \tx_crc_data[2]\, N_179_i, \tx_crc_data[3]\, 
        N_184_i, \tx_crc_data[4]\, N_183_i, N_181_i, N_182_i, 
        \tx_crc_data[7]\, N_185_i, \tx_crc_data[8]\, N_79_i_i, 
        \tx_crc_data[9]\, \lfsr_c[9]\, \tx_crc_data[10]\, 
        \tx_crc_data[11]\, \tx_crc_data[12]\, N_150_i
         : std_logic;

begin 

    tx_crc_data(15) <= \tx_crc_data[15]\;
    tx_crc_data(14) <= \tx_crc_data[14]\;
    tx_crc_data(13) <= \tx_crc_data[13]\;
    tx_crc_data(12) <= \tx_crc_data[12]\;
    tx_crc_data(11) <= \tx_crc_data[11]\;
    tx_crc_data(10) <= \tx_crc_data[10]\;
    tx_crc_data(9) <= \tx_crc_data[9]\;
    tx_crc_data(8) <= \tx_crc_data[8]\;
    tx_crc_data(7) <= \tx_crc_data[7]\;
    tx_crc_data(6) <= \tx_crc_data[6]\;
    tx_crc_data(5) <= \tx_crc_data[5]\;
    tx_crc_data(4) <= \tx_crc_data[4]\;
    tx_crc_data(3) <= \tx_crc_data[3]\;
    tx_crc_data(2) <= \tx_crc_data[2]\;
    tx_crc_data(1) <= \tx_crc_data[1]\;
    tx_crc_data(0) <= \tx_crc_data[0]\;

    \lfsr_q[9]\ : SLE
      port map(D => \lfsr_c[9]\, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[9]\);
    
    \lfsr_c_0_a2_0_x2_2_x2[7]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \tx_crc_data[14]\, B => \tx_crc_data[13]\, C
         => TX_FIFO_DOUT(6), D => TX_FIFO_DOUT(5), Y => N_185_i);
    
    \lfsr_q[6]\ : SLE
      port map(D => N_182_i, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[6]\);
    
    \lfsr_q[3]\ : SLE
      port map(D => N_184_i, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[3]\);
    
    \lfsr_q[10]\ : SLE
      port map(D => \tx_crc_data[2]\, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[10]\);
    
    \lfsr_c_0_a2_1_0_x2_0_x2[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => TX_FIFO_DOUT(7), B => \tx_crc_data[15]\, Y
         => N_150_i);
    
    \lfsr_q[2]\ : SLE
      port map(D => N_179_i, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[2]\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \lfsr_q[1]\ : SLE
      port map(D => \lfsr_c[1]\, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[1]\);
    
    \lfsr_q[7]\ : SLE
      port map(D => N_185_i, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[7]\);
    
    \lfsr_c_0_a2_0_x2_1_x2[3]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \tx_crc_data[9]\, B => \tx_crc_data[10]\, C
         => TX_FIFO_DOUT(2), D => TX_FIFO_DOUT(1), Y => N_184_i);
    
    \lfsr_q[4]\ : SLE
      port map(D => N_183_i, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[4]\);
    
    \lfsr_q[11]\ : SLE
      port map(D => \tx_crc_data[3]\, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[11]\);
    
    \lfsr_q[5]\ : SLE
      port map(D => N_181_i, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[5]\);
    
    \lfsr_c_0_a2[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => N_150_i, B => \tx_crc_data[1]\, Y => 
        \lfsr_c[9]\);
    
    \lfsr_c_0_a2[1]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => N_181_i, B => N_184_i, C => N_150_i, D => 
        N_185_i, Y => \lfsr_c[1]\);
    
    \lfsr_q[0]\ : SLE
      port map(D => \lfsr_c[0]\, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[0]\);
    
    \lfsr_c_0_a2[15]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => TX_FIFO_DOUT(0), B => \lfsr_c[1]\, C => 
        \tx_crc_data[7]\, D => \tx_crc_data[8]\, Y => 
        \lfsr_c[15]\);
    
    \lfsr_q[12]\ : SLE
      port map(D => \tx_crc_data[4]\, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[12]\);
    
    \lfsr_c_0_a2_2_x2_1_x2[4]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \tx_crc_data[11]\, B => \tx_crc_data[10]\, C
         => TX_FIFO_DOUT(3), D => TX_FIFO_DOUT(2), Y => N_183_i);
    
    \lfsr_c_0_a2_2_x2_1_x2[2]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \tx_crc_data[9]\, B => \tx_crc_data[8]\, C
         => TX_FIFO_DOUT(1), D => TX_FIFO_DOUT(0), Y => N_179_i);
    
    lfsr_q_0_sqmuxa : CFG2
      generic map(INIT => x"8")

      port map(A => byte_clk_en, B => tx_crc_gen, Y => 
        \lfsr_q_0_sqmuxa\);
    
    \lfsr_c_0_a2_0_x2_0_x2[5]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \tx_crc_data[12]\, B => \tx_crc_data[11]\, C
         => TX_FIFO_DOUT(4), D => TX_FIFO_DOUT(3), Y => N_181_i);
    
    \lfsr_q[14]\ : SLE
      port map(D => \tx_crc_data[6]\, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[14]\);
    
    \lfsr_c_0_a2_i_x2[8]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \tx_crc_data[14]\, B => \tx_crc_data[0]\, C
         => N_150_i, D => TX_FIFO_DOUT(6), Y => N_79_i_i);
    
    \lfsr_c_0_a2_2_x2_1_x2[6]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \tx_crc_data[13]\, B => \tx_crc_data[12]\, C
         => TX_FIFO_DOUT(5), D => TX_FIFO_DOUT(4), Y => N_182_i);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \lfsr_q[8]\ : SLE
      port map(D => N_79_i_i, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[8]\);
    
    \lfsr_q[13]\ : SLE
      port map(D => \tx_crc_data[5]\, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[13]\);
    
    \lfsr_c_0_a2[0]\ : CFG3
      generic map(INIT => x"96")

      port map(A => TX_FIFO_DOUT(0), B => \lfsr_c[1]\, C => 
        \tx_crc_data[8]\, Y => \lfsr_c[0]\);
    
    \lfsr_q[15]\ : SLE
      port map(D => \lfsr_c[15]\, CLK => BIT_CLK, EN => 
        \lfsr_q_0_sqmuxa\, ALn => tx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_crc_data[15]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity TX_Collision_Detector is

    port( RESET               : in    std_logic;
          external_loopback   : in    std_logic;
          internal_loopback   : in    std_logic;
          DRVR_EN_c           : in    std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          tx_col_detect_en    : out   std_logic
        );

end TX_Collision_Detector;

architecture DEF_ARCH of TX_Collision_Detector is 

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \tx_col_detect_en_0\, GND_net_1, 
        un10_reset : std_logic;

begin 


    tx_col_detect_en_0 : CFG2
      generic map(INIT => x"4")

      port map(A => un10_reset, B => DRVR_EN_c, Y => 
        \tx_col_detect_en_0\);
    
    \tx_col_detect_en\ : SLE
      port map(D => \tx_col_detect_en_0\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => tx_col_detect_en);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \SYNCH_PROC.un10_reset\ : CFG3
      generic map(INIT => x"FE")

      port map(A => internal_loopback, B => external_loopback, C
         => RESET, Y => un10_reset);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity IdleLineDetector_0 is

    port( manches_in_dly      : in    std_logic_vector(1 downto 0);
          idle_line5          : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          RESET_i             : in    std_logic;
          tx_idle_line        : out   std_logic
        );

end IdleLineDetector_0;

architecture DEF_ARCH of IdleLineDetector_0 is 

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \idle_line_cntr_0_sqmuxa\, GND_net_1, 
        \idle_line_cntr[0]_net_1\, \idle_line_cntr_s[0]\, 
        \idle_line_cntr[1]_net_1\, \idle_line_cntr_s[1]\, 
        \idle_line_cntr[2]_net_1\, \idle_line_cntr_s[2]\, 
        \idle_line_cntr[3]_net_1\, \idle_line_cntr_s[3]\, 
        \idle_line_cntr[4]_net_1\, \idle_line_cntr_s[4]\, 
        \idle_line_cntr[5]_net_1\, \idle_line_cntr_s[5]\, 
        \idle_line_cntr[6]_net_1\, \idle_line_cntr_s[6]\, 
        \idle_line_cntr[7]_net_1\, \idle_line_cntr_s[7]\, 
        \idle_line_cntr[8]_net_1\, \idle_line_cntr_s[8]\, 
        \idle_line_cntr[9]_net_1\, \idle_line_cntr_s[9]\, 
        \idle_line_cntr[10]_net_1\, \idle_line_cntr_s[10]\, 
        \idle_line_cntr[11]_net_1\, \idle_line_cntr_s[11]\, 
        \idle_line_cntr[12]_net_1\, \idle_line_cntr_s[12]\, 
        \idle_line_cntr[13]_net_1\, \idle_line_cntr_s[13]\, 
        \idle_line_cntr[14]_net_1\, \idle_line_cntr_s[14]\, 
        \idle_line_cntr[15]_net_1\, \idle_line_cntr_s[15]\, 
        idle_line_cntr_cry_cy, un5_manches_in_dly_9_RNIQSC51_Y, 
        \idle_line5\, un5_manches_in_dly_9, un5_manches_in_dly_10, 
        un5_manches_in_dly_11, \idle_line_cntr_cry[0]\, 
        \idle_line_cntr_cry[1]\, \idle_line_cntr_cry[2]\, 
        \idle_line_cntr_cry[3]\, \idle_line_cntr_cry[4]\, 
        \idle_line_cntr_cry[5]\, \idle_line_cntr_cry[6]\, 
        \idle_line_cntr_cry[7]\, \idle_line_cntr_cry[8]\, 
        \idle_line_cntr_cry[9]\, \idle_line_cntr_cry[10]\, 
        \idle_line_cntr_cry[11]\, \idle_line_cntr_cry[12]\, 
        \idle_line_cntr_cry[13]\, \idle_line_cntr_cry[14]\, 
        un5_manches_in_dly_8 : std_logic;

begin 

    idle_line5 <= \idle_line5\;

    \idle_line_cntr_RNICPKC7[3]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[3]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[2]\, S => \idle_line_cntr_s[3]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[3]\);
    
    idle_line : SLE
      port map(D => \idle_line_cntr_0_sqmuxa\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => tx_idle_line);
    
    \IDLE_LINE_DETECT_PROC.un5_manches_in_dly_11\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \idle_line_cntr[11]_net_1\, B => 
        \idle_line_cntr[8]_net_1\, C => \idle_line_cntr[7]_net_1\, 
        D => un5_manches_in_dly_8, Y => un5_manches_in_dly_11);
    
    idle_line_cntr_0_sqmuxa : CFG4
      generic map(INIT => x"4000")

      port map(A => \idle_line5\, B => un5_manches_in_dly_11, C
         => un5_manches_in_dly_10, D => un5_manches_in_dly_9, Y
         => \idle_line_cntr_0_sqmuxa\);
    
    \idle_line_cntr_RNIE6TJD[7]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[7]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[6]\, S => \idle_line_cntr_s[7]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[7]\);
    
    \idle_line_cntr_RNIV6IUO[14]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[14]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[13]\, S => \idle_line_cntr_s[14]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[14]\);
    
    \idle_line_cntr[4]\ : SLE
      port map(D => \idle_line_cntr_s[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[4]_net_1\);
    
    \idle_line_cntr[14]\ : SLE
      port map(D => \idle_line_cntr_s[14]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[14]_net_1\);
    
    \idle_line_cntr_RNIDQ6N2[0]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[0]_net_1\, D => GND_net_1, FCI => 
        idle_line_cntr_cry_cy, S => \idle_line_cntr_s[0]\, Y => 
        OPEN, FCO => \idle_line_cntr_cry[0]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \idle_line_cntr_RNIG5T0M[12]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[12]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[11]\, S => \idle_line_cntr_s[12]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[12]\);
    
    \IDLE_LINE_DETECT_PROC.un5_manches_in_dly_9\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \idle_line_cntr[10]_net_1\, B => 
        \idle_line_cntr[9]_net_1\, C => \idle_line_cntr[2]_net_1\, 
        D => \idle_line_cntr[1]_net_1\, Y => un5_manches_in_dly_9);
    
    \IDLE_LINE_DETECT_PROC.un5_manches_in_dly_10\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \idle_line_cntr[6]_net_1\, B => 
        \idle_line_cntr[5]_net_1\, C => \idle_line_cntr[4]_net_1\, 
        D => \idle_line_cntr[3]_net_1\, Y => 
        un5_manches_in_dly_10);
    
    \idle_line_cntr_RNINLNFN[13]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[13]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[12]\, S => \idle_line_cntr_s[13]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[13]\);
    
    \idle_line_cntr[9]\ : SLE
      port map(D => \idle_line_cntr_s[9]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[9]_net_1\);
    
    \idle_line_cntr[8]\ : SLE
      port map(D => \idle_line_cntr_s[8]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[8]_net_1\);
    
    \idle_line_cntr[7]\ : SLE
      port map(D => \idle_line_cntr_s[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[7]_net_1\);
    
    \idle_line_cntr[15]\ : SLE
      port map(D => \idle_line_cntr_s[15]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[15]_net_1\);
    
    \idle_line_cntr_RNIAM2IK[11]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[11]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[10]\, S => \idle_line_cntr_s[11]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[11]\);
    
    \idle_line_cntr_RNI5883J[10]\ : ARI1
      generic map(INIT => x"4D800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[10]_net_1\, D => 
        \idle_line_cntr_0_sqmuxa\, FCI => \idle_line_cntr_cry[9]\, 
        S => \idle_line_cntr_s[10]\, Y => OPEN, FCO => 
        \idle_line_cntr_cry[10]\);
    
    \idle_line_cntr[11]\ : SLE
      port map(D => \idle_line_cntr_s[11]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[11]_net_1\);
    
    \idle_line_cntr[10]\ : SLE
      port map(D => \idle_line_cntr_s[10]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[10]_net_1\);
    
    \idle_line_cntr[1]\ : SLE
      port map(D => \idle_line_cntr_s[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[1]_net_1\);
    
    \idle_line_cntr_RNIK132C[6]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[6]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[5]\, S => \idle_line_cntr_s[6]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[6]\);
    
    \IDLE_LINE_DETECT_PROC.un5_manches_in_dly_8\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \idle_line_cntr[15]_net_1\, B => 
        \idle_line_cntr[14]_net_1\, C => 
        \idle_line_cntr[13]_net_1\, D => 
        \idle_line_cntr[12]_net_1\, Y => un5_manches_in_dly_8);
    
    \idle_line_cntr_RNI9CN5F[8]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[8]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[7]\, S => \idle_line_cntr_s[8]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[8]\);
    
    \idle_line_cntr_RNO[15]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[15]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[14]\, S => \idle_line_cntr_s[15]\, Y
         => OPEN, FCO => OPEN);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \idle_line_cntr_RNI1P094[1]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[1]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[0]\, S => \idle_line_cntr_s[1]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[1]\);
    
    \idle_line_cntr[6]\ : SLE
      port map(D => \idle_line_cntr_s[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[6]_net_1\);
    
    \idle_line_cntr_RNIMOQQ5[2]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[2]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[1]\, S => \idle_line_cntr_s[2]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[2]\);
    
    \idle_line_cntr_RNI3REU8[4]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[4]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[3]\, S => \idle_line_cntr_s[4]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[4]\);
    
    \idle_line_cntr_RNIRT8GA[5]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[5]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[4]\, S => \idle_line_cntr_s[5]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[5]\);
    
    \idle_line_cntr[13]\ : SLE
      port map(D => \idle_line_cntr_s[13]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[13]_net_1\);
    
    \idle_line_cntr[0]\ : SLE
      port map(D => \idle_line_cntr_s[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[0]_net_1\);
    
    \idle_line_cntr_RNI3NV5H[9]\ : ARI1
      generic map(INIT => x"4D800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNIQSC51_Y, C => 
        \idle_line_cntr[9]_net_1\, D => \idle_line_cntr_0_sqmuxa\, 
        FCI => \idle_line_cntr_cry[8]\, S => 
        \idle_line_cntr_s[9]\, Y => OPEN, FCO => 
        \idle_line_cntr_cry[9]\);
    
    \IDLE_LINE_DETECT_PROC.un5_manches_in_dly_9_RNIQSC51\ : ARI1
      generic map(INIT => x"41555")

      port map(A => un5_manches_in_dly_11, B => \idle_line5\, C
         => un5_manches_in_dly_9, D => un5_manches_in_dly_10, FCI
         => VCC_net_1, S => OPEN, Y => 
        un5_manches_in_dly_9_RNIQSC51_Y, FCO => 
        idle_line_cntr_cry_cy);
    
    \idle_line_cntr[12]\ : SLE
      port map(D => \idle_line_cntr_s[12]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[12]_net_1\);
    
    \idle_line_cntr[3]\ : SLE
      port map(D => \idle_line_cntr_s[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[3]_net_1\);
    
    un4_manches_in_dly : CFG2
      generic map(INIT => x"6")

      port map(A => manches_in_dly(1), B => manches_in_dly(0), Y
         => \idle_line5\);
    
    \idle_line_cntr[5]\ : SLE
      port map(D => \idle_line_cntr_s[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[5]_net_1\);
    
    \idle_line_cntr[2]\ : SLE
      port map(D => \idle_line_cntr_s[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[2]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity TX_SM is

    port( manches_in_dly      : in    std_logic_vector(1 downto 0);
          TX_FIFO_DOUT        : in    std_logic_vector(7 downto 0);
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          idle_line5          : out   std_logic;
          N_114               : out   std_logic;
          TX_FIFO_Empty       : in    std_logic;
          TX_DataEn           : out   std_logic;
          TX_PreAmble         : out   std_logic;
          tx_crc_byte1_en     : out   std_logic;
          tx_crc_byte2_en     : out   std_logic;
          tx_packet_complt    : out   std_logic;
          tx_crc_gen          : out   std_logic;
          start_tx_FIFO       : in    std_logic;
          DRVR_EN_c           : out   std_logic;
          byte_clk_en         : in    std_logic;
          tx_preamble_pat_en  : out   std_logic;
          BIT_CLK             : in    std_logic;
          RESET_i             : in    std_logic
        );

end TX_SM;

architecture DEF_ARCH of TX_SM is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component IdleLineDetector_0
    port( manches_in_dly      : in    std_logic_vector(1 downto 0) := (others => 'U');
          idle_line5          : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          RESET_i             : in    std_logic := 'U';
          tx_idle_line        : out   std_logic
        );
  end component;

    signal \TX_STATE[8]_net_1\, \TX_STATE_i_0[8]\, 
        \un25_tx_byte_cntr_a_4[6]\, GND_net_1, 
        \un25_tx_byte_cntr_a_4_i[6]\, un1_byte_clk_en_inv_2_i, 
        VCC_net_1, \un25_tx_byte_cntr_a_4[7]\, 
        \un25_tx_byte_cntr_a_4_i[7]\, \un25_tx_byte_cntr_a_4[8]\, 
        \un25_tx_byte_cntr_a_4_i[8]\, \un25_tx_byte_cntr_a_4[9]\, 
        \un25_tx_byte_cntr_a_4_i[9]\, \un25_tx_byte_cntr_a_4[10]\, 
        \un25_tx_byte_cntr_a_4_i[10]\, 
        \un25_tx_byte_cntr_a_4[11]\, 
        \un25_tx_byte_cntr_a_4_i[11]\, 
        \tx_packet_length[1]_net_1\, 
        \un25_tx_byte_cntr_a_4_i_i[1]\, 
        \tx_packet_length[2]_net_1\, 
        un25_tx_byte_cntr_a_4_axb_1_i, 
        \tx_packet_length[3]_net_1\, 
        un25_tx_byte_cntr_a_4_axb_2_i, 
        \tx_packet_length[4]_net_1\, 
        un25_tx_byte_cntr_a_4_axb_3_i, 
        \tx_packet_length[5]_net_1\, N_49_i, 
        \tx_packet_length[6]_net_1\, 
        un25_tx_byte_cntr_a_4_axb_5_i, 
        \tx_packet_length[7]_net_1\, 
        un25_tx_byte_cntr_a_4_axb_6_i, 
        \tx_packet_length[8]_net_1\, N_10_i, 
        \tx_packet_length[9]_net_1\, 
        un25_tx_byte_cntr_a_4_axb_8_i, 
        \tx_packet_length[10]_net_1\, 
        un25_tx_byte_cntr_a_4_axb_9_i, \un25_tx_byte_cntr_a_4[1]\, 
        un25_tx_byte_cntr_a_4_cry_0_Y, \un25_tx_byte_cntr_a_4[2]\, 
        \un25_tx_byte_cntr_a_4_i[2]\, \un25_tx_byte_cntr_a_4[3]\, 
        \un25_tx_byte_cntr_a_4_i[3]\, \un25_tx_byte_cntr_a_4[4]\, 
        \un25_tx_byte_cntr_a_4_i[4]\, \un25_tx_byte_cntr_a_4[5]\, 
        \un25_tx_byte_cntr_a_4_i[5]\, \tx_packet_length[0]_net_1\, 
        N_12_i, TX_DataEn_1_m, \tx_idle_line_s\, tx_idle_line, 
        \start_tx_FIFO_s\, \TX_STATE[3]_net_1\, \TX_STATE_69\, 
        \TX_STATE[4]_net_1\, \TX_STATE_68\, \TX_STATE[5]_net_1\, 
        \TX_STATE_67\, \TX_STATE[6]_net_1\, \TX_STATE_66\, 
        \TX_STATE[7]_net_1\, \TX_STATE_65\, \TX_STATE_64\, 
        un1_tx_packet_length_0_sqmuxa_o, 
        \iTX_FIFO_rd_en_ret_1_RNO\, TX_DataEn_1_o, N_163, 
        \tx_byte_cntr_cry_cy_Y[0]\, \TX_STATE[0]_net_1\, 
        \TX_STATE[2]_net_1\, TX_PreAmble_net_1, \TX_PreAmble_34\, 
        TX_DataEn_7, \TX_STATE_72\, \TX_STATE[1]_net_1\, 
        \TX_STATE_71\, \TX_STATE_70\, \PostAmble_cntr[0]_net_1\, 
        \PostAmble_cntr_s[0]\, \PostAmble_cntr[1]_net_1\, 
        \PostAmble_cntr_s[1]\, \PostAmble_cntr[2]_net_1\, 
        \PostAmble_cntr_s[2]\, \PostAmble_cntr[3]_net_1\, 
        \PostAmble_cntr_s[3]\, \PostAmble_cntr[4]_net_1\, 
        \PostAmble_cntr_s[4]\, \PostAmble_cntr[5]_net_1\, 
        \PostAmble_cntr_s[5]\, \PostAmble_cntr[6]_net_1\, 
        \PostAmble_cntr_s[6]\, \PostAmble_cntr[7]_net_1\, 
        \PostAmble_cntr_s[7]\, \PostAmble_cntr[8]_net_1\, 
        \PostAmble_cntr_s[8]\, \PostAmble_cntr[9]_net_1\, 
        \PostAmble_cntr_s[9]\, \PostAmble_cntr[10]_net_1\, 
        \PostAmble_cntr_s[10]\, \PostAmble_cntr[11]_net_1\, 
        \PostAmble_cntr_s[11]\, \txen_early_cntr[0]_net_1\, 
        \txen_early_cntr_s[0]\, \txen_early_cntr[1]_net_1\, 
        \txen_early_cntr_s[1]\, \txen_early_cntr[2]_net_1\, 
        \txen_early_cntr_s[2]\, \txen_early_cntr[3]_net_1\, 
        \txen_early_cntr_s[3]\, \txen_early_cntr[4]_net_1\, 
        \txen_early_cntr_s[4]\, \txen_early_cntr[5]_net_1\, 
        \txen_early_cntr_s[5]\, \txen_early_cntr[6]_net_1\, 
        \txen_early_cntr_s[6]\, \txen_early_cntr[7]_net_1\, 
        \txen_early_cntr_s[7]\, \txen_early_cntr[8]_net_1\, 
        \txen_early_cntr_s[8]\, \txen_early_cntr[9]_net_1\, 
        \txen_early_cntr_s[9]\, \txen_early_cntr[10]_net_1\, 
        \txen_early_cntr_s[10]\, \txen_early_cntr[11]_net_1\, 
        \txen_early_cntr_s[11]\, \tx_byte_cntr[0]_net_1\, 
        \tx_byte_cntr_s[0]\, \tx_byte_cntr[1]_net_1\, 
        \tx_byte_cntr_s[1]\, \tx_byte_cntr[2]_net_1\, 
        \tx_byte_cntr_s[2]\, \tx_byte_cntr[3]_net_1\, 
        \tx_byte_cntr_s[3]\, \tx_byte_cntr[4]_net_1\, 
        \tx_byte_cntr_s[4]\, \tx_byte_cntr[5]_net_1\, 
        \tx_byte_cntr_s[5]\, \tx_byte_cntr[6]_net_1\, 
        \tx_byte_cntr_s[6]\, \tx_byte_cntr[7]_net_1\, 
        \tx_byte_cntr_s[7]\, \tx_byte_cntr[8]_net_1\, 
        \tx_byte_cntr_s[8]\, \tx_byte_cntr[9]_net_1\, 
        \tx_byte_cntr_s[9]\, \tx_byte_cntr[10]_net_1\, 
        \tx_byte_cntr_s[10]\, \tx_byte_cntr[11]_net_1\, 
        \tx_byte_cntr_s[11]_net_1\, \PreAmble_cntr[0]_net_1\, 
        \PreAmble_cntr_s[0]\, N_17_i, \PreAmble_cntr[1]_net_1\, 
        \PreAmble_cntr_s[1]\, \PreAmble_cntr[2]_net_1\, 
        \PreAmble_cntr_s[2]\, \PreAmble_cntr[3]_net_1\, 
        \PreAmble_cntr_s[3]\, \PreAmble_cntr[4]_net_1\, 
        \PreAmble_cntr_s[4]\, \PreAmble_cntr[5]_net_1\, 
        \PreAmble_cntr_s[5]\, \PreAmble_cntr[6]_net_1\, 
        \PreAmble_cntr_s[6]\, PostAmble_cntr_cry_cy, 
        tx_state29_6_RNI9SJ61_Y, tx_state29_6, tx_state29_7, 
        tx_state29_8, \PostAmble_cntr_cry[0]\, 
        \PostAmble_cntr_cry[1]\, \PostAmble_cntr_cry[2]\, 
        \PostAmble_cntr_cry[3]\, \PostAmble_cntr_cry[4]\, 
        \PostAmble_cntr_cry[5]\, \PostAmble_cntr_cry[6]\, 
        \PostAmble_cntr_cry[7]\, \PostAmble_cntr_cry[8]\, 
        \PostAmble_cntr_cry[9]\, \PostAmble_cntr_cry[10]\, 
        txen_early_cntr_cry_cy, \TX_STATE_RNIAIGV2_Y[7]\, m15_e_6, 
        m15_e_7, m15_e_8, \txen_early_cntr_cry[0]\, 
        \txen_early_cntr_cry[1]\, \txen_early_cntr_cry[2]\, 
        \txen_early_cntr_cry[3]\, \txen_early_cntr_cry[4]\, 
        \txen_early_cntr_cry[5]\, \txen_early_cntr_cry[6]\, 
        \txen_early_cntr_cry[7]\, \txen_early_cntr_cry[8]\, 
        \txen_early_cntr_cry[9]\, \txen_early_cntr_cry[10]\, 
        tx_byte_cntr_cry_cy, \tx_byte_cntr_cry[0]_net_1\, 
        \tx_byte_cntr_cry[1]_net_1\, \tx_byte_cntr_cry[2]_net_1\, 
        \tx_byte_cntr_cry[3]_net_1\, \tx_byte_cntr_cry[4]_net_1\, 
        \tx_byte_cntr_cry[5]_net_1\, \tx_byte_cntr_cry[6]_net_1\, 
        \tx_byte_cntr_cry[7]_net_1\, \tx_byte_cntr_cry[8]_net_1\, 
        \tx_byte_cntr_cry[9]_net_1\, \tx_byte_cntr_cry[10]_net_1\, 
        PreAmble_cntr_cry_cy, \PreAmble_cntr_RNIHNV31_Y[6]\, 
        PreAmble_cntr_0_sqmuxa_0_83_i_o3_0, 
        PreAmble_cntr_0_sqmuxa_0_83_i_o3_4, 
        \PreAmble_cntr_cry[0]\, \PreAmble_cntr_cry[1]\, 
        \PreAmble_cntr_cry[2]\, \PreAmble_cntr_cry[3]\, 
        \PreAmble_cntr_cry[4]\, \PreAmble_cntr_cry[5]\, 
        un25_tx_byte_cntr_a_4_cry_0, N_81, 
        un25_tx_byte_cntr_a_4_cry_1, un25_tx_byte_cntr_a_4_cry_2, 
        un25_tx_byte_cntr_a_4_cry_3, un25_tx_byte_cntr_a_4_cry_4, 
        un25_tx_byte_cntr_a_4_cry_5, un25_tx_byte_cntr_a_4_cry_6, 
        un25_tx_byte_cntr_a_4_cry_7, un25_tx_byte_cntr_a_4_cry_8, 
        \un25_tx_byte_cntr_1_data_tmp[0]\, 
        \un25_tx_byte_cntr_1_data_tmp[1]\, 
        \un25_tx_byte_cntr_1_data_tmp[2]\, 
        \un25_tx_byte_cntr_1_data_tmp[3]\, 
        \un25_tx_byte_cntr_1_data_tmp[4]\, un25_tx_byte_cntr, 
        un25_tx_byte_cntr_a_4_s_9_931_FCO, N_213_i, 
        un25_tx_byte_cntr_a_4_s_9_sf, m56_i_0_0, 
        un14_tx_byte_cntr_0_a2_8_a2_0_1_0, un9_start_tx_fifo_s, 
        N_360, \un1_byte_clk_en_inv_2_0_0_2\, N_403, N_402, 
        un14_tx_byte_cntr_0_a2_8_a2_0_5, N_80, N_513, N_471, 
        un14_tx_byte_cntr_0_a2_8_a2_0_6, N_554, N_362, N_511
         : std_logic;

    for all : IdleLineDetector_0
	Use entity work.IdleLineDetector_0(DEF_ARCH);
begin 

    TX_PreAmble <= TX_PreAmble_net_1;

    iTX_FIFO_rd_en_ret_1 : SLE
      port map(D => \iTX_FIFO_rd_en_ret_1_RNO\, CLK => BIT_CLK, 
        EN => VCC_net_1, ALn => RESET_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        un1_tx_packet_length_0_sqmuxa_o);
    
    \tx_packet_length_RNO[2]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => N_81, B => TX_FIFO_DOUT(2), C => 
        \tx_packet_length[2]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => un25_tx_byte_cntr_a_4_axb_1_i);
    
    \txen_early_cntr_RNIJFKLC[2]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \TX_STATE_RNIAIGV2_Y[7]\, C
         => \txen_early_cntr[2]_net_1\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[1]\, S => \txen_early_cntr_s[2]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[2]\);
    
    \TX_STATE_ns_8_0_.m56_i_0_a2\ : CFG4
      generic map(INIT => x"E000")

      port map(A => N_402, B => N_403, C => 
        un14_tx_byte_cntr_0_a2_8_a2_0_5, D => 
        un14_tx_byte_cntr_0_a2_8_a2_0_6, Y => N_554);
    
    \tx_byte_cntr[8]\ : SLE
      port map(D => \tx_byte_cntr_s[8]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \tx_byte_cntr[8]_net_1\);
    
    \tx_byte_cntr[2]\ : SLE
      port map(D => \tx_byte_cntr_s[2]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \tx_byte_cntr[2]_net_1\);
    
    \PreAmble_cntr[6]\ : SLE
      port map(D => \PreAmble_cntr_s[6]\, CLK => BIT_CLK, EN => 
        N_17_i, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PreAmble_cntr[6]_net_1\);
    
    \PreAmble_cntr_RNI4FPH8[5]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \PreAmble_cntr[5]_net_1\, C
         => \PreAmble_cntr_RNIHNV31_Y[6]\, D => GND_net_1, FCI
         => \PreAmble_cntr_cry[4]\, S => \PreAmble_cntr_s[5]\, Y
         => OPEN, FCO => \PreAmble_cntr_cry[5]\);
    
    \TX_SM.un14_tx_byte_cntr_0_a2_8_a2_0_5\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \tx_byte_cntr[10]_net_1\, B => 
        \tx_byte_cntr[8]_net_1\, C => \tx_byte_cntr[7]_net_1\, D
         => \tx_byte_cntr[3]_net_1\, Y => 
        un14_tx_byte_cntr_0_a2_8_a2_0_5);
    
    \PreAmble_cntr_RNI7UJB2[0]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \PreAmble_cntr[0]_net_1\, C
         => \PreAmble_cntr_RNIHNV31_Y[6]\, D => GND_net_1, FCI
         => PreAmble_cntr_cry_cy, S => \PreAmble_cntr_s[0]\, Y
         => OPEN, FCO => \PreAmble_cntr_cry[0]\);
    
    \TX_STATE[7]\ : SLE
      port map(D => \TX_STATE_65\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_STATE[7]_net_1\);
    
    \tx_packet_length_ret_0[10]\ : SLE
      port map(D => \un25_tx_byte_cntr_a_4_i[11]\, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => RESET_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \un25_tx_byte_cntr_a_4[11]\);
    
    \TX_STATE_ns_8_0_.m54_i_0_o2\ : CFG3
      generic map(INIT => x"F8")

      port map(A => \TX_STATE[5]_net_1\, B => un25_tx_byte_cntr, 
        C => \TX_STATE[4]_net_1\, Y => N_471);
    
    \tx_byte_cntr_cry[7]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[7]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[6]_net_1\, S => \tx_byte_cntr_s[7]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[7]_net_1\);
    
    start_tx_FIFO_s : SLE
      port map(D => start_tx_FIFO, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \start_tx_FIFO_s\);
    
    \tx_packet_length[4]\ : SLE
      port map(D => un25_tx_byte_cntr_a_4_axb_3_i, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_packet_length[4]_net_1\);
    
    \TX_SM.un25_tx_byte_cntr_a_4_s_10_RNO\ : CFG4
      generic map(INIT => x"1BFF")

      port map(A => N_81, B => TX_FIFO_DOUT(2), C => 
        \tx_packet_length[10]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => un25_tx_byte_cntr_a_4_s_9_sf);
    
    \TX_STATE_ns_8_0_.m56_i_0_0\ : CFG2
      generic map(INIT => x"B")

      port map(A => un25_tx_byte_cntr, B => \TX_STATE[5]_net_1\, 
        Y => m56_i_0_0);
    
    \tx_byte_cntr[0]\ : SLE
      port map(D => \tx_byte_cntr_s[0]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \tx_byte_cntr[0]_net_1\);
    
    \tx_packet_length[1]\ : SLE
      port map(D => \un25_tx_byte_cntr_a_4_i_i[1]\, CLK => 
        BIT_CLK, EN => un1_byte_clk_en_inv_2_i, ALn => RESET_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \tx_packet_length[1]_net_1\);
    
    \txen_early_cntr_RNI5MOBM[5]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \TX_STATE_RNIAIGV2_Y[7]\, C
         => \txen_early_cntr[5]_net_1\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[4]\, S => \txen_early_cntr_s[5]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[5]\);
    
    \TX_SM.un25_tx_byte_cntr_a_4_cry_7\ : ARI1
      generic map(INIT => x"63B7F")

      port map(A => TX_FIFO_DOUT(0), B => N_81, C => 
        \TX_STATE[5]_net_1\, D => \tx_packet_length[8]_net_1\, 
        FCI => un25_tx_byte_cntr_a_4_cry_6, S => 
        \un25_tx_byte_cntr_a_4_i[8]\, Y => OPEN, FCO => 
        un25_tx_byte_cntr_a_4_cry_7);
    
    \tx_packet_length_ret_0[1]\ : SLE
      port map(D => \un25_tx_byte_cntr_a_4_i[2]\, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => RESET_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \un25_tx_byte_cntr_a_4[2]\);
    
    \tx_byte_cntr_cry[4]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[4]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[3]_net_1\, S => \tx_byte_cntr_s[4]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[4]_net_1\);
    
    \PostAmble_cntr_RNIMPNEJ[10]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => tx_state29_6_RNI9SJ61_Y, C
         => \PostAmble_cntr[10]_net_1\, D => GND_net_1, FCI => 
        \PostAmble_cntr_cry[9]\, S => \PostAmble_cntr_s[10]\, Y
         => OPEN, FCO => \PostAmble_cntr_cry[10]\);
    
    TX_STATE_69 : CFG4
      generic map(INIT => x"11F0")

      port map(A => m56_i_0_0, B => N_554, C => 
        \TX_STATE[3]_net_1\, D => byte_clk_en, Y => \TX_STATE_69\);
    
    \tx_packet_length_RNO[6]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => N_81, B => TX_FIFO_DOUT(6), C => 
        \tx_packet_length[6]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => un25_tx_byte_cntr_a_4_axb_5_i);
    
    \tx_packet_length_RNO[3]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => N_81, B => TX_FIFO_DOUT(3), C => 
        \tx_packet_length[3]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => un25_tx_byte_cntr_a_4_axb_2_i);
    
    \TX_STATE[2]\ : SLE
      port map(D => \TX_STATE_70\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_STATE[2]_net_1\);
    
    \TX_PreAmble\ : SLE
      port map(D => \TX_PreAmble_34\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        TX_PreAmble_net_1);
    
    \tx_packet_length[9]\ : SLE
      port map(D => un25_tx_byte_cntr_a_4_axb_8_i, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_packet_length[9]_net_1\);
    
    \tx_packet_length_ret_0[6]\ : SLE
      port map(D => \un25_tx_byte_cntr_a_4_i[7]\, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => RESET_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \un25_tx_byte_cntr_a_4[7]\);
    
    \PreAmble_cntr_RNIH597[3]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \PreAmble_cntr[3]_net_1\, B => 
        \PreAmble_cntr[4]_net_1\, Y => 
        PreAmble_cntr_0_sqmuxa_0_83_i_o3_0);
    
    \txen_early_cntr_RNIFF8E9[1]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \TX_STATE_RNIAIGV2_Y[7]\, C
         => \txen_early_cntr[1]_net_1\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[0]\, S => \txen_early_cntr_s[1]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[1]\);
    
    \TX_SM.un25_tx_byte_cntr_a_4_s_10\ : CFG2
      generic map(INIT => x"4")

      port map(A => un25_tx_byte_cntr_a_4_cry_8, B => 
        un25_tx_byte_cntr_a_4_s_9_sf, Y => 
        \un25_tx_byte_cntr_a_4_i[11]\);
    
    \TX_SM.un25_tx_byte_cntr_a_4_s_9_931\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => un25_tx_byte_cntr_a_4_cry_8, 
        C => GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => 
        OPEN, Y => OPEN, FCO => un25_tx_byte_cntr_a_4_s_9_931_FCO);
    
    \txen_early_cntr[5]\ : SLE
      port map(D => \txen_early_cntr_s[5]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \txen_early_cntr[5]_net_1\);
    
    \PreAmble_cntr_RNI935A7[4]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \PreAmble_cntr[4]_net_1\, C
         => \PreAmble_cntr_RNIHNV31_Y[6]\, D => GND_net_1, FCI
         => \PreAmble_cntr_cry[3]\, S => \PreAmble_cntr_s[4]\, Y
         => OPEN, FCO => \PreAmble_cntr_cry[4]\);
    
    un1_byte_clk_en_inv_2_0_0_2_RNITD6M : CFG4
      generic map(INIT => x"3331")

      port map(A => \TX_STATE[5]_net_1\, B => 
        \un1_byte_clk_en_inv_2_0_0_2\, C => N_80, D => N_81, Y
         => un1_byte_clk_en_inv_2_i);
    
    TX_PreAmble_34 : CFG3
      generic map(INIT => x"AC")

      port map(A => \TX_STATE[6]_net_1\, B => TX_PreAmble_net_1, 
        C => byte_clk_en, Y => \TX_PreAmble_34\);
    
    \tx_packet_length_ret_0[7]\ : SLE
      port map(D => \un25_tx_byte_cntr_a_4_i[8]\, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => RESET_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \un25_tx_byte_cntr_a_4[8]\);
    
    \tx_byte_cntr[6]\ : SLE
      port map(D => \tx_byte_cntr_s[6]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \tx_byte_cntr[6]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \tx_crc_byte2_en\ : SLE
      port map(D => \TX_STATE[2]_net_1\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        tx_crc_byte2_en);
    
    \tx_packet_length_RNO[0]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => N_81, B => TX_FIFO_DOUT(0), C => 
        \tx_packet_length[0]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => N_12_i);
    
    \tx_byte_cntr_cry[10]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[10]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[9]_net_1\, S => \tx_byte_cntr_s[10]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[10]_net_1\);
    
    \PreAmble_cntr_RNO[6]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \PreAmble_cntr[6]_net_1\, C
         => \PreAmble_cntr_RNIHNV31_Y[6]\, D => GND_net_1, FCI
         => \PreAmble_cntr_cry[5]\, S => \PreAmble_cntr_s[6]\, Y
         => OPEN, FCO => OPEN);
    
    \tx_packet_length[3]\ : SLE
      port map(D => un25_tx_byte_cntr_a_4_axb_2_i, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_packet_length[3]_net_1\);
    
    \PreAmble_cntr[1]\ : SLE
      port map(D => \PreAmble_cntr_s[1]\, CLK => BIT_CLK, EN => 
        N_17_i, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PreAmble_cntr[1]_net_1\);
    
    \PostAmble_cntr[6]\ : SLE
      port map(D => \PostAmble_cntr_s[6]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PostAmble_cntr[6]_net_1\);
    
    \tx_byte_cntr_s[11]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[11]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[10]_net_1\, S => 
        \tx_byte_cntr_s[11]_net_1\, Y => OPEN, FCO => OPEN);
    
    \txen_early_cntr[8]\ : SLE
      port map(D => \txen_early_cntr_s[8]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \txen_early_cntr[8]_net_1\);
    
    \un3_i_0_i[1]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => N_81, B => TX_FIFO_DOUT(1), C => 
        \tx_packet_length[1]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => \un25_tx_byte_cntr_a_4_i_i[1]\);
    
    \tx_byte_cntr[5]\ : SLE
      port map(D => \tx_byte_cntr_s[5]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \tx_byte_cntr[5]_net_1\);
    
    \TX_STATE[0]\ : SLE
      port map(D => \TX_STATE_72\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_STATE[0]_net_1\);
    
    \TX_SM.TX_DataEn_7_iv\ : CFG3
      generic map(INIT => x"8F")

      port map(A => N_163, B => \TX_STATE[6]_net_1\, C => N_213_i, 
        Y => TX_DataEn_7);
    
    \PostAmble_cntr_RNI342U7[3]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => tx_state29_6_RNI9SJ61_Y, C
         => \PostAmble_cntr[3]_net_1\, D => GND_net_1, FCI => 
        \PostAmble_cntr_cry[2]\, S => \PostAmble_cntr_s[3]\, Y
         => OPEN, FCO => \PostAmble_cntr_cry[3]\);
    
    iTX_Enable : SLE
      port map(D => \TX_STATE_i_0[8]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        DRVR_EN_c);
    
    \TX_STATE_ns_8_0_.m38_i_0_a2_0\ : CFG4
      generic map(INIT => x"8000")

      port map(A => m15_e_7, B => m15_e_6, C => 
        \TX_STATE[7]_net_1\, D => m15_e_8, Y => N_362);
    
    \tx_byte_cntr_cry[2]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[2]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[1]_net_1\, S => \tx_byte_cntr_s[2]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[2]_net_1\);
    
    \PreAmble_cntr[3]\ : SLE
      port map(D => \PreAmble_cntr_s[3]\, CLK => BIT_CLK, EN => 
        N_17_i, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PreAmble_cntr[3]_net_1\);
    
    \tx_packet_length_ret_0[4]\ : SLE
      port map(D => \un25_tx_byte_cntr_a_4_i[5]\, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => RESET_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \un25_tx_byte_cntr_a_4[5]\);
    
    \tx_packet_length[10]\ : SLE
      port map(D => un25_tx_byte_cntr_a_4_axb_9_i, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_packet_length[10]_net_1\);
    
    \txen_early_cntr_RNIUP0C61[10]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \TX_STATE_RNIAIGV2_Y[7]\, C
         => \txen_early_cntr[10]_net_1\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[9]\, S => \txen_early_cntr_s[10]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[10]\);
    
    \tx_byte_cntr[11]\ : SLE
      port map(D => \tx_byte_cntr_s[11]_net_1\, CLK => BIT_CLK, 
        EN => byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \tx_byte_cntr[11]_net_1\);
    
    \TX_SM.un25_tx_byte_cntr_a_4_cry_4\ : ARI1
      generic map(INIT => x"637BF")

      port map(A => TX_FIFO_DOUT(5), B => N_81, C => 
        \TX_STATE[5]_net_1\, D => \tx_packet_length[5]_net_1\, 
        FCI => un25_tx_byte_cntr_a_4_cry_3, S => 
        \un25_tx_byte_cntr_a_4_i[5]\, Y => OPEN, FCO => 
        un25_tx_byte_cntr_a_4_cry_4);
    
    \tx_byte_cntr_cry_cy[0]\ : ARI1
      generic map(INIT => x"4EE00")

      port map(A => VCC_net_1, B => \TX_STATE[4]_net_1\, C => 
        \TX_STATE[5]_net_1\, D => GND_net_1, FCI => VCC_net_1, S
         => OPEN, Y => \tx_byte_cntr_cry_cy_Y[0]\, FCO => 
        tx_byte_cntr_cry_cy);
    
    \tx_packet_length[5]\ : SLE
      port map(D => N_49_i, CLK => BIT_CLK, EN => 
        un1_byte_clk_en_inv_2_i, ALn => RESET_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_packet_length[5]_net_1\);
    
    \tx_packet_length_ret_0[0]\ : SLE
      port map(D => un25_tx_byte_cntr_a_4_cry_0_Y, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => RESET_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \un25_tx_byte_cntr_a_4[1]\);
    
    \PreAmble_cntr_RNIFOG26[3]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \PreAmble_cntr[3]_net_1\, C
         => \PreAmble_cntr_RNIHNV31_Y[6]\, D => GND_net_1, FCI
         => \PreAmble_cntr_cry[2]\, S => \PreAmble_cntr_s[3]\, Y
         => OPEN, FCO => \PreAmble_cntr_cry[3]\);
    
    \txen_early_cntr_RNIOG0TF[3]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \TX_STATE_RNIAIGV2_Y[7]\, C
         => \txen_early_cntr[3]_net_1\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[2]\, S => \txen_early_cntr_s[3]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[3]\);
    
    \PostAmble_cntr_RNI6EP9B[5]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => tx_state29_6_RNI9SJ61_Y, C
         => \PostAmble_cntr[5]_net_1\, D => GND_net_1, FCI => 
        \PostAmble_cntr_cry[4]\, S => \PostAmble_cntr_s[5]\, Y
         => OPEN, FCO => \PostAmble_cntr_cry[5]\);
    
    \txen_early_cntr[9]\ : SLE
      port map(D => \txen_early_cntr_s[9]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \txen_early_cntr[9]_net_1\);
    
    \TX_STATE_RNIAIGV2[7]\ : ARI1
      generic map(INIT => x"42AAA")

      port map(A => m15_e_8, B => \TX_STATE[7]_net_1\, C => 
        m15_e_6, D => m15_e_7, FCI => VCC_net_1, S => OPEN, Y => 
        \TX_STATE_RNIAIGV2_Y[7]\, FCO => txen_early_cntr_cry_cy);
    
    \PostAmble_cntr[11]\ : SLE
      port map(D => \PostAmble_cntr_s[11]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PostAmble_cntr[11]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \tx_byte_cntr[4]\ : SLE
      port map(D => \tx_byte_cntr_s[4]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \tx_byte_cntr[4]_net_1\);
    
    \txen_early_cntr[1]\ : SLE
      port map(D => \txen_early_cntr_s[1]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \txen_early_cntr[1]_net_1\);
    
    \tx_byte_cntr_cry[0]\ : ARI1
      generic map(INIT => x"4A800")

      port map(A => VCC_net_1, B => \tx_byte_cntr[0]_net_1\, C
         => \TX_STATE[5]_net_1\, D => \TX_STATE[4]_net_1\, FCI
         => tx_byte_cntr_cry_cy, S => \tx_byte_cntr_s[0]\, Y => 
        OPEN, FCO => \tx_byte_cntr_cry[0]_net_1\);
    
    \TX_STATE_ns_8_0_.m56_i_0_a2_0\ : CFG3
      generic map(INIT => x"40")

      port map(A => \tx_byte_cntr[2]_net_1\, B => 
        \tx_byte_cntr[1]_net_1\, C => \tx_byte_cntr[0]_net_1\, Y
         => N_402);
    
    \TX_SM.un25_tx_byte_cntr_a_4_cry_6\ : ARI1
      generic map(INIT => x"637BF")

      port map(A => TX_FIFO_DOUT(7), B => N_81, C => 
        \TX_STATE[5]_net_1\, D => \tx_packet_length[7]_net_1\, 
        FCI => un25_tx_byte_cntr_a_4_cry_5, S => 
        \un25_tx_byte_cntr_a_4_i[7]\, Y => OPEN, FCO => 
        un25_tx_byte_cntr_a_4_cry_6);
    
    un1_tx_packet_length_0_sqmuxa_0_0_a2 : CFG3
      generic map(INIT => x"C8")

      port map(A => N_81, B => \TX_STATE[5]_net_1\, C => N_80, Y
         => N_513);
    
    \TX_STATE_ns_8_0_.m15_e_6\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \txen_early_cntr[9]_net_1\, B => 
        \txen_early_cntr[8]_net_1\, C => 
        \txen_early_cntr[7]_net_1\, D => 
        \txen_early_cntr[6]_net_1\, Y => m15_e_6);
    
    \txen_early_cntr_RNIBD9931[9]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \TX_STATE_RNIAIGV2_Y[7]\, C
         => \txen_early_cntr[9]_net_1\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[8]\, S => \txen_early_cntr_s[9]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[9]\);
    
    \PostAmble_cntr_RNIDSGLE[7]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => tx_state29_6_RNI9SJ61_Y, C
         => \PostAmble_cntr[7]_net_1\, D => GND_net_1, FCI => 
        \PostAmble_cntr_cry[6]\, S => \PostAmble_cntr_s[7]\, Y
         => OPEN, FCO => \PostAmble_cntr_cry[7]\);
    
    \tx_packet_length_ret_0_RNIOF324[7]\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \tx_byte_cntr[9]_net_1\, B => 
        \un25_tx_byte_cntr_a_4[8]\, C => 
        \un25_tx_byte_cntr_a_4[9]\, D => \tx_byte_cntr[8]_net_1\, 
        FCI => \un25_tx_byte_cntr_1_data_tmp[3]\, S => OPEN, Y
         => OPEN, FCO => \un25_tx_byte_cntr_1_data_tmp[4]\);
    
    \tx_packet_length[8]\ : SLE
      port map(D => N_10_i, CLK => BIT_CLK, EN => 
        un1_byte_clk_en_inv_2_i, ALn => RESET_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_packet_length[8]_net_1\);
    
    \PostAmble_cntr_RNIJG686[2]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => tx_state29_6_RNI9SJ61_Y, C
         => \PostAmble_cntr[2]_net_1\, D => GND_net_1, FCI => 
        \PostAmble_cntr_cry[1]\, S => \PostAmble_cntr_s[2]\, Y
         => OPEN, FCO => \PostAmble_cntr_cry[2]\);
    
    \tx_byte_cntr_cry[1]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[1]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[0]_net_1\, S => \tx_byte_cntr_s[1]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[1]_net_1\);
    
    \TX_DataEn\ : SLE
      port map(D => TX_DataEn_7, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        TX_DataEn);
    
    \tx_byte_cntr[3]\ : SLE
      port map(D => \tx_byte_cntr_s[3]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \tx_byte_cntr[3]_net_1\);
    
    \tx_byte_cntr[7]\ : SLE
      port map(D => \tx_byte_cntr_s[7]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \tx_byte_cntr[7]_net_1\);
    
    \tx_packet_length_ret_0_RNI8D2S[0]\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \tx_packet_length[0]_net_1\, B => 
        \un25_tx_byte_cntr_a_4[1]\, C => \tx_byte_cntr[0]_net_1\, 
        D => \tx_byte_cntr[1]_net_1\, FCI => GND_net_1, S => OPEN, 
        Y => OPEN, FCO => \un25_tx_byte_cntr_1_data_tmp[0]\);
    
    \TX_STATE[8]\ : SLE
      port map(D => \TX_STATE_64\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => RESET_i, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_STATE[8]_net_1\);
    
    \TX_SM.un25_tx_byte_cntr_a_4_cry_8\ : ARI1
      generic map(INIT => x"63B7F")

      port map(A => TX_FIFO_DOUT(1), B => N_81, C => 
        \TX_STATE[5]_net_1\, D => \tx_packet_length[9]_net_1\, 
        FCI => un25_tx_byte_cntr_a_4_cry_7, S => 
        \un25_tx_byte_cntr_a_4_i[9]\, Y => OPEN, FCO => 
        un25_tx_byte_cntr_a_4_cry_8);
    
    \txen_early_cntr_RNIDQ4JP[6]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \TX_STATE_RNIAIGV2_Y[7]\, C
         => \txen_early_cntr[6]_net_1\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[5]\, S => \txen_early_cntr_s[6]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[6]\);
    
    \TX_SM.op_eq.tx_state29_6\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \PostAmble_cntr[9]_net_1\, B => 
        \PostAmble_cntr[8]_net_1\, C => \PostAmble_cntr[7]_net_1\, 
        D => \PostAmble_cntr[6]_net_1\, Y => tx_state29_6);
    
    \txen_early_cntr_RNO[11]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \TX_STATE_RNIAIGV2_Y[7]\, C
         => \txen_early_cntr[11]_net_1\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[10]\, S => \txen_early_cntr_s[11]\, 
        Y => OPEN, FCO => OPEN);
    
    \txen_early_cntr_RNICGS66[0]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \TX_STATE_RNIAIGV2_Y[7]\, C
         => \txen_early_cntr[0]_net_1\, D => GND_net_1, FCI => 
        txen_early_cntr_cry_cy, S => \txen_early_cntr_s[0]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[0]\);
    
    \PreAmble_cntr_RNIU58J3[1]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \PreAmble_cntr[1]_net_1\, C
         => \PreAmble_cntr_RNIHNV31_Y[6]\, D => GND_net_1, FCI
         => \PreAmble_cntr_cry[0]\, S => \PreAmble_cntr_s[1]\, Y
         => OPEN, FCO => \PreAmble_cntr_cry[1]\);
    
    \TX_SM.un25_tx_byte_cntr_a_4_cry_1\ : ARI1
      generic map(INIT => x"637BF")

      port map(A => TX_FIFO_DOUT(2), B => N_81, C => 
        \TX_STATE[5]_net_1\, D => \tx_packet_length[2]_net_1\, 
        FCI => un25_tx_byte_cntr_a_4_cry_0, S => 
        \un25_tx_byte_cntr_a_4_i[2]\, Y => OPEN, FCO => 
        un25_tx_byte_cntr_a_4_cry_1);
    
    \TX_STATE_ns_8_0_.m16_i_0_a2_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => un9_start_tx_fifo_s, B => \TX_STATE[8]_net_1\, 
        Y => N_360);
    
    TX_STATE_68 : CFG4
      generic map(INIT => x"CA0A")

      port map(A => \TX_STATE[4]_net_1\, B => \TX_STATE[6]_net_1\, 
        C => byte_clk_en, D => N_163, Y => \TX_STATE_68\);
    
    \tx_packet_complt\ : SLE
      port map(D => \TX_STATE[0]_net_1\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        tx_packet_complt);
    
    \txen_early_cntr[0]\ : SLE
      port map(D => \txen_early_cntr_s[0]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \txen_early_cntr[0]_net_1\);
    
    \TX_STATE_ns_8_0_.m15_e_7\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \txen_early_cntr[11]_net_1\, B => 
        \txen_early_cntr[10]_net_1\, C => 
        \txen_early_cntr[1]_net_1\, D => 
        \txen_early_cntr[0]_net_1\, Y => m15_e_7);
    
    TX_STATE_71 : CFG4
      generic map(INIT => x"FAD8")

      port map(A => byte_clk_en, B => tx_state29_6_RNI9SJ61_Y, C
         => \TX_STATE[1]_net_1\, D => \TX_STATE[2]_net_1\, Y => 
        \TX_STATE_71\);
    
    \TX_SM.un14_tx_byte_cntr_0_a2_8_a2_0_6_1\ : CFG2
      generic map(INIT => x"1")

      port map(A => \tx_byte_cntr[4]_net_1\, B => 
        \tx_byte_cntr[9]_net_1\, Y => 
        un14_tx_byte_cntr_0_a2_8_a2_0_1_0);
    
    \PreAmble_cntr[2]\ : SLE
      port map(D => \PreAmble_cntr_s[2]\, CLK => BIT_CLK, EN => 
        N_17_i, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PreAmble_cntr[2]_net_1\);
    
    \PostAmble_cntr[8]\ : SLE
      port map(D => \PostAmble_cntr_s[8]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PostAmble_cntr[8]_net_1\);
    
    un1_byte_clk_en_inv_2_0_0_2 : CFG4
      generic map(INIT => x"FFFB")

      port map(A => \TX_STATE[2]_net_1\, B => byte_clk_en, C => 
        \TX_STATE[4]_net_1\, D => \TX_STATE[3]_net_1\, Y => 
        \un1_byte_clk_en_inv_2_0_0_2\);
    
    \TX_STATE_ns_8_0_.m56_i_0_a2_1\ : CFG3
      generic map(INIT => x"02")

      port map(A => \tx_byte_cntr[2]_net_1\, B => 
        \tx_byte_cntr[1]_net_1\, C => \tx_byte_cntr[0]_net_1\, Y
         => N_403);
    
    \tx_packet_length[6]\ : SLE
      port map(D => un25_tx_byte_cntr_a_4_axb_5_i, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_packet_length[6]_net_1\);
    
    \tx_byte_cntr[10]\ : SLE
      port map(D => \tx_byte_cntr_s[10]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \tx_byte_cntr[10]_net_1\);
    
    \TX_STATE_ns_8_0_.m15_e_8\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \txen_early_cntr[5]_net_1\, B => 
        \txen_early_cntr[4]_net_1\, C => 
        \txen_early_cntr[3]_net_1\, D => 
        \txen_early_cntr[2]_net_1\, Y => m15_e_8);
    
    TX_STATE_72 : CFG3
      generic map(INIT => x"AC")

      port map(A => N_511, B => \TX_STATE[0]_net_1\, C => 
        byte_clk_en, Y => \TX_STATE_72\);
    
    \TX_STATE_ns_8_0_.m55_0_a3_0_a2\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_163, B => \TX_STATE[6]_net_1\, Y => 
        TX_DataEn_1_m);
    
    \txen_early_cntr[4]\ : SLE
      port map(D => \txen_early_cntr_s[4]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \txen_early_cntr[4]_net_1\);
    
    \PostAmble_cntr[10]\ : SLE
      port map(D => \PostAmble_cntr_s[10]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PostAmble_cntr[10]_net_1\);
    
    \TX_SM.un14_tx_byte_cntr_0_a2_8_a2_0_6\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \tx_byte_cntr[11]_net_1\, B => 
        \tx_byte_cntr[6]_net_1\, C => \tx_byte_cntr[5]_net_1\, D
         => un14_tx_byte_cntr_0_a2_8_a2_0_1_0, Y => 
        un14_tx_byte_cntr_0_a2_8_a2_0_6);
    
    \PreAmble_cntr_RNIS4IE[0]\ : CFG4
      generic map(INIT => x"BFFF")

      port map(A => \PreAmble_cntr[5]_net_1\, B => 
        \PreAmble_cntr[2]_net_1\, C => \PreAmble_cntr[1]_net_1\, 
        D => \PreAmble_cntr[0]_net_1\, Y => 
        PreAmble_cntr_0_sqmuxa_0_83_i_o3_4);
    
    \tx_crc_byte1_en\ : SLE
      port map(D => \TX_STATE[3]_net_1\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        tx_crc_byte1_en);
    
    \PostAmble_cntr[5]\ : SLE
      port map(D => \PostAmble_cntr_s[5]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PostAmble_cntr[5]_net_1\);
    
    \tx_byte_cntr_cry[5]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[5]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[4]_net_1\, S => \tx_byte_cntr_s[5]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[5]_net_1\);
    
    \PreAmble_cntr_RNI07741[6]\ : CFG4
      generic map(INIT => x"0001")

      port map(A => PreAmble_cntr_0_sqmuxa_0_83_i_o3_0, B => 
        PreAmble_cntr_0_sqmuxa_0_83_i_o3_4, C => 
        \PreAmble_cntr[6]_net_1\, D => TX_FIFO_Empty, Y => N_163);
    
    \TX_SM.op_eq.tx_state29_7\ : CFG4
      generic map(INIT => x"4000")

      port map(A => \PostAmble_cntr[10]_net_1\, B => 
        \PostAmble_cntr[3]_net_1\, C => \PostAmble_cntr[1]_net_1\, 
        D => \PostAmble_cntr[0]_net_1\, Y => tx_state29_7);
    
    \TX_SM.un25_tx_byte_cntr_a_4_s_9\ : ARI1
      generic map(INIT => x"43B7F")

      port map(A => TX_FIFO_DOUT(2), B => N_81, C => 
        \TX_STATE[5]_net_1\, D => \tx_packet_length[10]_net_1\, 
        FCI => un25_tx_byte_cntr_a_4_s_9_931_FCO, S => 
        \un25_tx_byte_cntr_a_4_i[10]\, Y => OPEN, FCO => OPEN);
    
    \PostAmble_cntr[2]\ : SLE
      port map(D => \PostAmble_cntr_s[2]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PostAmble_cntr[2]_net_1\);
    
    TX_STATE_65 : CFG4
      generic map(INIT => x"EEF0")

      port map(A => N_360, B => \TX_STATE_RNIAIGV2_Y[7]\, C => 
        \TX_STATE[7]_net_1\, D => byte_clk_en, Y => \TX_STATE_65\);
    
    \TX_SM.op_eq.tx_state29_8\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \PostAmble_cntr[11]_net_1\, B => 
        \PostAmble_cntr[5]_net_1\, C => \PostAmble_cntr[4]_net_1\, 
        D => \PostAmble_cntr[2]_net_1\, Y => tx_state29_8);
    
    \PostAmble_cntr[1]\ : SLE
      port map(D => \PostAmble_cntr_s[1]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PostAmble_cntr[1]_net_1\);
    
    \tx_packet_length_ret_0[3]\ : SLE
      port map(D => \un25_tx_byte_cntr_a_4_i[4]\, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => RESET_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \un25_tx_byte_cntr_a_4[4]\);
    
    \txen_early_cntr[2]\ : SLE
      port map(D => \txen_early_cntr_s[2]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \txen_early_cntr[2]_net_1\);
    
    \tx_packet_length[2]\ : SLE
      port map(D => un25_tx_byte_cntr_a_4_axb_1_i, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_packet_length[2]_net_1\);
    
    \txen_early_cntr_RNIUIC4J[4]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \TX_STATE_RNIAIGV2_Y[7]\, C
         => \txen_early_cntr[4]_net_1\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[3]\, S => \txen_early_cntr_s[4]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[4]\);
    
    \tx_byte_cntr_cry[6]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[6]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[5]_net_1\, S => \tx_byte_cntr_s[6]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[6]_net_1\);
    
    \txen_early_cntr[7]\ : SLE
      port map(D => \txen_early_cntr_s[7]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \txen_early_cntr[7]_net_1\);
    
    \txen_early_cntr[3]\ : SLE
      port map(D => \txen_early_cntr_s[3]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \txen_early_cntr[3]_net_1\);
    
    \PreAmble_cntr_RNIHNV31[6]\ : ARI1
      generic map(INIT => x"4FE00")

      port map(A => \TX_STATE[6]_net_1\, B => 
        \PreAmble_cntr[6]_net_1\, C => 
        PreAmble_cntr_0_sqmuxa_0_83_i_o3_0, D => 
        PreAmble_cntr_0_sqmuxa_0_83_i_o3_4, FCI => VCC_net_1, S
         => OPEN, Y => \PreAmble_cntr_RNIHNV31_Y[6]\, FCO => 
        PreAmble_cntr_cry_cy);
    
    \PreAmble_cntr[5]\ : SLE
      port map(D => \PreAmble_cntr_s[5]\, CLK => BIT_CLK, EN => 
        N_17_i, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PreAmble_cntr[5]_net_1\);
    
    \TX_SM.un25_tx_byte_cntr_a_4_cry_2\ : ARI1
      generic map(INIT => x"637BF")

      port map(A => TX_FIFO_DOUT(3), B => N_81, C => 
        \TX_STATE[5]_net_1\, D => \tx_packet_length[3]_net_1\, 
        FCI => un25_tx_byte_cntr_a_4_cry_1, S => 
        \un25_tx_byte_cntr_a_4_i[3]\, Y => OPEN, FCO => 
        un25_tx_byte_cntr_a_4_cry_2);
    
    \tx_packet_length_RNO[8]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => N_81, B => TX_FIFO_DOUT(0), C => 
        \tx_packet_length[8]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => N_10_i);
    
    TX_FIFO_rd_en_i : CFG4
      generic map(INIT => x"EC00")

      port map(A => TX_DataEn_1_o, B => 
        un1_tx_packet_length_0_sqmuxa_o, C => TX_PreAmble_net_1, 
        D => byte_clk_en, Y => N_114);
    
    \PostAmble_cntr_RNO[11]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => tx_state29_6_RNI9SJ61_Y, C
         => \PostAmble_cntr[11]_net_1\, D => GND_net_1, FCI => 
        \PostAmble_cntr_cry[10]\, S => \PostAmble_cntr_s[11]\, Y
         => OPEN, FCO => OPEN);
    
    \TX_STATE_RNIC0CR[6]\ : CFG3
      generic map(INIT => x"4C")

      port map(A => TX_FIFO_Empty, B => byte_clk_en, C => 
        \TX_STATE[6]_net_1\, Y => N_17_i);
    
    \PostAmble_cntr_RNIP4LVC[6]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => tx_state29_6_RNI9SJ61_Y, C
         => \PostAmble_cntr[6]_net_1\, D => GND_net_1, FCI => 
        \PostAmble_cntr_cry[5]\, S => \PostAmble_cntr_s[6]\, Y
         => OPEN, FCO => \PostAmble_cntr_cry[6]\);
    
    TX_STATE_70 : CFG3
      generic map(INIT => x"E2")

      port map(A => \TX_STATE[2]_net_1\, B => byte_clk_en, C => 
        \TX_STATE[3]_net_1\, Y => \TX_STATE_70\);
    
    \tx_packet_length_RNO[5]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => N_81, B => TX_FIFO_DOUT(5), C => 
        \tx_packet_length[5]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => N_49_i);
    
    TX_STATE_67 : CFG4
      generic map(INIT => x"EAF0")

      port map(A => N_471, B => N_554, C => \TX_STATE[5]_net_1\, 
        D => byte_clk_en, Y => \TX_STATE_67\);
    
    \tx_packet_length_RNO[7]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => N_81, B => TX_FIFO_DOUT(7), C => 
        \tx_packet_length[7]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => un25_tx_byte_cntr_a_4_axb_6_i);
    
    \PostAmble_cntr[9]\ : SLE
      port map(D => \PostAmble_cntr_s[9]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PostAmble_cntr[9]_net_1\);
    
    \PostAmble_cntr_RNI4UAI4[1]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => tx_state29_6_RNI9SJ61_Y, C
         => \PostAmble_cntr[1]_net_1\, D => GND_net_1, FCI => 
        \PostAmble_cntr_cry[0]\, S => \PostAmble_cntr_s[1]\, Y
         => OPEN, FCO => \PostAmble_cntr_cry[1]\);
    
    \TX_SM.un25_tx_byte_cntr_a_4_cry_3\ : ARI1
      generic map(INIT => x"637BF")

      port map(A => TX_FIFO_DOUT(4), B => N_81, C => 
        \TX_STATE[5]_net_1\, D => \tx_packet_length[4]_net_1\, 
        FCI => un25_tx_byte_cntr_a_4_cry_2, S => 
        \un25_tx_byte_cntr_a_4_i[4]\, Y => OPEN, FCO => 
        un25_tx_byte_cntr_a_4_cry_3);
    
    \tx_packet_length_RNO[9]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => N_81, B => TX_FIFO_DOUT(1), C => 
        \tx_packet_length[9]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => un25_tx_byte_cntr_a_4_axb_8_i);
    
    \PostAmble_cntr_RNIOE81I[9]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => tx_state29_6_RNI9SJ61_Y, C
         => \PostAmble_cntr[9]_net_1\, D => GND_net_1, FCI => 
        \PostAmble_cntr_cry[8]\, S => \PostAmble_cntr_s[9]\, Y
         => OPEN, FCO => \PostAmble_cntr_cry[9]\);
    
    \tx_packet_length_ret_0_RNILDS25[9]\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \tx_byte_cntr[11]_net_1\, B => 
        \un25_tx_byte_cntr_a_4[10]\, C => 
        \un25_tx_byte_cntr_a_4[11]\, D => 
        \tx_byte_cntr[10]_net_1\, FCI => 
        \un25_tx_byte_cntr_1_data_tmp[4]\, S => OPEN, Y => OPEN, 
        FCO => un25_tx_byte_cntr);
    
    \PostAmble_cntr_RNIMCFS2[0]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => tx_state29_6_RNI9SJ61_Y, C
         => \PostAmble_cntr[0]_net_1\, D => GND_net_1, FCI => 
        PostAmble_cntr_cry_cy, S => \PostAmble_cntr_s[0]\, Y => 
        OPEN, FCO => \PostAmble_cntr_cry[0]\);
    
    \tx_byte_cntr[1]\ : SLE
      port map(D => \tx_byte_cntr_s[1]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \tx_byte_cntr[1]_net_1\);
    
    \PostAmble_cntr[4]\ : SLE
      port map(D => \PostAmble_cntr_s[4]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PostAmble_cntr[4]_net_1\);
    
    iTX_FIFO_rd_en_ret_0 : SLE
      port map(D => N_163, CLK => BIT_CLK, EN => byte_clk_en, ALn
         => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => TX_DataEn_1_o);
    
    TX_STATE_64 : CFG4
      generic map(INIT => x"FC70")

      port map(A => un9_start_tx_fifo_s, B => byte_clk_en, C => 
        \TX_STATE[8]_net_1\, D => \TX_STATE[0]_net_1\, Y => 
        \TX_STATE_64\);
    
    \txen_early_cntr_RNI06T101[8]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \TX_STATE_RNIAIGV2_Y[7]\, C
         => \txen_early_cntr[8]_net_1\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[7]\, S => \txen_early_cntr_s[8]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[8]\);
    
    \PreAmble_cntr[4]\ : SLE
      port map(D => \PreAmble_cntr_s[4]\, CLK => BIT_CLK, EN => 
        N_17_i, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PreAmble_cntr[4]_net_1\);
    
    TX_STATE_66 : CFG4
      generic map(INIT => x"BAF0")

      port map(A => N_362, B => N_163, C => \TX_STATE[6]_net_1\, 
        D => byte_clk_en, Y => \TX_STATE_66\);
    
    \PreAmble_cntr[0]\ : SLE
      port map(D => \PreAmble_cntr_s[0]\, CLK => BIT_CLK, EN => 
        N_17_i, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PreAmble_cntr[0]_net_1\);
    
    \tx_packet_length_ret_0_RNIG9IL1[1]\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \tx_byte_cntr[3]_net_1\, B => 
        \un25_tx_byte_cntr_a_4[2]\, C => 
        \un25_tx_byte_cntr_a_4[3]\, D => \tx_byte_cntr[2]_net_1\, 
        FCI => \un25_tx_byte_cntr_1_data_tmp[0]\, S => OPEN, Y
         => OPEN, FCO => \un25_tx_byte_cntr_1_data_tmp[1]\);
    
    \PostAmble_cntr[0]\ : SLE
      port map(D => \PostAmble_cntr_s[0]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PostAmble_cntr[0]_net_1\);
    
    \TX_SM.un25_tx_byte_cntr_a_4_cry_5\ : ARI1
      generic map(INIT => x"637BF")

      port map(A => TX_FIFO_DOUT(6), B => N_81, C => 
        \TX_STATE[5]_net_1\, D => \tx_packet_length[6]_net_1\, 
        FCI => un25_tx_byte_cntr_a_4_cry_4, S => 
        \un25_tx_byte_cntr_a_4_i[6]\, Y => OPEN, FCO => 
        un25_tx_byte_cntr_a_4_cry_5);
    
    iTX_FIFO_rd_en_ret_1_RNO : CFG4
      generic map(INIT => x"EEF0")

      port map(A => N_471, B => N_513, C => 
        un1_tx_packet_length_0_sqmuxa_o, D => byte_clk_en, Y => 
        \iTX_FIFO_rd_en_ret_1_RNO\);
    
    \tx_crc_gen\ : SLE
      port map(D => \tx_byte_cntr_cry_cy_Y[0]\, CLK => BIT_CLK, 
        EN => byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        tx_crc_gen);
    
    iTX_Enable_RNO : CFG1
      generic map(INIT => "01")

      port map(A => \TX_STATE[8]_net_1\, Y => \TX_STATE_i_0[8]\);
    
    \PostAmble_cntr_RNI2LCBG[8]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => tx_state29_6_RNI9SJ61_Y, C
         => \PostAmble_cntr[8]_net_1\, D => GND_net_1, FCI => 
        \PostAmble_cntr_cry[7]\, S => \PostAmble_cntr_s[8]\, Y
         => OPEN, FCO => \PostAmble_cntr_cry[8]\);
    
    \TX_STATE[4]\ : SLE
      port map(D => \TX_STATE_68\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_STATE[4]_net_1\);
    
    \tx_packet_length_ret_0[5]\ : SLE
      port map(D => \un25_tx_byte_cntr_a_4_i[6]\, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => RESET_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \un25_tx_byte_cntr_a_4[6]\);
    
    \tx_packet_length[7]\ : SLE
      port map(D => un25_tx_byte_cntr_a_4_axb_6_i, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_packet_length[7]_net_1\);
    
    \TX_STATE[5]\ : SLE
      port map(D => \TX_STATE_67\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_STATE[5]_net_1\);
    
    \tx_packet_length_RNO[4]\ : CFG4
      generic map(INIT => x"D800")

      port map(A => N_81, B => TX_FIFO_DOUT(4), C => 
        \tx_packet_length[4]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => un25_tx_byte_cntr_a_4_axb_3_i);
    
    \tx_packet_length_ret_0_RNIOQI83[5]\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \tx_byte_cntr[7]_net_1\, B => 
        \un25_tx_byte_cntr_a_4[6]\, C => 
        \un25_tx_byte_cntr_a_4[7]\, D => \tx_byte_cntr[6]_net_1\, 
        FCI => \un25_tx_byte_cntr_1_data_tmp[2]\, S => OPEN, Y
         => OPEN, FCO => \un25_tx_byte_cntr_1_data_tmp[3]\);
    
    \txen_early_cntr[10]\ : SLE
      port map(D => \txen_early_cntr_s[10]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \txen_early_cntr[10]_net_1\);
    
    \TX_STATE[3]\ : SLE
      port map(D => \TX_STATE_69\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_STATE[3]_net_1\);
    
    \tx_packet_length_RNO[10]\ : CFG4
      generic map(INIT => x"E400")

      port map(A => N_81, B => TX_FIFO_DOUT(2), C => 
        \tx_packet_length[10]_net_1\, D => \TX_STATE[5]_net_1\, Y
         => un25_tx_byte_cntr_a_4_axb_9_i);
    
    \tx_byte_cntr_cry[9]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[9]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[8]_net_1\, S => \tx_byte_cntr_s[9]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[9]_net_1\);
    
    \TX_SM.op_eq.tx_state29_6_RNI9SJ61\ : ARI1
      generic map(INIT => x"47F00")

      port map(A => \TX_STATE[1]_net_1\, B => tx_state29_6, C => 
        tx_state29_7, D => tx_state29_8, FCI => VCC_net_1, S => 
        OPEN, Y => tx_state29_6_RNI9SJ61_Y, FCO => 
        PostAmble_cntr_cry_cy);
    
    \PostAmble_cntr_RNIKOTJ9[4]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => tx_state29_6_RNI9SJ61_Y, C
         => \PostAmble_cntr[4]_net_1\, D => GND_net_1, FCI => 
        \PostAmble_cntr_cry[3]\, S => \PostAmble_cntr_s[4]\, Y
         => OPEN, FCO => \PostAmble_cntr_cry[4]\);
    
    TX_IDLE_LINE_DETECTOR : IdleLineDetector_0
      port map(manches_in_dly(1) => manches_in_dly(1), 
        manches_in_dly(0) => manches_in_dly(0), idle_line5 => 
        idle_line5, CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, 
        RESET_i => RESET_i, tx_idle_line => tx_idle_line);
    
    tx_idle_line_s : SLE
      port map(D => tx_idle_line, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \tx_idle_line_s\);
    
    \tx_packet_length[0]\ : SLE
      port map(D => N_12_i, CLK => BIT_CLK, EN => 
        un1_byte_clk_en_inv_2_i, ALn => RESET_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \tx_packet_length[0]_net_1\);
    
    \TX_SM.un9_start_tx_fifo_s\ : CFG2
      generic map(INIT => x"8")

      port map(A => \start_tx_FIFO_s\, B => \tx_idle_line_s\, Y
         => un9_start_tx_fifo_s);
    
    \TX_SM.un14_tx_byte_cntr_0_a2_8_a2\ : CFG3
      generic map(INIT => x"80")

      port map(A => un14_tx_byte_cntr_0_a2_8_a2_0_6, B => N_403, 
        C => un14_tx_byte_cntr_0_a2_8_a2_0_5, Y => N_81);
    
    \txen_early_cntr[6]\ : SLE
      port map(D => \txen_early_cntr_s[6]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \txen_early_cntr[6]_net_1\);
    
    \PostAmble_cntr[7]\ : SLE
      port map(D => \PostAmble_cntr_s[7]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PostAmble_cntr[7]_net_1\);
    
    \tx_packet_length_ret_0[2]\ : SLE
      port map(D => \un25_tx_byte_cntr_a_4_i[3]\, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => RESET_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \un25_tx_byte_cntr_a_4[3]\);
    
    \tx_byte_cntr[9]\ : SLE
      port map(D => \tx_byte_cntr_s[9]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \tx_byte_cntr[9]_net_1\);
    
    \tx_packet_length_ret_0[9]\ : SLE
      port map(D => \un25_tx_byte_cntr_a_4_i[10]\, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => RESET_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \un25_tx_byte_cntr_a_4[10]\);
    
    \tx_byte_cntr_cry[8]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[8]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[7]_net_1\, S => \tx_byte_cntr_s[8]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[8]_net_1\);
    
    \TX_STATE_ns_8_0_.m72_i_i_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \TX_STATE[1]_net_1\, B => tx_state29_7, C => 
        tx_state29_8, D => tx_state29_6, Y => N_511);
    
    \tx_byte_cntr_cry[3]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \tx_byte_cntr_cry_cy_Y[0]\, C
         => \tx_byte_cntr[3]_net_1\, D => GND_net_1, FCI => 
        \tx_byte_cntr_cry[2]_net_1\, S => \tx_byte_cntr_s[3]\, Y
         => OPEN, FCO => \tx_byte_cntr_cry[3]_net_1\);
    
    \PostAmble_cntr[3]\ : SLE
      port map(D => \PostAmble_cntr_s[3]\, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \PostAmble_cntr[3]_net_1\);
    
    un1_TX_STATE_7_i_a2_0_a2_0_a2 : CFG4
      generic map(INIT => x"0001")

      port map(A => \TX_STATE[2]_net_1\, B => \TX_STATE[5]_net_1\, 
        C => \TX_STATE[4]_net_1\, D => \TX_STATE[3]_net_1\, Y => 
        N_213_i);
    
    \txen_early_cntr_RNIMVGQS[7]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \TX_STATE_RNIAIGV2_Y[7]\, C
         => \txen_early_cntr[7]_net_1\, D => GND_net_1, FCI => 
        \txen_early_cntr_cry[6]\, S => \txen_early_cntr_s[7]\, Y
         => OPEN, FCO => \txen_early_cntr_cry[7]\);
    
    \TX_SM.un25_tx_byte_cntr_a_4_cry_0\ : ARI1
      generic map(INIT => x"637BF")

      port map(A => TX_FIFO_DOUT(1), B => N_81, C => 
        \TX_STATE[5]_net_1\, D => \tx_packet_length[1]_net_1\, 
        FCI => GND_net_1, S => OPEN, Y => 
        un25_tx_byte_cntr_a_4_cry_0_Y, FCO => 
        un25_tx_byte_cntr_a_4_cry_0);
    
    \TX_STATE[6]\ : SLE
      port map(D => \TX_STATE_66\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_STATE[6]_net_1\);
    
    \tx_preamble_pat_en\ : SLE
      port map(D => TX_DataEn_1_m, CLK => BIT_CLK, EN => 
        byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        tx_preamble_pat_en);
    
    \TX_STATE[1]\ : SLE
      port map(D => \TX_STATE_71\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_STATE[1]_net_1\);
    
    \TX_SM.un9_tx_byte_cntr_0_a2_0_a2\ : CFG3
      generic map(INIT => x"80")

      port map(A => un14_tx_byte_cntr_0_a2_8_a2_0_6, B => N_402, 
        C => un14_tx_byte_cntr_0_a2_8_a2_0_5, Y => N_80);
    
    \PreAmble_cntr_RNIMESQ4[2]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => \PreAmble_cntr[2]_net_1\, C
         => \PreAmble_cntr_RNIHNV31_Y[6]\, D => GND_net_1, FCI
         => \PreAmble_cntr_cry[1]\, S => \PreAmble_cntr_s[2]\, Y
         => OPEN, FCO => \PreAmble_cntr_cry[2]\);
    
    \tx_packet_length_ret_0_RNI0E2F2[3]\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \tx_byte_cntr[5]_net_1\, B => 
        \un25_tx_byte_cntr_a_4[4]\, C => 
        \un25_tx_byte_cntr_a_4[5]\, D => \tx_byte_cntr[4]_net_1\, 
        FCI => \un25_tx_byte_cntr_1_data_tmp[1]\, S => OPEN, Y
         => OPEN, FCO => \un25_tx_byte_cntr_1_data_tmp[2]\);
    
    \tx_packet_length_ret_0[8]\ : SLE
      port map(D => \un25_tx_byte_cntr_a_4_i[9]\, CLK => BIT_CLK, 
        EN => un1_byte_clk_en_inv_2_i, ALn => RESET_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \un25_tx_byte_cntr_a_4[9]\);
    
    \txen_early_cntr[11]\ : SLE
      port map(D => \txen_early_cntr_s[11]\, CLK => BIT_CLK, EN
         => byte_clk_en, ALn => RESET_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \txen_early_cntr[11]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity ManchesEncoder is

    port( manches_in_dly      : in    std_logic_vector(1 downto 0);
          TX_FIFO_DOUT        : in    std_logic_vector(7 downto 0);
          p2s_data            : out   std_logic_vector(7 downto 0);
          start_tx_FIFO       : in    std_logic;
          TX_FIFO_Empty       : in    std_logic;
          N_114               : out   std_logic;
          idle_line5          : out   std_logic;
          tx_col_detect_en    : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          DRVR_EN_c           : out   std_logic;
          internal_loopback   : in    std_logic;
          external_loopback   : in    std_logic;
          tx_packet_complt    : out   std_logic;
          RESET               : in    std_logic;
          TX_PreAmble         : out   std_logic;
          CommsFPGA_CCC_0_GL1 : in    std_logic;
          byte_clk_en         : in    std_logic;
          BIT_CLK             : in    std_logic;
          RESET_i             : in    std_logic;
          MANCH_OUT_P_c_i     : out   std_logic;
          MANCH_OUT_P_c       : out   std_logic
        );

end ManchesEncoder;

architecture DEF_ARCH of ManchesEncoder is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CRC16_Generator_0
    port( TX_FIFO_DOUT   : in    std_logic_vector(7 downto 0) := (others => 'U');
          tx_crc_data    : out   std_logic_vector(15 downto 0);
          tx_crc_gen     : in    std_logic := 'U';
          byte_clk_en    : in    std_logic := 'U';
          BIT_CLK        : in    std_logic := 'U';
          tx_crc_reset_i : in    std_logic := 'U'
        );
  end component;

  component TX_Collision_Detector
    port( RESET               : in    std_logic := 'U';
          external_loopback   : in    std_logic := 'U';
          internal_loopback   : in    std_logic := 'U';
          DRVR_EN_c           : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          tx_col_detect_en    : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component TX_SM
    port( manches_in_dly      : in    std_logic_vector(1 downto 0) := (others => 'U');
          TX_FIFO_DOUT        : in    std_logic_vector(7 downto 0) := (others => 'U');
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          idle_line5          : out   std_logic;
          N_114               : out   std_logic;
          TX_FIFO_Empty       : in    std_logic := 'U';
          TX_DataEn           : out   std_logic;
          TX_PreAmble         : out   std_logic;
          tx_crc_byte1_en     : out   std_logic;
          tx_crc_byte2_en     : out   std_logic;
          tx_packet_complt    : out   std_logic;
          tx_crc_gen          : out   std_logic;
          start_tx_FIFO       : in    std_logic := 'U';
          DRVR_EN_c           : out   std_logic;
          byte_clk_en         : in    std_logic := 'U';
          tx_preamble_pat_en  : out   std_logic;
          BIT_CLK             : in    std_logic := 'U';
          RESET_i             : in    std_logic := 'U'
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal tx_crc_reset_i, \tx_crc_reset\, \MANCH_OUT_P_c\, 
        \p2s_data[5]_net_1\, VCC_net_1, \p2s_data_9[5]\, 
        GND_net_1, \p2s_data[6]_net_1\, N_296_i, 
        \p2s_data[7]_net_1\, N_295_i, \byte_clk_en_d[0]_net_1\, 
        \TX_PreAmble_d[0]_net_1\, \TX_PreAmble\, 
        \TX_PreAmble_d[1]_net_1\, \p2s_data[0]_net_1\, N_299_i, 
        \p2s_data[1]_net_1\, \p2s_data_9[1]\, \p2s_data[2]_net_1\, 
        N_298_i, \p2s_data[3]_net_1\, \p2s_data_9[3]\, 
        \p2s_data[4]_net_1\, N_297_i, \TX_DataEn_d1\, TX_DataEn, 
        MANCHESTER_OUT_5, tx_preamble_pat_en, N_339, 
        \p2s_data_9_i_0_m2_1_1[0]\, tx_crc_byte1_en, N_487, N_468, 
        \tx_crc_data[8]\, \tx_crc_data[0]\, 
        \p2s_data_9_m2_1_0[1]\, \p2s_data_9_m2[1]\, N_300_1, 
        \tx_crc_data[1]\, \p2s_data_9_m2_1_0[6]\, 
        \p2s_data_9_m2[6]\, \tx_crc_data[6]\, 
        \p2s_data_9_m2_1_0[5]\, \p2s_data_9_m2[5]\, 
        \tx_crc_data[5]\, \p2s_data_9_m2_1_0[7]\, 
        \p2s_data_9_m2[7]\, \tx_crc_data[7]\, 
        \p2s_data_9_m2_1_0[4]\, \p2s_data_9_m2[4]\, 
        \tx_crc_data[4]\, \p2s_data_9_m2_1_0[3]\, 
        \p2s_data_9_m2[3]\, \tx_crc_data[3]\, 
        \p2s_data_9_m2_1_0[2]\, \p2s_data_9_m2[2]\, 
        \tx_crc_data[2]\, un24_tx_dataen, N_460, N_549, 
        \un1_TX_PreAmble_d_i[0]\, tx_crc_byte2_en, 
        \tx_packet_complt\, N_422, N_125, \tx_crc_data[13]\, 
        \tx_crc_data[11]\, \tx_crc_data[9]\, \tx_crc_data[12]\, 
        \tx_crc_data[10]\, \tx_crc_data[15]\, \tx_crc_data[14]\, 
        \DRVR_EN_c\, tx_crc_gen : std_logic;

    for all : CRC16_Generator_0
	Use entity work.CRC16_Generator_0(DEF_ARCH);
    for all : TX_Collision_Detector
	Use entity work.TX_Collision_Detector(DEF_ARCH);
    for all : TX_SM
	Use entity work.TX_SM(DEF_ARCH);
begin 

    p2s_data(7) <= \p2s_data[7]_net_1\;
    p2s_data(6) <= \p2s_data[6]_net_1\;
    p2s_data(5) <= \p2s_data[5]_net_1\;
    p2s_data(4) <= \p2s_data[4]_net_1\;
    p2s_data(3) <= \p2s_data[3]_net_1\;
    p2s_data(2) <= \p2s_data[2]_net_1\;
    p2s_data(1) <= \p2s_data[1]_net_1\;
    p2s_data(0) <= \p2s_data[0]_net_1\;
    DRVR_EN_c <= \DRVR_EN_c\;
    tx_packet_complt <= \tx_packet_complt\;
    TX_PreAmble <= \TX_PreAmble\;
    MANCH_OUT_P_c <= \MANCH_OUT_P_c\;

    \byte_clk_en_d[0]\ : SLE
      port map(D => byte_clk_en, CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \byte_clk_en_d[0]_net_1\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_m2[3]\ : CFG4
      generic map(INIT => x"AAC5")

      port map(A => \p2s_data_9_m2_1_0[3]\, B => TX_FIFO_DOUT(3), 
        C => N_487, D => N_339, Y => \p2s_data_9_m2[3]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_m2_1_0[4]\ : CFG4
      generic map(INIT => x"2075")

      port map(A => N_339, B => N_300_1, C => \p2s_data[3]_net_1\, 
        D => \tx_crc_data[4]\, Y => \p2s_data_9_m2_1_0[4]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_0_a2_3[1]\ : CFG4
      generic map(INIT => x"0020")

      port map(A => TX_DataEn, B => N_460, C => 
        \byte_clk_en_d[0]_net_1\, D => tx_preamble_pat_en, Y => 
        N_422);
    
    \TX_PreAmble_d[0]\ : SLE
      port map(D => \TX_PreAmble\, CLK => CommsFPGA_CCC_0_GL1, EN
         => VCC_net_1, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_PreAmble_d[0]_net_1\);
    
    \un1_TX_PreAmble_d_0_o2_0_o2[0]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => N_549, B => \TX_PreAmble\, C => 
        tx_preamble_pat_en, Y => \un1_TX_PreAmble_d_i[0]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_m2_1_0[5]\ : CFG4
      generic map(INIT => x"2075")

      port map(A => N_339, B => N_300_1, C => \p2s_data[4]_net_1\, 
        D => \tx_crc_data[5]\, Y => \p2s_data_9_m2_1_0[5]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_0_0[1]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => N_422, B => \tx_crc_data[9]\, C => 
        \p2s_data_9_m2[1]\, D => N_125, Y => \p2s_data_9[1]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_m2[4]\ : CFG4
      generic map(INIT => x"AAC5")

      port map(A => \p2s_data_9_m2_1_0[4]\, B => TX_FIFO_DOUT(4), 
        C => N_487, D => N_339, Y => \p2s_data_9_m2[4]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_0_o2_0[1]\ : CFG2
      generic map(INIT => x"D")

      port map(A => tx_crc_byte1_en, B => 
        \TX_PreAmble_d[1]_net_1\, Y => N_460);
    
    \p2s_data[0]\ : SLE
      port map(D => N_299_i, CLK => BIT_CLK, EN => VCC_net_1, ALn
         => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \p2s_data[0]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \p2s_data[6]\ : SLE
      port map(D => N_296_i, CLK => BIT_CLK, EN => VCC_net_1, ALn
         => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \p2s_data[6]_net_1\);
    
    \MAN_OUT_DATA_PROC.un24_tx_dataen\ : CFG2
      generic map(INIT => x"E")

      port map(A => TX_DataEn, B => \TX_DataEn_d1\, Y => 
        un24_tx_dataen);
    
    tx_crc_reset_RNI5CLE : CLKINT
      port map(A => \tx_crc_reset\, Y => tx_crc_reset_i);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_i_0_m2[0]\ : CFG4
      generic map(INIT => x"7455")

      port map(A => \p2s_data_9_i_0_m2_1_1[0]\, B => 
        tx_crc_byte1_en, C => TX_FIFO_DOUT(0), D => N_487, Y => 
        N_468);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_0_0[3]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => N_422, B => \tx_crc_data[11]\, C => 
        \p2s_data_9_m2[3]\, D => N_125, Y => \p2s_data_9[3]\);
    
    TX_CRC_GEN_INST : CRC16_Generator_0
      port map(TX_FIFO_DOUT(7) => TX_FIFO_DOUT(7), 
        TX_FIFO_DOUT(6) => TX_FIFO_DOUT(6), TX_FIFO_DOUT(5) => 
        TX_FIFO_DOUT(5), TX_FIFO_DOUT(4) => TX_FIFO_DOUT(4), 
        TX_FIFO_DOUT(3) => TX_FIFO_DOUT(3), TX_FIFO_DOUT(2) => 
        TX_FIFO_DOUT(2), TX_FIFO_DOUT(1) => TX_FIFO_DOUT(1), 
        TX_FIFO_DOUT(0) => TX_FIFO_DOUT(0), tx_crc_data(15) => 
        \tx_crc_data[15]\, tx_crc_data(14) => \tx_crc_data[14]\, 
        tx_crc_data(13) => \tx_crc_data[13]\, tx_crc_data(12) => 
        \tx_crc_data[12]\, tx_crc_data(11) => \tx_crc_data[11]\, 
        tx_crc_data(10) => \tx_crc_data[10]\, tx_crc_data(9) => 
        \tx_crc_data[9]\, tx_crc_data(8) => \tx_crc_data[8]\, 
        tx_crc_data(7) => \tx_crc_data[7]\, tx_crc_data(6) => 
        \tx_crc_data[6]\, tx_crc_data(5) => \tx_crc_data[5]\, 
        tx_crc_data(4) => \tx_crc_data[4]\, tx_crc_data(3) => 
        \tx_crc_data[3]\, tx_crc_data(2) => \tx_crc_data[2]\, 
        tx_crc_data(1) => \tx_crc_data[1]\, tx_crc_data(0) => 
        \tx_crc_data[0]\, tx_crc_gen => tx_crc_gen, byte_clk_en
         => byte_clk_en, BIT_CLK => BIT_CLK, tx_crc_reset_i => 
        tx_crc_reset_i);
    
    TX_COLLISION_DETECTOR_INST : TX_Collision_Detector
      port map(RESET => RESET, external_loopback => 
        external_loopback, internal_loopback => internal_loopback, 
        DRVR_EN_c => \DRVR_EN_c\, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, tx_col_detect_en => tx_col_detect_en);
    
    \p2s_data[2]\ : SLE
      port map(D => N_298_i, CLK => BIT_CLK, EN => VCC_net_1, ALn
         => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \p2s_data[2]_net_1\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_m2[7]\ : CFG4
      generic map(INIT => x"AAC5")

      port map(A => \p2s_data_9_m2_1_0[7]\, B => TX_FIFO_DOUT(7), 
        C => N_487, D => N_339, Y => \p2s_data_9_m2[7]\);
    
    \MAN_OUT_DATA_PROC.MANCHESTER_OUT_5_u\ : CFG4
      generic map(INIT => x"36CC")

      port map(A => un24_tx_dataen, B => \p2s_data[7]_net_1\, C
         => \un1_TX_PreAmble_d_i[0]\, D => BIT_CLK, Y => 
        MANCHESTER_OUT_5);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_ss0_i_0_a2_1\ : CFG3
      generic map(INIT => x"40")

      port map(A => tx_crc_byte2_en, B => 
        \byte_clk_en_d[0]_net_1\, C => TX_DataEn, Y => N_487);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_i_0_m2_1_1[0]\ : CFG3
      generic map(INIT => x"27")

      port map(A => tx_crc_byte1_en, B => \tx_crc_data[8]\, C => 
        \tx_crc_data[0]\, Y => \p2s_data_9_i_0_m2_1_1[0]\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \PARALLEL_2_SERIAL_PROC.un5_tx_dataen_i_o2_0_o2\ : CFG4
      generic map(INIT => x"73FF")

      port map(A => tx_preamble_pat_en, B => TX_DataEn, C => 
        \TX_PreAmble_d[1]_net_1\, D => \byte_clk_en_d[0]_net_1\, 
        Y => N_339);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_m2_1_0[2]\ : CFG4
      generic map(INIT => x"2075")

      port map(A => N_339, B => N_300_1, C => \p2s_data[1]_net_1\, 
        D => \tx_crc_data[2]\, Y => \p2s_data_9_m2_1_0[2]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_m2_1_0[6]\ : CFG4
      generic map(INIT => x"2075")

      port map(A => N_339, B => N_300_1, C => \p2s_data[5]_net_1\, 
        D => \tx_crc_data[6]\, Y => \p2s_data_9_m2_1_0[6]\);
    
    \p2s_data_RNO[6]\ : CFG4
      generic map(INIT => x"D0DD")

      port map(A => N_422, B => \tx_crc_data[14]\, C => 
        \p2s_data_9_m2[6]\, D => N_125, Y => N_296_i);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_m2_1_0[1]\ : CFG4
      generic map(INIT => x"2705")

      port map(A => N_339, B => N_300_1, C => \tx_crc_data[1]\, D
         => \p2s_data[0]_net_1\, Y => \p2s_data_9_m2_1_0[1]\);
    
    \p2s_data[4]\ : SLE
      port map(D => N_297_i, CLK => BIT_CLK, EN => VCC_net_1, ALn
         => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \p2s_data[4]_net_1\);
    
    TRANSMIT_SM : TX_SM
      port map(manches_in_dly(1) => manches_in_dly(1), 
        manches_in_dly(0) => manches_in_dly(0), TX_FIFO_DOUT(7)
         => TX_FIFO_DOUT(7), TX_FIFO_DOUT(6) => TX_FIFO_DOUT(6), 
        TX_FIFO_DOUT(5) => TX_FIFO_DOUT(5), TX_FIFO_DOUT(4) => 
        TX_FIFO_DOUT(4), TX_FIFO_DOUT(3) => TX_FIFO_DOUT(3), 
        TX_FIFO_DOUT(2) => TX_FIFO_DOUT(2), TX_FIFO_DOUT(1) => 
        TX_FIFO_DOUT(1), TX_FIFO_DOUT(0) => TX_FIFO_DOUT(0), 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, idle_line5
         => idle_line5, N_114 => N_114, TX_FIFO_Empty => 
        TX_FIFO_Empty, TX_DataEn => TX_DataEn, TX_PreAmble => 
        \TX_PreAmble\, tx_crc_byte1_en => tx_crc_byte1_en, 
        tx_crc_byte2_en => tx_crc_byte2_en, tx_packet_complt => 
        \tx_packet_complt\, tx_crc_gen => tx_crc_gen, 
        start_tx_FIFO => start_tx_FIFO, DRVR_EN_c => \DRVR_EN_c\, 
        byte_clk_en => byte_clk_en, tx_preamble_pat_en => 
        tx_preamble_pat_en, BIT_CLK => BIT_CLK, RESET_i => 
        RESET_i);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_m2_1_0[7]\ : CFG4
      generic map(INIT => x"2705")

      port map(A => N_339, B => N_300_1, C => \tx_crc_data[7]\, D
         => \p2s_data[6]_net_1\, Y => \p2s_data_9_m2_1_0[7]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_m2[2]\ : CFG4
      generic map(INIT => x"AAC5")

      port map(A => \p2s_data_9_m2_1_0[2]\, B => TX_FIFO_DOUT(2), 
        C => N_487, D => N_339, Y => \p2s_data_9_m2[2]\);
    
    \p2s_data_RNO[2]\ : CFG4
      generic map(INIT => x"D0DD")

      port map(A => N_422, B => \tx_crc_data[10]\, C => 
        \p2s_data_9_m2[2]\, D => N_125, Y => N_298_i);
    
    \p2s_data_RNO[4]\ : CFG4
      generic map(INIT => x"D0DD")

      port map(A => N_422, B => \tx_crc_data[12]\, C => 
        \p2s_data_9_m2[4]\, D => N_125, Y => N_297_i);
    
    \p2s_data[1]\ : SLE
      port map(D => \p2s_data_9[1]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \p2s_data[1]_net_1\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_m2_1_0[3]\ : CFG4
      generic map(INIT => x"2075")

      port map(A => N_339, B => N_300_1, C => \p2s_data[2]_net_1\, 
        D => \tx_crc_data[3]\, Y => \p2s_data_9_m2_1_0[3]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_0_0[5]\ : CFG4
      generic map(INIT => x"F888")

      port map(A => N_422, B => \tx_crc_data[13]\, C => 
        \p2s_data_9_m2[5]\, D => N_125, Y => \p2s_data_9[5]\);
    
    \p2s_data_RNO[0]\ : CFG3
      generic map(INIT => x"32")

      port map(A => tx_preamble_pat_en, B => N_339, C => N_468, Y
         => N_299_i);
    
    \p2s_data[3]\ : SLE
      port map(D => \p2s_data_9[3]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \p2s_data[3]_net_1\);
    
    MANCHESTER_OUT : SLE
      port map(D => MANCHESTER_OUT_5, CLK => CommsFPGA_CCC_0_GL1, 
        EN => VCC_net_1, ALn => RESET_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \MANCH_OUT_P_c\);
    
    \TX_PreAmble_d[1]\ : SLE
      port map(D => \TX_PreAmble_d[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL1, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \TX_PreAmble_d[1]_net_1\);
    
    MANCHESTER_OUT_RNI19ND : CFG1
      generic map(INIT => "01")

      port map(A => \MANCH_OUT_P_c\, Y => MANCH_OUT_P_c_i);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_m2[5]\ : CFG4
      generic map(INIT => x"AAC5")

      port map(A => \p2s_data_9_m2_1_0[5]\, B => TX_FIFO_DOUT(5), 
        C => N_487, D => N_339, Y => \p2s_data_9_m2[5]\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_ss0_i_0_1\ : CFG4
      generic map(INIT => x"AB03")

      port map(A => \byte_clk_en_d[0]_net_1\, B => \TX_PreAmble\, 
        C => TX_DataEn, D => N_549, Y => N_300_1);
    
    \p2s_data[5]\ : SLE
      port map(D => \p2s_data_9[5]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => RESET_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \p2s_data[5]_net_1\);
    
    TX_DataEn_d1 : SLE
      port map(D => TX_DataEn, CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \TX_DataEn_d1\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_ss0_i_0_a2_2\ : CFG2
      generic map(INIT => x"4")

      port map(A => tx_preamble_pat_en, B => 
        \TX_PreAmble_d[1]_net_1\, Y => N_549);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_0_0_o2[1]\ : CFG4
      generic map(INIT => x"5FDF")

      port map(A => TX_DataEn, B => N_460, C => 
        \byte_clk_en_d[0]_net_1\, D => tx_preamble_pat_en, Y => 
        N_125);
    
    tx_crc_reset : CFG2
      generic map(INIT => x"1")

      port map(A => RESET, B => \tx_packet_complt\, Y => 
        \tx_crc_reset\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_m2[1]\ : CFG4
      generic map(INIT => x"AAC5")

      port map(A => \p2s_data_9_m2_1_0[1]\, B => TX_FIFO_DOUT(1), 
        C => N_487, D => N_339, Y => \p2s_data_9_m2[1]\);
    
    \p2s_data_RNO[7]\ : CFG4
      generic map(INIT => x"D0DD")

      port map(A => N_422, B => \tx_crc_data[15]\, C => 
        \p2s_data_9_m2[7]\, D => N_125, Y => N_295_i);
    
    \p2s_data[7]\ : SLE
      port map(D => N_295_i, CLK => BIT_CLK, EN => VCC_net_1, ALn
         => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \p2s_data[7]_net_1\);
    
    \PARALLEL_2_SERIAL_PROC.p2s_data_9_m2[6]\ : CFG4
      generic map(INIT => x"AAC5")

      port map(A => \p2s_data_9_m2_1_0[6]\, B => TX_FIFO_DOUT(6), 
        C => N_487, D => N_339, Y => \p2s_data_9_m2[6]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity IdleLineDetector_1 is

    port( idle_line5          : in    std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          RESET_i             : in    std_logic;
          idle_line           : out   std_logic
        );

end IdleLineDetector_1;

architecture DEF_ARCH of IdleLineDetector_1 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \idle_line_cntr_0_sqmuxa\, GND_net_1, 
        \idle_line_cntr[0]_net_1\, \idle_line_cntr_s[0]\, 
        \idle_line_cntr[1]_net_1\, \idle_line_cntr_s[1]\, 
        \idle_line_cntr[2]_net_1\, \idle_line_cntr_s[2]\, 
        \idle_line_cntr[3]_net_1\, \idle_line_cntr_s[3]\, 
        \idle_line_cntr[4]_net_1\, \idle_line_cntr_s[4]\, 
        \idle_line_cntr[5]_net_1\, \idle_line_cntr_s[5]\, 
        \idle_line_cntr[6]_net_1\, \idle_line_cntr_s[6]\, 
        \idle_line_cntr[7]_net_1\, \idle_line_cntr_s[7]\, 
        \idle_line_cntr[8]_net_1\, \idle_line_cntr_s[8]\, 
        \idle_line_cntr[9]_net_1\, \idle_line_cntr_s[9]\, 
        \idle_line_cntr[10]_net_1\, \idle_line_cntr_s[10]\, 
        \idle_line_cntr[11]_net_1\, \idle_line_cntr_s[11]\, 
        \idle_line_cntr[12]_net_1\, \idle_line_cntr_s[12]\, 
        \idle_line_cntr[13]_net_1\, \idle_line_cntr_s[13]\, 
        \idle_line_cntr[14]_net_1\, \idle_line_cntr_s[14]\, 
        \idle_line_cntr[15]_net_1\, \idle_line_cntr_s[15]\, 
        idle_line_cntr_cry_cy, un5_manches_in_dly_9_RNINM8S_Y, 
        un5_manches_in_dly_9, un5_manches_in_dly_10, 
        un5_manches_in_dly_11, \idle_line_cntr_cry[0]\, 
        \idle_line_cntr_cry[1]\, \idle_line_cntr_cry[2]\, 
        \idle_line_cntr_cry[3]\, \idle_line_cntr_cry[4]\, 
        \idle_line_cntr_cry[5]\, \idle_line_cntr_cry[6]\, 
        \idle_line_cntr_cry[7]\, \idle_line_cntr_cry[8]\, 
        \idle_line_cntr_cry[9]\, \idle_line_cntr_cry[10]\, 
        \idle_line_cntr_cry[11]\, \idle_line_cntr_cry[12]\, 
        \idle_line_cntr_cry[13]\, \idle_line_cntr_cry[14]\, 
        un5_manches_in_dly_8 : std_logic;

begin 


    \idle_line\ : SLE
      port map(D => \idle_line_cntr_0_sqmuxa\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => idle_line);
    
    \IDLE_LINE_DETECT_PROC.un5_manches_in_dly_11\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \idle_line_cntr[11]_net_1\, B => 
        \idle_line_cntr[8]_net_1\, C => \idle_line_cntr[7]_net_1\, 
        D => un5_manches_in_dly_8, Y => un5_manches_in_dly_11);
    
    \idle_line_cntr_RNILB687[6]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[6]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[5]\, S => \idle_line_cntr_s[6]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[6]\);
    
    idle_line_cntr_0_sqmuxa : CFG4
      generic map(INIT => x"0800")

      port map(A => un5_manches_in_dly_10, B => 
        un5_manches_in_dly_9, C => idle_line5, D => 
        un5_manches_in_dly_11, Y => \idle_line_cntr_0_sqmuxa\);
    
    \idle_line_cntr_RNIN3V8E[12]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[12]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[11]\, S => \idle_line_cntr_s[12]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[12]\);
    
    \idle_line_cntr_RNI24F29[8]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[8]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[7]\, S => \idle_line_cntr_s[8]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[8]\);
    
    \idle_line_cntr[4]\ : SLE
      port map(D => \idle_line_cntr_s[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[4]_net_1\);
    
    \idle_line_cntr[14]\ : SLE
      port map(D => \idle_line_cntr_s[14]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[14]_net_1\);
    
    \idle_line_cntr_RNIM0HM2[1]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[1]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[0]\, S => \idle_line_cntr_s[1]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[1]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \IDLE_LINE_DETECT_PROC.un5_manches_in_dly_9\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \idle_line_cntr[10]_net_1\, B => 
        \idle_line_cntr[9]_net_1\, C => \idle_line_cntr[2]_net_1\, 
        D => \idle_line_cntr[1]_net_1\, Y => un5_manches_in_dly_9);
    
    \IDLE_LINE_DETECT_PROC.un5_manches_in_dly_10\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \idle_line_cntr[6]_net_1\, B => 
        \idle_line_cntr[5]_net_1\, C => \idle_line_cntr[4]_net_1\, 
        D => \idle_line_cntr[3]_net_1\, Y => 
        un5_manches_in_dly_10);
    
    \idle_line_cntr_RNICNTD5[4]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[4]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[3]\, S => \idle_line_cntr_s[4]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[4]\);
    
    \idle_line_cntr[9]\ : SLE
      port map(D => \idle_line_cntr_s[9]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[9]_net_1\);
    
    \idle_line_cntr[8]\ : SLE
      port map(D => \idle_line_cntr_s[8]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[8]_net_1\);
    
    \idle_line_cntr[7]\ : SLE
      port map(D => \idle_line_cntr_s[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[7]_net_1\);
    
    \idle_line_cntr[15]\ : SLE
      port map(D => \idle_line_cntr_s[15]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[15]_net_1\);
    
    \idle_line_cntr[11]\ : SLE
      port map(D => \idle_line_cntr_s[11]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[11]_net_1\);
    
    \idle_line_cntr[10]\ : SLE
      port map(D => \idle_line_cntr_s[10]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[10]_net_1\);
    
    \idle_line_cntr[1]\ : SLE
      port map(D => \idle_line_cntr_s[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[1]_net_1\);
    
    \IDLE_LINE_DETECT_PROC.un5_manches_in_dly_8\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \idle_line_cntr[15]_net_1\, B => 
        \idle_line_cntr[14]_net_1\, C => 
        \idle_line_cntr[13]_net_1\, D => 
        \idle_line_cntr[12]_net_1\, Y => un5_manches_in_dly_8);
    
    \idle_line_cntr_RNO[15]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[15]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[14]\, S => \idle_line_cntr_s[15]\, Y
         => OPEN, FCO => OPEN);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \idle_line_cntr_RNI77LJ3[2]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[2]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[1]\, S => \idle_line_cntr_s[2]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[2]\);
    
    \IDLE_LINE_DETECT_PROC.un5_manches_in_dly_9_RNINM8S\ : ARI1
      generic map(INIT => x"4007F")

      port map(A => idle_line5, B => un5_manches_in_dly_9, C => 
        un5_manches_in_dly_10, D => un5_manches_in_dly_11, FCI
         => VCC_net_1, S => OPEN, Y => 
        un5_manches_in_dly_9_RNINM8S_Y, FCO => 
        idle_line_cntr_cry_cy);
    
    \idle_line_cntr_RNI6RCP1[0]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[0]_net_1\, D => GND_net_1, FCI => 
        idle_line_cntr_cry_cy, S => \idle_line_cntr_s[0]\, Y => 
        OPEN, FCO => \idle_line_cntr_cry[0]\);
    
    \idle_line_cntr_RNILED0D[11]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[11]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[10]\, S => \idle_line_cntr_s[11]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[11]\);
    
    \idle_line_cntr[6]\ : SLE
      port map(D => \idle_line_cntr_s[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[6]_net_1\);
    
    \idle_line_cntr_RNIPEPG4[3]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[3]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[2]\, S => \idle_line_cntr_s[3]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[3]\);
    
    \idle_line_cntr[13]\ : SLE
      port map(D => \idle_line_cntr_s[13]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[13]_net_1\);
    
    \idle_line_cntr[0]\ : SLE
      port map(D => \idle_line_cntr_s[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[0]_net_1\);
    
    \idle_line_cntr_RNIUG2QG[14]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[14]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[13]\, S => \idle_line_cntr_s[14]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[14]\);
    
    \idle_line_cntr_RNI012B6[5]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[5]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[4]\, S => \idle_line_cntr_s[5]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[5]\);
    
    \idle_line_cntr[12]\ : SLE
      port map(D => \idle_line_cntr_s[12]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[12]_net_1\);
    
    \idle_line_cntr[3]\ : SLE
      port map(D => \idle_line_cntr_s[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[3]_net_1\);
    
    \idle_line_cntr_RNINSE7A[9]\ : ARI1
      generic map(INIT => x"4D800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[9]_net_1\, D => \idle_line_cntr_0_sqmuxa\, 
        FCI => \idle_line_cntr_cry[8]\, S => 
        \idle_line_cntr_s[9]\, Y => OPEN, FCO => 
        \idle_line_cntr_cry[9]\);
    
    \idle_line_cntr_RNIKQRNB[10]\ : ARI1
      generic map(INIT => x"4D800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[10]_net_1\, D => 
        \idle_line_cntr_0_sqmuxa\, FCI => \idle_line_cntr_cry[9]\, 
        S => \idle_line_cntr_s[10]\, Y => OPEN, FCO => 
        \idle_line_cntr_cry[10]\);
    
    \idle_line_cntr_RNIQPGHF[13]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[13]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[12]\, S => \idle_line_cntr_s[13]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[13]\);
    
    \idle_line_cntr[5]\ : SLE
      port map(D => \idle_line_cntr_s[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[5]_net_1\);
    
    \idle_line_cntr_RNIBNA58[7]\ : ARI1
      generic map(INIT => x"48800")

      port map(A => VCC_net_1, B => 
        un5_manches_in_dly_9_RNINM8S_Y, C => 
        \idle_line_cntr[7]_net_1\, D => GND_net_1, FCI => 
        \idle_line_cntr_cry[6]\, S => \idle_line_cntr_s[7]\, Y
         => OPEN, FCO => \idle_line_cntr_cry[7]\);
    
    \idle_line_cntr[2]\ : SLE
      port map(D => \idle_line_cntr_s[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \idle_line_cntr[2]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity ManchesDecoder_Adapter is

    port( clkdiv              : out   std_logic_vector(3 downto 0);
          RX_FIFO_DIN         : out   std_logic_vector(7 downto 0);
          manches_in_dly      : out   std_logic_vector(1 downto 0);
          idle_line5          : in    std_logic;
          RESET               : in    std_logic;
          MANCHESTER_IN_c     : in    std_logic;
          MANCH_OUT_P_c       : in    std_logic;
          internal_loopback   : in    std_logic;
          rx_packet_end_all   : in    std_logic;
          idle_line           : out   std_logic;
          irx_center_sample   : out   std_logic;
          sampler_clk1x_en    : out   std_logic;
          iNRZ_data           : out   std_logic;
          clk1x_enable        : in    std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          RESET_i             : in    std_logic
        );

end ManchesDecoder_Adapter;

architecture DEF_ARCH of ManchesDecoder_Adapter is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component IdleLineDetector_1
    port( idle_line5          : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          RESET_i             : in    std_logic := 'U';
          idle_line           : out   std_logic
        );
  end component;

    signal \clock_adjust\, clock_adjust_i, \manches_in_dly[0]\, 
        GND_net_1, \un1_manches_in[0]_net_1\, VCC_net_1, 
        \manches_in_dly[1]\, \decoder_Transition_d[0]_net_1\, 
        un2_rst_i, \decoder_Transition\, 
        \decoder_Transition_d[1]_net_1\, 
        \decoder_Transition_d[2]_net_1\, \RX_FIFO_DIN[0]\, 
        iNRZ_data_net_1, \sampler_clk1x_en\, \RX_FIFO_DIN[1]\, 
        \RX_FIFO_DIN[2]\, \RX_FIFO_DIN[3]\, \RX_FIFO_DIN[4]\, 
        \RX_FIFO_DIN[5]\, \RX_FIFO_DIN[6]\, 
        \decoder_ShiftReg[0]_net_1\, \clkdiv[3]_net_1\, 
        \manches_ShiftReg[0]_net_1\, un18_rst_i, iNRZ_data_1, 
        irx_center_sample_net_1, isampler_clk1x_en_1, 
        decoder_Transition_1, \manches_Transition\, 
        manches_Transition_1, un16_irx_center_sample, 
        un16_clk1x_enable, \clkdiv[0]_net_1\, \clkdiv_3[0]_net_1\, 
        \clkdiv[1]_net_1\, \clkdiv_3[1]_net_1\, \clkdiv[2]_net_1\, 
        \clkdiv_3[2]_net_1\, \clkdiv_3[3]_net_1\, \idle_line\, 
        \un1_iidle_line\, CO1 : std_logic;

    for all : IdleLineDetector_1
	Use entity work.IdleLineDetector_1(DEF_ARCH);
begin 

    clkdiv(3) <= \clkdiv[3]_net_1\;
    clkdiv(2) <= \clkdiv[2]_net_1\;
    clkdiv(1) <= \clkdiv[1]_net_1\;
    clkdiv(0) <= \clkdiv[0]_net_1\;
    RX_FIFO_DIN(6) <= \RX_FIFO_DIN[6]\;
    RX_FIFO_DIN(5) <= \RX_FIFO_DIN[5]\;
    RX_FIFO_DIN(4) <= \RX_FIFO_DIN[4]\;
    RX_FIFO_DIN(3) <= \RX_FIFO_DIN[3]\;
    RX_FIFO_DIN(2) <= \RX_FIFO_DIN[2]\;
    RX_FIFO_DIN(1) <= \RX_FIFO_DIN[1]\;
    RX_FIFO_DIN(0) <= \RX_FIFO_DIN[0]\;
    manches_in_dly(1) <= \manches_in_dly[1]\;
    manches_in_dly(0) <= \manches_in_dly[0]\;
    idle_line <= \idle_line\;
    irx_center_sample <= irx_center_sample_net_1;
    sampler_clk1x_en <= \sampler_clk1x_en\;
    iNRZ_data <= iNRZ_data_net_1;

    \s2p_data[2]\ : SLE
      port map(D => \RX_FIFO_DIN[1]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => \sampler_clk1x_en\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN[2]\);
    
    \imanches_in_dly[0]\ : SLE
      port map(D => \un1_manches_in[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \manches_in_dly[0]\);
    
    \RX_CENTER_SAMPLE_PROC.un16_irx_center_sample\ : CFG3
      generic map(INIT => x"40")

      port map(A => \clkdiv[2]_net_1\, B => \clkdiv[1]_net_1\, C
         => \clkdiv[0]_net_1\, Y => un16_irx_center_sample);
    
    \decoder_Transition_d[2]\ : SLE
      port map(D => \decoder_Transition_d[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clk1x_enable, ALn => un2_rst_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \decoder_Transition_d[2]_net_1\);
    
    \NRZ_DATA_PROC.un18_rst\ : CFG2
      generic map(INIT => x"1")

      port map(A => \idle_line\, B => RESET, Y => un18_rst_i);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \s2p_data[4]\ : SLE
      port map(D => \RX_FIFO_DIN[3]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => \sampler_clk1x_en\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN[4]\);
    
    clock_adjust_RNIMA1A : CFG1
      generic map(INIT => "01")

      port map(A => \clock_adjust\, Y => clock_adjust_i);
    
    \TRANISTION_DETECT_SHIFTREG_PROC.un2_rst\ : CFG2
      generic map(INIT => x"1")

      port map(A => rx_packet_end_all, B => RESET, Y => un2_rst_i);
    
    \SAMPLE_CLK1X_EN_PROC.isampler_clk1x_en_1\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \clkdiv[3]_net_1\, B => \clkdiv[0]_net_1\, C
         => \clkdiv[2]_net_1\, D => \clkdiv[1]_net_1\, Y => 
        isampler_clk1x_en_1);
    
    \irx_center_sample\ : SLE
      port map(D => un16_irx_center_sample, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clock_adjust_i, ALn => RESET_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => irx_center_sample_net_1);
    
    \clkdiv_3[2]\ : CFG3
      generic map(INIT => x"12")

      port map(A => \clkdiv[2]_net_1\, B => \un1_iidle_line\, C
         => CO1, Y => \clkdiv_3[2]_net_1\);
    
    \s2p_data[1]\ : SLE
      port map(D => \RX_FIFO_DIN[0]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => \sampler_clk1x_en\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN[1]\);
    
    \decoder_ShiftReg[0]\ : SLE
      port map(D => \clkdiv[3]_net_1\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => clk1x_enable, ALn => un2_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \decoder_ShiftReg[0]_net_1\);
    
    \clkdiv_3[1]\ : CFG4
      generic map(INIT => x"006A")

      port map(A => \clkdiv[1]_net_1\, B => \clkdiv[0]_net_1\, C
         => clk1x_enable, D => \un1_iidle_line\, Y => 
        \clkdiv_3[1]_net_1\);
    
    \manches_ShiftReg[0]\ : SLE
      port map(D => \manches_in_dly[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clk1x_enable, ALn => un2_rst_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \manches_ShiftReg[0]_net_1\);
    
    \iNRZ_data\ : SLE
      port map(D => iNRZ_data_1, CLK => CommsFPGA_CCC_0_GL0, EN
         => irx_center_sample_net_1, ALn => un18_rst_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => iNRZ_data_net_1);
    
    \clkdiv[2]\ : SLE
      port map(D => \clkdiv_3[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clock_adjust_i, ALn => RESET_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \clkdiv[2]_net_1\);
    
    \s2p_data[3]\ : SLE
      port map(D => \RX_FIFO_DIN[2]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => \sampler_clk1x_en\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN[3]\);
    
    \decoder_Transition_d[0]\ : SLE
      port map(D => \decoder_Transition\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clk1x_enable, ALn => un2_rst_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \decoder_Transition_d[0]_net_1\);
    
    decoder_Transition : SLE
      port map(D => decoder_Transition_1, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clk1x_enable, ALn => un2_rst_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \decoder_Transition\);
    
    \clkdiv_3[3]\ : CFG4
      generic map(INIT => x"FF6A")

      port map(A => \clkdiv[3]_net_1\, B => \clkdiv[2]_net_1\, C
         => CO1, D => \un1_iidle_line\, Y => \clkdiv_3[3]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \clkdiv[1]\ : SLE
      port map(D => \clkdiv_3[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clock_adjust_i, ALn => RESET_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \clkdiv[1]_net_1\);
    
    \s2p_data[5]\ : SLE
      port map(D => \RX_FIFO_DIN[4]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => \sampler_clk1x_en\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN[5]\);
    
    RX_IDLE_LINE_DETECTOR : IdleLineDetector_1
      port map(idle_line5 => idle_line5, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, RESET_i => RESET_i, idle_line => 
        \idle_line\);
    
    un10_clk1x_enable : CFG2
      generic map(INIT => x"6")

      port map(A => \clkdiv[3]_net_1\, B => 
        \decoder_ShiftReg[0]_net_1\, Y => decoder_Transition_1);
    
    clock_adjust : SLE
      port map(D => un16_clk1x_enable, CLK => CommsFPGA_CCC_0_GL0, 
        EN => clk1x_enable, ALn => un2_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \clock_adjust\);
    
    \un1_manches_in[0]\ : CFG3
      generic map(INIT => x"8D")

      port map(A => internal_loopback, B => MANCH_OUT_P_c, C => 
        MANCHESTER_IN_c, Y => \un1_manches_in[0]_net_1\);
    
    manches_Transition : SLE
      port map(D => manches_Transition_1, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clk1x_enable, ALn => un2_rst_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \manches_Transition\);
    
    \CLOCK_ADJUST_PROC.un16_clk1x_enable\ : CFG2
      generic map(INIT => x"8")

      port map(A => \decoder_Transition_d[2]_net_1\, B => 
        \manches_Transition\, Y => un16_clk1x_enable);
    
    \s2p_data[7]\ : SLE
      port map(D => \RX_FIFO_DIN[6]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => \sampler_clk1x_en\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => RX_FIFO_DIN(7));
    
    \clkdiv[0]\ : SLE
      port map(D => \clkdiv_3[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clock_adjust_i, ALn => RESET_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \clkdiv[0]_net_1\);
    
    \clkdiv[3]\ : SLE
      port map(D => \clkdiv_3[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clock_adjust_i, ALn => RESET_i, 
        ADn => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \clkdiv[3]_net_1\);
    
    un1_iidle_line : CFG2
      generic map(INIT => x"E")

      port map(A => \idle_line\, B => rx_packet_end_all, Y => 
        \un1_iidle_line\);
    
    \clkdiv_3[0]\ : CFG3
      generic map(INIT => x"06")

      port map(A => \clkdiv[0]_net_1\, B => clk1x_enable, C => 
        \un1_iidle_line\, Y => \clkdiv_3[0]_net_1\);
    
    \imanches_in_dly[1]\ : SLE
      port map(D => \manches_in_dly[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \manches_in_dly[1]\);
    
    \un1_clkdiv_1.CO1\ : CFG3
      generic map(INIT => x"80")

      port map(A => \clkdiv[1]_net_1\, B => \clkdiv[0]_net_1\, C
         => clk1x_enable, Y => CO1);
    
    \decoder_Transition_d[1]\ : SLE
      port map(D => \decoder_Transition_d[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clk1x_enable, ALn => un2_rst_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \decoder_Transition_d[1]_net_1\);
    
    \s2p_data[0]\ : SLE
      port map(D => iNRZ_data_net_1, CLK => CommsFPGA_CCC_0_GL0, 
        EN => \sampler_clk1x_en\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN[0]\);
    
    \NRZ_DATA_PROC.iNRZ_data_1\ : CFG2
      generic map(INIT => x"6")

      port map(A => \clkdiv[3]_net_1\, B => \manches_in_dly[1]\, 
        Y => iNRZ_data_1);
    
    \s2p_data[6]\ : SLE
      port map(D => \RX_FIFO_DIN[5]\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => \sampler_clk1x_en\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN[6]\);
    
    un4_clk1x_enable : CFG2
      generic map(INIT => x"6")

      port map(A => \manches_in_dly[1]\, B => 
        \manches_ShiftReg[0]_net_1\, Y => manches_Transition_1);
    
    isampler_clk1x_en : SLE
      port map(D => isampler_clk1x_en_1, CLK => 
        CommsFPGA_CCC_0_GL0, EN => clock_adjust_i, ALn => RESET_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \sampler_clk1x_en\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CRC16_Generator_1 is

    port( RX_FIFO_DIN         : in    std_logic_vector(7 downto 0);
          rx_crc_data_calc    : out   std_logic_vector(15 downto 0);
          rx_crc_gen          : in    std_logic;
          sampler_clk1x_en    : in    std_logic;
          iRX_FIFO_wr_en      : in    std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          rx_crc_reset_i      : in    std_logic
        );

end CRC16_Generator_1;

architecture DEF_ARCH of CRC16_Generator_1 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \rx_crc_data_calc[13]\, GND_net_1, 
        \rx_crc_data_calc[5]\, \lfsr_q_0_sqmuxa\, VCC_net_1, 
        \rx_crc_data_calc[14]\, \rx_crc_data_calc[6]\, 
        \rx_crc_data_calc[15]\, \lfsr_c[15]\, 
        \rx_crc_data_calc[0]\, \lfsr_c[0]\, \rx_crc_data_calc[1]\, 
        \lfsr_c[1]\, \rx_crc_data_calc[2]\, \lfsr_c[2]\, 
        \rx_crc_data_calc[3]\, \lfsr_c[3]\, \rx_crc_data_calc[4]\, 
        \lfsr_c[4]\, \lfsr_c[5]\, \lfsr_c[6]\, 
        \rx_crc_data_calc[7]\, \lfsr_c[7]\, \rx_crc_data_calc[8]\, 
        \lfsr_c[8]\, \rx_crc_data_calc[9]\, \lfsr_c[9]\, 
        \rx_crc_data_calc[10]\, \rx_crc_data_calc[11]\, 
        \rx_crc_data_calc[12]\, N_33 : std_logic;

begin 

    rx_crc_data_calc(15) <= \rx_crc_data_calc[15]\;
    rx_crc_data_calc(14) <= \rx_crc_data_calc[14]\;
    rx_crc_data_calc(13) <= \rx_crc_data_calc[13]\;
    rx_crc_data_calc(12) <= \rx_crc_data_calc[12]\;
    rx_crc_data_calc(11) <= \rx_crc_data_calc[11]\;
    rx_crc_data_calc(10) <= \rx_crc_data_calc[10]\;
    rx_crc_data_calc(9) <= \rx_crc_data_calc[9]\;
    rx_crc_data_calc(8) <= \rx_crc_data_calc[8]\;
    rx_crc_data_calc(7) <= \rx_crc_data_calc[7]\;
    rx_crc_data_calc(6) <= \rx_crc_data_calc[6]\;
    rx_crc_data_calc(5) <= \rx_crc_data_calc[5]\;
    rx_crc_data_calc(4) <= \rx_crc_data_calc[4]\;
    rx_crc_data_calc(3) <= \rx_crc_data_calc[3]\;
    rx_crc_data_calc(2) <= \rx_crc_data_calc[2]\;
    rx_crc_data_calc(1) <= \rx_crc_data_calc[1]\;
    rx_crc_data_calc(0) <= \rx_crc_data_calc[0]\;

    \lfsr_q[9]\ : SLE
      port map(D => \lfsr_c[9]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \lfsr_q_0_sqmuxa\, ALn => rx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_data_calc[9]\);
    
    \lfsr_q[6]\ : SLE
      port map(D => \lfsr_c[6]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \lfsr_q_0_sqmuxa\, ALn => rx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_data_calc[6]\);
    
    \lfsr_q[3]\ : SLE
      port map(D => \lfsr_c[3]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \lfsr_q_0_sqmuxa\, ALn => rx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_data_calc[3]\);
    
    \lfsr_q[10]\ : SLE
      port map(D => \rx_crc_data_calc[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \lfsr_q_0_sqmuxa\, ALn => 
        rx_crc_reset_i, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_calc[10]\);
    
    \lfsr_q[2]\ : SLE
      port map(D => \lfsr_c[2]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \lfsr_q_0_sqmuxa\, ALn => rx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_data_calc[2]\);
    
    \lfsr_c_0_a2_1[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => RX_FIFO_DIN(7), B => \rx_crc_data_calc[15]\, 
        Y => N_33);
    
    \lfsr_c_0_a2[5]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \rx_crc_data_calc[12]\, B => 
        \rx_crc_data_calc[11]\, C => RX_FIFO_DIN(4), D => 
        RX_FIFO_DIN(3), Y => \lfsr_c[5]\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \lfsr_q[1]\ : SLE
      port map(D => \lfsr_c[1]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \lfsr_q_0_sqmuxa\, ALn => rx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_data_calc[1]\);
    
    \lfsr_c_0_a2[4]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \rx_crc_data_calc[11]\, B => 
        \rx_crc_data_calc[10]\, C => RX_FIFO_DIN(3), D => 
        RX_FIFO_DIN(2), Y => \lfsr_c[4]\);
    
    \lfsr_q[7]\ : SLE
      port map(D => \lfsr_c[7]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \lfsr_q_0_sqmuxa\, ALn => rx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_data_calc[7]\);
    
    \lfsr_c_0_a2[3]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \rx_crc_data_calc[10]\, B => 
        \rx_crc_data_calc[9]\, C => RX_FIFO_DIN(2), D => 
        RX_FIFO_DIN(1), Y => \lfsr_c[3]\);
    
    \lfsr_q[4]\ : SLE
      port map(D => \lfsr_c[4]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \lfsr_q_0_sqmuxa\, ALn => rx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_data_calc[4]\);
    
    \lfsr_q[11]\ : SLE
      port map(D => \rx_crc_data_calc[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \lfsr_q_0_sqmuxa\, ALn => 
        rx_crc_reset_i, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_calc[11]\);
    
    \lfsr_q[5]\ : SLE
      port map(D => \lfsr_c[5]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \lfsr_q_0_sqmuxa\, ALn => rx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_data_calc[5]\);
    
    \lfsr_c_0_a2[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => N_33, B => \rx_crc_data_calc[1]\, Y => 
        \lfsr_c[9]\);
    
    \lfsr_c_0_a2[1]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => N_33, B => \lfsr_c[7]\, C => \lfsr_c[5]\, D
         => \lfsr_c[3]\, Y => \lfsr_c[1]\);
    
    \lfsr_q[0]\ : SLE
      port map(D => \lfsr_c[0]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \lfsr_q_0_sqmuxa\, ALn => rx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_data_calc[0]\);
    
    \lfsr_c_0_a2[7]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \rx_crc_data_calc[13]\, B => 
        \rx_crc_data_calc[14]\, C => RX_FIFO_DIN(6), D => 
        RX_FIFO_DIN(5), Y => \lfsr_c[7]\);
    
    \lfsr_c_0_a2[15]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \lfsr_c[0]\, B => \rx_crc_data_calc[7]\, Y
         => \lfsr_c[15]\);
    
    \lfsr_q[12]\ : SLE
      port map(D => \rx_crc_data_calc[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \lfsr_q_0_sqmuxa\, ALn => 
        rx_crc_reset_i, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_calc[12]\);
    
    \lfsr_c_0_a2[8]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \rx_crc_data_calc[14]\, B => 
        \rx_crc_data_calc[0]\, C => N_33, D => RX_FIFO_DIN(6), Y
         => \lfsr_c[8]\);
    
    \lfsr_c_0_a2[2]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \rx_crc_data_calc[9]\, B => 
        \rx_crc_data_calc[8]\, C => RX_FIFO_DIN(1), D => 
        RX_FIFO_DIN(0), Y => \lfsr_c[2]\);
    
    lfsr_q_0_sqmuxa : CFG3
      generic map(INIT => x"80")

      port map(A => iRX_FIFO_wr_en, B => sampler_clk1x_en, C => 
        rx_crc_gen, Y => \lfsr_q_0_sqmuxa\);
    
    \lfsr_q[14]\ : SLE
      port map(D => \rx_crc_data_calc[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \lfsr_q_0_sqmuxa\, ALn => 
        rx_crc_reset_i, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_calc[14]\);
    
    \lfsr_c_0_a2[6]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => \rx_crc_data_calc[13]\, B => 
        \rx_crc_data_calc[12]\, C => RX_FIFO_DIN(5), D => 
        RX_FIFO_DIN(4), Y => \lfsr_c[6]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \lfsr_q[8]\ : SLE
      port map(D => \lfsr_c[8]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \lfsr_q_0_sqmuxa\, ALn => rx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_data_calc[8]\);
    
    \lfsr_q[13]\ : SLE
      port map(D => \rx_crc_data_calc[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \lfsr_q_0_sqmuxa\, ALn => 
        rx_crc_reset_i, ADn => GND_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_calc[13]\);
    
    \lfsr_c_0_a2[0]\ : CFG3
      generic map(INIT => x"96")

      port map(A => RX_FIFO_DIN(0), B => \lfsr_c[1]\, C => 
        \rx_crc_data_calc[8]\, Y => \lfsr_c[0]\);
    
    \lfsr_q[15]\ : SLE
      port map(D => \lfsr_c[15]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \lfsr_q_0_sqmuxa\, ALn => rx_crc_reset_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_data_calc[15]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity ReadFIFO_Write_SM is

    port( consumer_type4_reg                 : in    std_logic_vector(9 downto 0);
          consumer_type3_reg                 : in    std_logic_vector(9 downto 0);
          consumer_type1_reg                 : in    std_logic_vector(9 downto 0);
          consumer_type2_reg                 : in    std_logic_vector(9 downto 0);
          CoreAPB3_0_APBmslave0_PRDATA_m     : out   std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PRDATA       : in    std_logic_vector(7 downto 0);
          un15                               : out   std_logic_vector(10 downto 0);
          RX_FIFO_DIN                        : in    std_logic_vector(7 downto 0);
          RX_FIFO_DIN_pipe                   : out   std_logic_vector(8 downto 0);
          DRVR_EN_c                          : in    std_logic;
          clk1x_enable                       : in    std_logic;
          CoreAPB3_0_APBmslave0_PREADY_i_m_i : out   std_logic;
          CoreAPB3_0_APBmslave0_PREADY       : in    std_logic;
          RESET                              : in    std_logic;
          RX_FIFO_TxColDetDis_wr_en          : out   std_logic;
          tx_col_detect_en                   : in    std_logic;
          idle_line                          : in    std_logic;
          CoreAPB3_0_APBmslave0_PSELx        : in    std_logic;
          sampler_clk1x_en                   : in    std_logic;
          packet_avail                       : in    std_logic;
          rx_packet_complt                   : out   std_logic;
          RX_EarlyTerm                       : out   std_logic;
          RESET_i                            : in    std_logic;
          CommsFPGA_CCC_0_GL0                : in    std_logic;
          rx_CRC_error_i                     : out   std_logic;
          rx_CRC_error                       : out   std_logic
        );

end ReadFIFO_Write_SM;

architecture DEF_ARCH of ReadFIFO_Write_SM is 

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CRC16_Generator_1
    port( RX_FIFO_DIN         : in    std_logic_vector(7 downto 0) := (others => 'U');
          rx_crc_data_calc    : out   std_logic_vector(15 downto 0);
          rx_crc_gen          : in    std_logic := 'U';
          sampler_clk1x_en    : in    std_logic := 'U';
          iRX_FIFO_wr_en      : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          rx_crc_reset_i      : in    std_logic := 'U'
        );
  end component;

    signal rx_crc_reset_i, \rx_crc_reset\, un9_rst, un9_rst_i, 
        rx_CRC_error_net_1, \bit_cntr[0]_net_1\, VCC_net_1, 
        un16_rst_i, N_44_i, GND_net_1, \bit_cntr[1]_net_1\, N_116, 
        \bit_cntr[2]_net_1\, N_117, \SM_advancebit_cntr[0]_net_1\, 
        N_45_i, \SM_advancebit_cntr[1]_net_1\, N_121, 
        \SM_advancebit_cntr[2]_net_1\, N_122, 
        \un65_sm_advance_i[4]\, \un65_sm_advance_i_i[4]\, 
        un1_ReadFIFO_WR_STATE_14, \un65_sm_advance_i[3]\, 
        \un65_sm_advance_i_i[3]\, \un65_sm_advance_i[2]\, 
        \un65_sm_advance_i_i[2]\, \un65_sm_advance_i[1]\, 
        \un65_sm_advance_i_i[1]\, \un56_sm_advance_i[11]\, 
        un56_sm_advance_i_cry_0_0_Y, \un56_sm_advance_i[10]\, 
        \un56_sm_advance_i_i[10]\, \un56_sm_advance_i[9]\, 
        \un56_sm_advance_i_i[9]\, \un56_sm_advance_i[8]\, 
        \un56_sm_advance_i_i[8]\, \un56_sm_advance_i[7]\, 
        \un56_sm_advance_i_i[7]\, \un56_sm_advance_i[6]\, 
        \un56_sm_advance_i_i[6]\, \un56_sm_advance_i[5]\, 
        \un56_sm_advance_i_i[5]\, \un56_sm_advance_i[4]\, 
        \un56_sm_advance_i_i[4]\, \un56_sm_advance_i[3]\, 
        \un56_sm_advance_i_i[3]\, \un56_sm_advance_i[2]\, 
        \un56_sm_advance_i_i[2]\, \un56_sm_advance_i[1]\, 
        \un56_sm_advance_i_i[1]\, \rx_packet_length[1]_net_1\, 
        \rx_packet_length_13[1]_net_1\, 
        \rx_packet_length[2]_net_1\, 
        \rx_packet_length_13[2]_net_1\, 
        \rx_packet_length[3]_net_1\, 
        \rx_packet_length_13[3]_net_1\, 
        \rx_packet_length[4]_net_1\, 
        \rx_packet_length_13[4]_net_1\, 
        \rx_packet_length[5]_net_1\, 
        \rx_packet_length_13[5]_net_1\, 
        \rx_packet_length[6]_net_1\, 
        \rx_packet_length_13[6]_net_1\, 
        \rx_packet_length[7]_net_1\, 
        \rx_packet_length_13[7]_net_1\, 
        \rx_packet_length[8]_net_1\, 
        \rx_packet_length_13[8]_net_1\, 
        \rx_packet_length[9]_net_1\, 
        \rx_packet_length_13[9]_net_1\, 
        \rx_packet_length[10]_net_1\, 
        \rx_packet_length_13[10]_net_1\, \un65_sm_advance_i[9]\, 
        \un65_sm_advance_i_i[9]\, \un65_sm_advance_i[8]\, 
        \un65_sm_advance_i_i[8]\, \un65_sm_advance_i[7]\, 
        \un65_sm_advance_i_i[7]\, \un65_sm_advance_i[6]\, 
        \un65_sm_advance_i_i[6]\, \un65_sm_advance_i[5]\, 
        \un65_sm_advance_i_i[5]\, \rx_crc_data_store[12]_net_1\, 
        \RX_FIFO_DIN_pipe[4]\, rx_crc_data_store_151, 
        \rx_crc_data_store[13]_net_1\, \RX_FIFO_DIN_pipe[5]\, 
        \rx_crc_data_store[14]_net_1\, \RX_FIFO_DIN_pipe[6]\, 
        \rx_crc_data_store[15]_net_1\, \RX_FIFO_DIN_pipe[7]\, 
        \consumer_type[0]_net_1\, \consumer_type_12[0]\, 
        un1_ReadFIFO_WR_STATE_12, \consumer_type[1]_net_1\, 
        \consumer_type_12[1]\, \consumer_type[2]_net_1\, 
        \consumer_type_12[2]\, \consumer_type[3]_net_1\, 
        \consumer_type_12[3]\, \consumer_type[4]_net_1\, 
        \consumer_type_12[4]\, \consumer_type[5]_net_1\, 
        \consumer_type_12[5]\, \consumer_type[6]_net_1\, 
        \consumer_type_12[6]\, \consumer_type[7]_net_1\, 
        \consumer_type_12[7]\, \consumer_type[8]_net_1\, 
        \consumer_type_12[8]\, \consumer_type[9]_net_1\, 
        \consumer_type_12[9]\, \rx_packet_length[0]_net_1\, 
        \rx_packet_length_13[0]_net_1\, 
        \rx_crc_data_store[0]_net_1\, 
        \un1_rx_fifo_din_d3[0]_net_1\, un1_sampler_clk1x_en_inv_i, 
        \rx_crc_data_store[1]_net_1\, 
        \un1_rx_fifo_din_d3[1]_net_1\, 
        \rx_crc_data_store[2]_net_1\, 
        \un1_rx_fifo_din_d3[2]_net_1\, 
        \rx_crc_data_store[3]_net_1\, 
        \un1_rx_fifo_din_d3[3]_net_1\, 
        \rx_crc_data_store[4]_net_1\, 
        \un1_rx_fifo_din_d3[4]_net_1\, 
        \rx_crc_data_store[5]_net_1\, 
        \un1_rx_fifo_din_d3[5]_net_1\, 
        \rx_crc_data_store[6]_net_1\, 
        \un1_rx_fifo_din_d3[6]_net_1\, 
        \rx_crc_data_store[7]_net_1\, 
        \un1_rx_fifo_din_d3[7]_net_1\, 
        \rx_crc_data_store[8]_net_1\, \RX_FIFO_DIN_pipe[0]\, 
        \rx_crc_data_store[9]_net_1\, \RX_FIFO_DIN_pipe[1]\, 
        \rx_crc_data_store[10]_net_1\, \RX_FIFO_DIN_pipe[2]\, 
        \rx_crc_data_store[11]_net_1\, \RX_FIFO_DIN_pipe[3]\, N_6, 
        \un1_sampler_clk1x_en_inv_0\, N_3, \iRX_FIFO_wr_en\, 
        un5_packet_avail, N_221, rx_packet_end, N_689_i, 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0\, \RX_FIFO_DIN_pipe[8]\, 
        \un15[3]\, \rx_crc_HighByte_en\, N_225_i, \rx_crc_gen\, 
        \un1_ReadFIFO_WR_STATE_15\, \SM_advance_i\, 
        un2_packet_avail, \rx_end_rst\, N_279_i, \RX_EarlyTerm\, 
        \un15[4]\, N_2, N_24, N_23, N_21, N_20, N_18, N_17, N_15, 
        N_14, N_12, N_11, N_9, N_8, N_5, \un65_sm_advance_i[10]\, 
        \un65_sm_advance_i_i[10]\, \rx_packet_complt_1_sqmuxa\, 
        N_676, \RX_InProcess\, N_314, 
        \ReadFIFO_WR_STATE_ns[5]_net_1\, 
        \ReadFIFO_WR_STATE_ns[6]_net_1\, \un15[2]\, \un15[1]\, 
        \ReadFIFO_WR_STATE_ns[8]_net_1\, \un15[0]\, 
        \ReadFIFO_WR_STATE_ns[9]_net_1\, \RX_InProcess_d1\, 
        \un15[10]\, N_253_i, \un15[9]\, 
        \ReadFIFO_WR_STATE_ns[1]_net_1\, \un15[8]\, 
        \ReadFIFO_WR_STATE_208\, \un15[7]\, 
        \ReadFIFO_WR_STATE_ns[3]\, \un15[5]\, 
        \ReadFIFO_WR_STATE_ns[4]_net_1\, \rx_byte_cntr[0]_net_1\, 
        \rx_byte_cntr_lm[0]\, rx_byte_cntre, 
        \rx_byte_cntr[1]_net_1\, \rx_byte_cntr_lm[1]\, 
        \rx_byte_cntr[2]_net_1\, \rx_byte_cntr_lm[2]\, 
        \rx_byte_cntr[3]_net_1\, \rx_byte_cntr_lm[3]\, 
        \rx_byte_cntr[4]_net_1\, \rx_byte_cntr_lm[4]\, 
        \rx_byte_cntr[5]_net_1\, \rx_byte_cntr_lm[5]\, 
        \rx_byte_cntr[6]_net_1\, \rx_byte_cntr_lm[6]\, 
        \rx_byte_cntr[7]_net_1\, \rx_byte_cntr_lm[7]\, 
        \rx_byte_cntr[8]_net_1\, \rx_byte_cntr_lm[8]\, 
        \rx_byte_cntr[9]_net_1\, \rx_byte_cntr_lm[9]\, 
        \rx_byte_cntr[10]_net_1\, \rx_byte_cntr_lm[10]\, 
        \rx_byte_cntr[11]_net_1\, \rx_byte_cntr_lm[11]\, 
        un56_sm_advance_i_cry_0, N_658_mux, 
        un56_sm_advance_i_cry_1, N_657_mux, 
        un56_sm_advance_i_cry_2, N_656_mux, 
        un56_sm_advance_i_cry_3, N_655_mux, 
        un56_sm_advance_i_cry_4, N_654_mux, 
        un56_sm_advance_i_cry_5, N_653_mux, 
        un56_sm_advance_i_cry_6, N_652_mux, 
        un56_sm_advance_i_cry_7, N_651_mux, 
        un56_sm_advance_i_cry_8, N_650_mux, 
        un65_sm_advance_i_cry_0, un65_sm_advance_i_cry_1, 
        un65_sm_advance_i_cry_2, un65_sm_advance_i_cry_3, 
        un65_sm_advance_i_cry_4, un65_sm_advance_i_cry_5, 
        un65_sm_advance_i_cry_6, un65_sm_advance_i_cry_7, 
        un65_sm_advance_i_cry_8, un67_sm_advance_i_cry_0, 
        un67_sm_advance_i_cry_1, un67_sm_advance_i_cry_2, 
        un67_sm_advance_i_cry_3, un67_sm_advance_i_cry_4, 
        un67_sm_advance_i_cry_5, un67_sm_advance_i_cry_6, 
        un67_sm_advance_i_cry_7, un67_sm_advance_i_cry_8, 
        un67_sm_advance_i_cry_9, un67_sm_advance_i_cry_10, 
        un67_sm_advance_i, \un58_sm_advance_i_0_data_tmp[0]\, 
        \un58_sm_advance_i_0_data_tmp[1]\, 
        \un58_sm_advance_i_0_data_tmp[2]\, 
        \un58_sm_advance_i_0_data_tmp[3]\, 
        \un58_sm_advance_i_0_data_tmp[4]\, 
        \un58_sm_advance_i_0_data_tmp[5]\, 
        \un1_sampler_clk1x_en_0_data_tmp[0]\, 
        \rx_crc_data_calc[0]\, \rx_crc_data_calc[1]\, 
        \un1_sampler_clk1x_en_0_data_tmp[1]\, 
        \rx_crc_data_calc[2]\, \rx_crc_data_calc[3]\, 
        \un1_sampler_clk1x_en_0_data_tmp[2]\, 
        \rx_crc_data_calc[4]\, \rx_crc_data_calc[5]\, 
        \un1_sampler_clk1x_en_0_data_tmp[3]\, 
        \rx_crc_data_calc[6]\, \rx_crc_data_calc[7]\, 
        \un1_sampler_clk1x_en_0_data_tmp[4]\, 
        \rx_crc_data_calc[8]\, \rx_crc_data_calc[9]\, 
        \un1_sampler_clk1x_en_0_data_tmp[5]\, 
        \rx_crc_data_calc[10]\, \rx_crc_data_calc[11]\, 
        \un1_sampler_clk1x_en_0_data_tmp[6]\, 
        \rx_crc_data_calc[12]\, \rx_crc_data_calc[13]\, 
        \un1_sampler_clk1x_en_0_data_tmp[7]\, 
        \rx_crc_data_calc[14]\, \rx_crc_data_calc[15]\, 
        rx_byte_cntr_s_916_FCO, \rx_byte_cntr_cry[1]_net_1\, 
        \rx_byte_cntr_s[1]\, \rx_byte_cntr_cry[2]_net_1\, 
        \rx_byte_cntr_s[2]\, \rx_byte_cntr_cry[3]_net_1\, 
        \rx_byte_cntr_s[3]\, \rx_byte_cntr_cry[4]_net_1\, 
        \rx_byte_cntr_s[4]\, \rx_byte_cntr_cry[5]_net_1\, 
        \rx_byte_cntr_s[5]\, \rx_byte_cntr_cry[6]_net_1\, 
        \rx_byte_cntr_s[6]\, \rx_byte_cntr_cry[7]_net_1\, 
        \rx_byte_cntr_s[7]\, \rx_byte_cntr_cry[8]_net_1\, 
        \rx_byte_cntr_s[8]\, \rx_byte_cntr_cry[9]_net_1\, 
        \rx_byte_cntr_s[9]\, \rx_byte_cntr_s[11]_net_1\, 
        \rx_byte_cntr_cry[10]_net_1\, \rx_byte_cntr_s[10]\, 
        un1_ReadFIFO_WR_STATE_6_i, N_649_mux, 
        un56_sm_advance_i_s_9_921_FCO, 
        un65_sm_advance_i_s_9_922_FCO, 
        \un65_sm_advance_i_cry_9_ma\, 
        \un56_sm_advance_i_cry_9_ma\, consumer_type_0_sqmuxa, 
        N_294, un1_iRX_EarlyTerm_0_sqmuxa, N_299, N_4706_i, 
        N_4729_i, un35_sm_advance_i_5, un38_sm_advance_i_5, 
        un29_sm_advance_i_5, un32_sm_advance_i_1, 
        consumer_type_12_sn_N_2, N_320, N_315, N_276, 
        un32_sm_advance_i_NE_4, un32_sm_advance_i_NE_3, 
        un32_sm_advance_i_NE_2, un32_sm_advance_i_NE_1, 
        un29_sm_advance_i_NE_4, un29_sm_advance_i_NE_3, 
        un29_sm_advance_i_NE_1, un29_sm_advance_i_NE_0, 
        un35_sm_advance_i_NE_4, un35_sm_advance_i_NE_3, 
        un35_sm_advance_i_NE_1, un35_sm_advance_i_NE_0, 
        un38_sm_advance_i_NE_4, un38_sm_advance_i_NE_3, 
        un38_sm_advance_i_NE_1, un38_sm_advance_i_NE_0, 
        \rx_crc_gen_3_sqmuxa\, 
        \ReadFIFO_WR_STATE_ns_a3_0_0[3]_net_1\, N_661, N_321, 
        \ReadFIFO_WR_STATE_ns_0[5]_net_1\, un32_sm_advance_i_NE_5, 
        un29_sm_advance_i_NE_6, un35_sm_advance_i_NE_6, 
        un38_sm_advance_i_NE_6, N_308, un29_sm_advance_i_NE_7, 
        un35_sm_advance_i_NE_7, un38_sm_advance_i_NE_7, 
        un33_sm_advance_i, un40_sm_advance_i_1, 
        un40_sm_advance_i_2, 
        \ReadFIFO_WR_STATE_ns_a3_0_1_0[3]_net_1\ : std_logic;

    for all : CRC16_Generator_1
	Use entity work.CRC16_Generator_1(DEF_ARCH);
begin 

    un15(10) <= \un15[10]\;
    un15(9) <= \un15[9]\;
    un15(8) <= \un15[8]\;
    un15(7) <= \un15[7]\;
    un15(5) <= \un15[5]\;
    un15(4) <= \un15[4]\;
    un15(3) <= \un15[3]\;
    un15(2) <= \un15[2]\;
    un15(1) <= \un15[1]\;
    un15(0) <= \un15[0]\;
    RX_FIFO_DIN_pipe(8) <= \RX_FIFO_DIN_pipe[8]\;
    RX_FIFO_DIN_pipe(7) <= \RX_FIFO_DIN_pipe[7]\;
    RX_FIFO_DIN_pipe(6) <= \RX_FIFO_DIN_pipe[6]\;
    RX_FIFO_DIN_pipe(5) <= \RX_FIFO_DIN_pipe[5]\;
    RX_FIFO_DIN_pipe(4) <= \RX_FIFO_DIN_pipe[4]\;
    RX_FIFO_DIN_pipe(3) <= \RX_FIFO_DIN_pipe[3]\;
    RX_FIFO_DIN_pipe(2) <= \RX_FIFO_DIN_pipe[2]\;
    RX_FIFO_DIN_pipe(1) <= \RX_FIFO_DIN_pipe[1]\;
    RX_FIFO_DIN_pipe(0) <= \RX_FIFO_DIN_pipe[0]\;
    RX_EarlyTerm <= \RX_EarlyTerm\;
    rx_CRC_error <= rx_CRC_error_net_1;

    un65_sm_advance_i_s_9_922 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => un65_sm_advance_i_cry_8, C
         => GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => 
        OPEN, Y => OPEN, FCO => un65_sm_advance_i_s_9_922_FCO);
    
    \ReadFIFO_WR_STATE_RNIL7N4[3]\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \un15[5]\, B => \un15[3]\, C => \un15[7]\, D
         => \un15[8]\, Y => N_314);
    
    \rx_packet_length[5]\ : SLE
      port map(D => \rx_packet_length_13[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rx_packet_length[5]_net_1\);
    
    \rx_packet_length_RNI4CTA1[2]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => RX_FIFO_DIN(2), B => N_299, C => 
        \rx_packet_length[2]_net_1\, Y => N_657_mux);
    
    \ReadFIFO_WR_SM.un35_sm_advance_i_NE_4\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type3_reg(9), B => 
        consumer_type3_reg(8), C => \consumer_type[9]_net_1\, D
         => \consumer_type[8]_net_1\, Y => un35_sm_advance_i_NE_4);
    
    \rx_packet_length_ret[4]\ : SLE
      port map(D => \un56_sm_advance_i_i[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \un56_sm_advance_i[7]\);
    
    un56_sm_advance_i_cry_5_0 : ARI1
      generic map(INIT => x"511FF")

      port map(A => N_653_mux, B => \un15[7]\, C => \un15[8]\, D
         => GND_net_1, FCI => un56_sm_advance_i_cry_4, S => 
        \un56_sm_advance_i_i[6]\, Y => OPEN, FCO => 
        un56_sm_advance_i_cry_5);
    
    rx_crc_LowByte_en : SLE
      port map(D => \un15[3]\, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN_pipe[8]\);
    
    \ReadFIFO_WR_STATE_ns[4]\ : CFG4
      generic map(INIT => x"FF8C")

      port map(A => \un58_sm_advance_i_0_data_tmp[5]\, B => 
        \un15[5]\, C => \un1_sampler_clk1x_en_inv_0\, D => N_299, 
        Y => \ReadFIFO_WR_STATE_ns[4]_net_1\);
    
    \ReadFIFO_WR_SM.un38_sm_advance_i_NE_7\ : CFG3
      generic map(INIT => x"FE")

      port map(A => un38_sm_advance_i_NE_4, B => 
        un38_sm_advance_i_NE_1, C => un38_sm_advance_i_NE_0, Y
         => un38_sm_advance_i_NE_7);
    
    \ReadFIFO_WR_SM.un58_sm_advance_i_0_I_27\ : ARI1
      generic map(INIT => x"68241")

      port map(A => \un56_sm_advance_i[4]\, B => 
        \rx_byte_cntr[8]_net_1\, C => \rx_byte_cntr[9]_net_1\, D
         => \un56_sm_advance_i[3]\, FCI => 
        \un58_sm_advance_i_0_data_tmp[3]\, S => OPEN, Y => OPEN, 
        FCO => \un58_sm_advance_i_0_data_tmp[4]\);
    
    un1_iRX_EarlyTerm_0_sqmuxa_0_a3 : CFG3
      generic map(INIT => x"2A")

      port map(A => \un15[10]\, B => \un1_sampler_clk1x_en_inv_0\, 
        C => packet_avail, Y => N_308);
    
    \rx_byte_cntr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rx_byte_cntr[10]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \rx_byte_cntr_cry[9]_net_1\, S => \rx_byte_cntr_s[10]\, Y
         => OPEN, FCO => \rx_byte_cntr_cry[10]_net_1\);
    
    \rx_packet_length_ret[0]\ : SLE
      port map(D => un56_sm_advance_i_cry_0_0_Y, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \un56_sm_advance_i[11]\);
    
    \rx_byte_cntr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rx_byte_cntr[9]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \rx_byte_cntr_cry[8]_net_1\, S => \rx_byte_cntr_s[9]\, Y
         => OPEN, FCO => \rx_byte_cntr_cry[9]_net_1\);
    
    \ReadFIFO_WR_SM.un32_sm_advance_i_NE_2\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type2_reg(5), B => 
        consumer_type2_reg(4), C => \consumer_type[5]_net_1\, D
         => \consumer_type[4]_net_1\, Y => un32_sm_advance_i_NE_2);
    
    un56_sm_advance_i_cry_3_0 : ARI1
      generic map(INIT => x"511FF")

      port map(A => N_655_mux, B => \un15[7]\, C => \un15[8]\, D
         => GND_net_1, FCI => un56_sm_advance_i_cry_2, S => 
        \un56_sm_advance_i_i[8]\, Y => OPEN, FCO => 
        un56_sm_advance_i_cry_3);
    
    un65_sm_advance_i_s_10_RNO : CFG2
      generic map(INIT => x"7")

      port map(A => N_649_mux, B => un1_ReadFIFO_WR_STATE_6_i, Y
         => N_4706_i);
    
    \SM_advancebit_cntr_RNO[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => N_221, B => \SM_advancebit_cntr[0]_net_1\, Y
         => N_45_i);
    
    \rx_packet_length[10]\ : SLE
      port map(D => \rx_packet_length_13[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rx_packet_length[10]_net_1\);
    
    \rx_byte_cntr[11]\ : SLE
      port map(D => \rx_byte_cntr_lm[11]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => rx_byte_cntre, ALn => RESET_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \rx_byte_cntr[11]_net_1\);
    
    \ReadFIFO_WR_SM.un58_sm_advance_i_0_I_33\ : ARI1
      generic map(INIT => x"68241")

      port map(A => \un56_sm_advance_i[8]\, B => 
        \rx_byte_cntr[4]_net_1\, C => \rx_byte_cntr[5]_net_1\, D
         => \un56_sm_advance_i[7]\, FCI => 
        \un58_sm_advance_i_0_data_tmp[1]\, S => OPEN, Y => OPEN, 
        FCO => \un58_sm_advance_i_0_data_tmp[2]\);
    
    \ReadFIFO_WR_STATE[4]\ : SLE
      port map(D => \ReadFIFO_WR_STATE_ns[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \un15[4]\);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_6\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[6]_net_1\, B => 
        \un65_sm_advance_i[6]\, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_5, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_6);
    
    rx_end_rst : SLE
      port map(D => N_279_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0\, ALn => RESET_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_end_rst\);
    
    \ReadFIFO_WR_STATE_ns_a3_0_1[3]\ : CFG3
      generic map(INIT => x"DC")

      port map(A => un40_sm_advance_i_2, B => 
        \ReadFIFO_WR_STATE_ns_a3_0_1_0[3]_net_1\, C => 
        \ReadFIFO_WR_STATE_ns_a3_0_0[3]_net_1\, Y => 
        \ReadFIFO_WR_STATE_ns[3]\);
    
    \rx_packet_length_ret[5]\ : SLE
      port map(D => \un56_sm_advance_i_i[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \un56_sm_advance_i[6]\);
    
    \rx_fifo_din_d3[2]\ : SLE
      port map(D => N_9, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_sampler_clk1x_en_inv_0\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN_pipe[2]\);
    
    \SM_advancebit_cntr[0]\ : SLE
      port map(D => N_45_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => un9_rst_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SM_advancebit_cntr[0]_net_1\);
    
    \rx_byte_cntr_lm_0[1]\ : CFG2
      generic map(INIT => x"4")

      port map(A => un1_iRX_EarlyTerm_0_sqmuxa, B => 
        \rx_byte_cntr_s[1]\, Y => \rx_byte_cntr_lm[1]\);
    
    iRX_FIFO_wr_en : SLE
      port map(D => un5_packet_avail, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_221, ALn => un16_rst_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \iRX_FIFO_wr_en\);
    
    \rx_packet_length[8]\ : SLE
      port map(D => \rx_packet_length_13[8]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rx_packet_length[8]_net_1\);
    
    \ReadFIFO_WR_STATE_ns[8]\ : CFG4
      generic map(INIT => x"E222")

      port map(A => \un15[1]\, B => sampler_clk1x_en, C => 
        \SM_advance_i\, D => \un15[2]\, Y => 
        \ReadFIFO_WR_STATE_ns[8]_net_1\);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_1\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[1]_net_1\, B => 
        \un56_sm_advance_i[11]\, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_0, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_1);
    
    \rx_packet_length_ret[2]\ : SLE
      port map(D => \un56_sm_advance_i_i[9]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \un56_sm_advance_i[9]\);
    
    consumer_type_0_sqmuxa_0_a3 : CFG3
      generic map(INIT => x"80")

      port map(A => \un15[10]\, B => \un1_sampler_clk1x_en_inv_0\, 
        C => packet_avail, Y => consumer_type_0_sqmuxa);
    
    \consumer_type[4]\ : SLE
      port map(D => \consumer_type_12[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_12, ALn
         => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type[4]_net_1\);
    
    \rx_byte_cntr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rx_byte_cntr[8]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \rx_byte_cntr_cry[7]_net_1\, S => \rx_byte_cntr_s[8]\, Y
         => OPEN, FCO => \rx_byte_cntr_cry[8]_net_1\);
    
    \CoreAPB3_0_APBmslave0_PRDATA_m[3]\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        CoreAPB3_0_APBmslave0_PRDATA(3), Y => 
        CoreAPB3_0_APBmslave0_PRDATA_m(3));
    
    \rx_packet_length_ret_1[6]\ : SLE
      port map(D => \un65_sm_advance_i_i[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \un65_sm_advance_i[3]\);
    
    \rx_fifo_din_d1[0]\ : SLE
      port map(D => RX_FIFO_DIN(0), CLK => CommsFPGA_CCC_0_GL0, 
        EN => \un1_sampler_clk1x_en_inv_0\, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => N_2);
    
    \rx_packet_length_13[10]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_649_mux, B => un1_ReadFIFO_WR_STATE_6_i, Y
         => \rx_packet_length_13[10]_net_1\);
    
    \rx_byte_cntr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rx_byte_cntr[3]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \rx_byte_cntr_cry[2]_net_1\, S => \rx_byte_cntr_s[3]\, Y
         => OPEN, FCO => \rx_byte_cntr_cry[3]_net_1\);
    
    \ReadFIFO_WR_SM.un38_sm_advance_i_NE_0\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type4_reg(1), B => 
        consumer_type4_reg(0), C => \consumer_type[1]_net_1\, D
         => \consumer_type[0]_net_1\, Y => un38_sm_advance_i_NE_0);
    
    \SM_ADVANCE_PROC.un2_packet_avail\ : CFG3
      generic map(INIT => x"80")

      port map(A => \SM_advancebit_cntr[2]_net_1\, B => 
        \SM_advancebit_cntr[1]_net_1\, C => 
        \SM_advancebit_cntr[0]_net_1\, Y => un2_packet_avail);
    
    \ReadFIFO_WR_STATE_ns_i_a2[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \un15[0]\, B => \un15[4]\, Y => N_320);
    
    \rx_crc_data_store[1]\ : SLE
      port map(D => \un1_rx_fifo_din_d3[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_sampler_clk1x_en_inv_i, 
        ALn => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[1]_net_1\);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_11\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[11]_net_1\, B => 
        \un65_sm_advance_i[1]\, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_10, S => OPEN, Y => OPEN, 
        FCO => un67_sm_advance_i);
    
    \ReadFIFO_WRITE_PROC.un16_rst\ : CFG2
      generic map(INIT => x"1")

      port map(A => un9_rst, B => rx_packet_end, Y => un16_rst_i);
    
    \rx_packet_length_RNIVC031[10]\ : CFG4
      generic map(INIT => x"CCAC")

      port map(A => RX_FIFO_DIN(2), B => 
        \rx_packet_length[10]_net_1\, C => 
        \un1_sampler_clk1x_en_inv_0\, D => \un15[7]\, Y => 
        N_649_mux);
    
    un56_sm_advance_i_s_10 : CFG3
      generic map(INIT => x"27")

      port map(A => N_4729_i, B => un56_sm_advance_i_cry_8, C => 
        \un56_sm_advance_i_cry_9_ma\, Y => 
        \un56_sm_advance_i_i[1]\);
    
    \rx_byte_cntr_lm_0[0]\ : CFG2
      generic map(INIT => x"1")

      port map(A => un1_iRX_EarlyTerm_0_sqmuxa, B => 
        \rx_byte_cntr[0]_net_1\, Y => \rx_byte_cntr_lm[0]\);
    
    \ReadFIFO_WR_SM.un58_sm_advance_i_0_I_9\ : ARI1
      generic map(INIT => x"68241")

      port map(A => \un56_sm_advance_i[2]\, B => 
        \rx_byte_cntr[10]_net_1\, C => \rx_byte_cntr[11]_net_1\, 
        D => \un56_sm_advance_i[1]\, FCI => 
        \un58_sm_advance_i_0_data_tmp[4]\, S => OPEN, Y => OPEN, 
        FCO => \un58_sm_advance_i_0_data_tmp[5]\);
    
    \un1_rx_fifo_din_d3[4]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \RX_FIFO_DIN_pipe[4]\, B => 
        \rx_crc_HighByte_en\, Y => \un1_rx_fifo_din_d3[4]_net_1\);
    
    \rx_byte_cntr_lm_0[6]\ : CFG2
      generic map(INIT => x"4")

      port map(A => un1_iRX_EarlyTerm_0_sqmuxa, B => 
        \rx_byte_cntr_s[6]\, Y => \rx_byte_cntr_lm[6]\);
    
    \CoreAPB3_0_APBmslave0_PRDATA_m[2]\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        CoreAPB3_0_APBmslave0_PRDATA(2), Y => 
        CoreAPB3_0_APBmslave0_PRDATA_m(2));
    
    \rx_fifo_din_d3[4]\ : SLE
      port map(D => N_15, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_sampler_clk1x_en_inv_0\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN_pipe[4]\);
    
    \consumer_type[7]\ : SLE
      port map(D => \consumer_type_12[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_12, ALn
         => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type[7]_net_1\);
    
    \ReadFIFO_WR_STATE_RNO[9]\ : CFG4
      generic map(INIT => x"00AE")

      port map(A => \un15[10]\, B => idle_line, C => N_320, D => 
        N_294, Y => N_253_i);
    
    un65_sm_advance_i_cry_3_0 : ARI1
      generic map(INIT => x"511FF")

      port map(A => N_655_mux, B => \un15[7]\, C => \un15[8]\, D
         => GND_net_1, FCI => un65_sm_advance_i_cry_2, S => 
        \un65_sm_advance_i_i[8]\, Y => OPEN, FCO => 
        un65_sm_advance_i_cry_3);
    
    \ReadFIFO_WR_SM.consumer_type_12[9]\ : CFG4
      generic map(INIT => x"E4A0")

      port map(A => \un15[9]\, B => consumer_type_0_sqmuxa, C => 
        \consumer_type[9]_net_1\, D => RX_FIFO_DIN(7), Y => 
        \consumer_type_12[9]\);
    
    un56_sm_advance_i_cry_0_0 : ARI1
      generic map(INIT => x"511FF")

      port map(A => N_658_mux, B => \un15[7]\, C => \un15[8]\, D
         => GND_net_1, FCI => GND_net_1, S => OPEN, Y => 
        un56_sm_advance_i_cry_0_0_Y, FCO => 
        un56_sm_advance_i_cry_0);
    
    \rx_fifo_din_d1[5]\ : SLE
      port map(D => RX_FIFO_DIN(5), CLK => CommsFPGA_CCC_0_GL0, 
        EN => \un1_sampler_clk1x_en_inv_0\, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => N_17);
    
    \ReadFIFO_WR_STATE_ns[5]\ : CFG4
      generic map(INIT => x"EAAA")

      port map(A => \ReadFIFO_WR_STATE_ns_0[5]_net_1\, B => 
        un40_sm_advance_i_1, C => 
        \ReadFIFO_WR_STATE_ns_a3_0_0[3]_net_1\, D => 
        un40_sm_advance_i_2, Y => \ReadFIFO_WR_STATE_ns[5]_net_1\);
    
    \ReadFIFO_WR_SM.un1_sampler_clk1x_en_0_I_45\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \rx_crc_data_store[9]_net_1\, B => 
        \rx_crc_data_calc[8]\, C => \rx_crc_data_calc[9]\, D => 
        \rx_crc_data_store[8]_net_1\, FCI => 
        \un1_sampler_clk1x_en_0_data_tmp[3]\, S => OPEN, Y => 
        OPEN, FCO => \un1_sampler_clk1x_en_0_data_tmp[4]\);
    
    \CoreAPB3_0_APBmslave0_PRDATA_m[7]\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        CoreAPB3_0_APBmslave0_PRDATA(7), Y => 
        CoreAPB3_0_APBmslave0_PRDATA_m(7));
    
    \rx_crc_data_store[12]\ : SLE
      port map(D => \RX_FIFO_DIN_pipe[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => rx_crc_data_store_151, ALn => 
        RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[12]_net_1\);
    
    un56_sm_advance_i_cry_6_0 : ARI1
      generic map(INIT => x"511FF")

      port map(A => N_652_mux, B => \un15[7]\, C => \un15[8]\, D
         => GND_net_1, FCI => un56_sm_advance_i_cry_5, S => 
        \un56_sm_advance_i_i[5]\, Y => OPEN, FCO => 
        un56_sm_advance_i_cry_6);
    
    rx_crc_HighByte_en : SLE
      port map(D => N_225_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_HighByte_en\);
    
    \rx_byte_cntr_lm_0[5]\ : CFG2
      generic map(INIT => x"4")

      port map(A => un1_iRX_EarlyTerm_0_sqmuxa, B => 
        \rx_byte_cntr_s[5]\, Y => \rx_byte_cntr_lm[5]\);
    
    \ReadFIFO_WR_SM.un29_sm_advance_i_NE_7\ : CFG3
      generic map(INIT => x"FE")

      port map(A => un29_sm_advance_i_NE_4, B => 
        un29_sm_advance_i_NE_1, C => un29_sm_advance_i_NE_0, Y
         => un29_sm_advance_i_NE_7);
    
    \rx_packet_length_RNIKI731[8]\ : CFG4
      generic map(INIT => x"CCAC")

      port map(A => RX_FIFO_DIN(0), B => 
        \rx_packet_length[8]_net_1\, C => 
        \un1_sampler_clk1x_en_inv_0\, D => \un15[7]\, Y => 
        N_651_mux);
    
    un65_sm_advance_i_cry_4_0 : ARI1
      generic map(INIT => x"511FF")

      port map(A => N_654_mux, B => \un15[7]\, C => \un15[8]\, D
         => GND_net_1, FCI => un65_sm_advance_i_cry_3, S => 
        \un65_sm_advance_i_i[7]\, Y => OPEN, FCO => 
        un65_sm_advance_i_cry_4);
    
    \rx_CRC_error\ : SLE
      port map(D => N_676, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => rx_CRC_error_net_1);
    
    \rx_crc_data_store[8]\ : SLE
      port map(D => \RX_FIFO_DIN_pipe[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => rx_crc_data_store_151, ALn => 
        RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[8]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    un56_sm_advance_i_s_10_RNO : CFG2
      generic map(INIT => x"7")

      port map(A => N_649_mux, B => un1_ReadFIFO_WR_STATE_6_i, Y
         => N_4729_i);
    
    \rx_fifo_din_d1[2]\ : SLE
      port map(D => RX_FIFO_DIN(2), CLK => CommsFPGA_CCC_0_GL0, 
        EN => \un1_sampler_clk1x_en_inv_0\, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => N_8);
    
    ReadFIFO_WR_STATE_208 : CFG3
      generic map(INIT => x"AC")

      port map(A => \un15[9]\, B => \un15[8]\, C => 
        \un1_sampler_clk1x_en_inv_0\, Y => 
        \ReadFIFO_WR_STATE_208\);
    
    \consumer_type[6]\ : SLE
      port map(D => \consumer_type_12[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_12, ALn
         => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type[6]_net_1\);
    
    \rx_crc_data_store[5]\ : SLE
      port map(D => \un1_rx_fifo_din_d3[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_sampler_clk1x_en_inv_i, 
        ALn => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[5]_net_1\);
    
    \ReadFIFO_WR_SM.un1_sampler_clk1x_en_0_I_9\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \rx_crc_data_store[3]_net_1\, B => 
        \rx_crc_data_calc[2]\, C => \rx_crc_data_calc[3]\, D => 
        \rx_crc_data_store[2]_net_1\, FCI => 
        \un1_sampler_clk1x_en_0_data_tmp[0]\, S => OPEN, Y => 
        OPEN, FCO => \un1_sampler_clk1x_en_0_data_tmp[1]\);
    
    \rx_packet_length_RNI8GTA1[4]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => RX_FIFO_DIN(4), B => N_299, C => 
        \rx_packet_length[4]_net_1\, Y => N_655_mux);
    
    \rx_packet_length[6]\ : SLE
      port map(D => \rx_packet_length_13[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rx_packet_length[6]_net_1\);
    
    \ReadFIFO_WR_STATE[2]\ : SLE
      port map(D => \un15[3]\, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_sampler_clk1x_en_inv_0\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \un15[2]\);
    
    un65_sm_advance_i_cry_9_ma : CFG2
      generic map(INIT => x"8")

      port map(A => N_649_mux, B => un1_ReadFIFO_WR_STATE_6_i, Y
         => \un65_sm_advance_i_cry_9_ma\);
    
    un56_sm_advance_i_s_9_921 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => un56_sm_advance_i_cry_8, C
         => GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => 
        OPEN, Y => OPEN, FCO => un56_sm_advance_i_s_9_921_FCO);
    
    \rx_byte_cntr[1]\ : SLE
      port map(D => \rx_byte_cntr_lm[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => rx_byte_cntre, ALn => RESET_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \rx_byte_cntr[1]_net_1\);
    
    \ReadFIFO_WR_SM.un58_sm_advance_i_0_I_1\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \un56_sm_advance_i[11]\, B => 
        \rx_byte_cntr[0]_net_1\, C => \rx_byte_cntr[1]_net_1\, D
         => \rx_packet_length[0]_net_1\, FCI => GND_net_1, S => 
        OPEN, Y => OPEN, FCO => \un58_sm_advance_i_0_data_tmp[0]\);
    
    \ReadFIFO_WR_STATE_RNIEGKD[8]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \un1_sampler_clk1x_en_inv_0\, B => \un15[9]\, 
        Y => N_661);
    
    \ReadFIFO_WR_SM.un38_sm_advance_i_NE_1\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type4_reg(3), B => 
        consumer_type4_reg(2), C => \consumer_type[3]_net_1\, D
         => \consumer_type[2]_net_1\, Y => un38_sm_advance_i_NE_1);
    
    \rx_byte_cntr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rx_byte_cntr[7]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \rx_byte_cntr_cry[6]_net_1\, S => \rx_byte_cntr_s[7]\, Y
         => OPEN, FCO => \rx_byte_cntr_cry[7]_net_1\);
    
    \rx_packet_complt\ : SLE
      port map(D => \rx_packet_complt_1_sqmuxa\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => rx_packet_complt);
    
    iRX_EarlyTerm : SLE
      port map(D => \un15[4]\, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_EarlyTerm\);
    
    \rx_packet_length_13[0]\ : CFG4
      generic map(INIT => x"CA00")

      port map(A => \rx_packet_length[0]_net_1\, B => 
        RX_FIFO_DIN(0), C => N_299, D => 
        un1_ReadFIFO_WR_STATE_6_i, Y => 
        \rx_packet_length_13[0]_net_1\);
    
    \ReadFIFO_WR_SM.consumer_type_12[4]\ : CFG4
      generic map(INIT => x"E4A0")

      port map(A => \un15[9]\, B => consumer_type_0_sqmuxa, C => 
        \consumer_type[4]_net_1\, D => RX_FIFO_DIN(2), Y => 
        \consumer_type_12[4]\);
    
    \ReadFIFO_WR_SM.un58_sm_advance_i_0_I_21\ : ARI1
      generic map(INIT => x"68241")

      port map(A => \un56_sm_advance_i[6]\, B => 
        \rx_byte_cntr[6]_net_1\, C => \rx_byte_cntr[7]_net_1\, D
         => \un56_sm_advance_i[5]\, FCI => 
        \un58_sm_advance_i_0_data_tmp[2]\, S => OPEN, Y => OPEN, 
        FCO => \un58_sm_advance_i_0_data_tmp[3]\);
    
    \rx_packet_length_ret[8]\ : SLE
      port map(D => \un56_sm_advance_i_i[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \un56_sm_advance_i[3]\);
    
    \ReadFIFO_WR_SM.un38_sm_advance_i_NE_4\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type4_reg(9), B => 
        consumer_type4_reg(8), C => \consumer_type[9]_net_1\, D
         => \consumer_type[8]_net_1\, Y => un38_sm_advance_i_NE_4);
    
    \ReadFIFO_WR_SM.un1_sampler_clk1x_en_0_I_21\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \rx_crc_data_store[15]_net_1\, B => 
        \rx_crc_data_calc[14]\, C => \rx_crc_data_calc[15]\, D
         => \rx_crc_data_store[14]_net_1\, FCI => 
        \un1_sampler_clk1x_en_0_data_tmp[6]\, S => OPEN, Y => 
        OPEN, FCO => \un1_sampler_clk1x_en_0_data_tmp[7]\);
    
    \bit_cntr[2]\ : SLE
      port map(D => N_117, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => un16_rst_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \bit_cntr[2]_net_1\);
    
    \rx_packet_length_ret_1[0]\ : SLE
      port map(D => \un65_sm_advance_i_i[9]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \un65_sm_advance_i[9]\);
    
    \rx_packet_length_13[3]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_656_mux, B => un1_ReadFIFO_WR_STATE_6_i, Y
         => \rx_packet_length_13[3]_net_1\);
    
    \ReadFIFO_WR_SM.un35_sm_advance_i_5\ : CFG2
      generic map(INIT => x"6")

      port map(A => \consumer_type[5]_net_1\, B => 
        consumer_type3_reg(5), Y => un35_sm_advance_i_5);
    
    \bit_cntr[0]\ : SLE
      port map(D => N_44_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => un16_rst_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \bit_cntr[0]_net_1\);
    
    \ReadFIFO_WR_SM.un32_sm_advance_i_NE\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => un32_sm_advance_i_NE_2, B => 
        un32_sm_advance_i_NE_5, C => un32_sm_advance_i_NE_4, D
         => un32_sm_advance_i_NE_3, Y => un33_sm_advance_i);
    
    \ReadFIFO_WR_SM.un29_sm_advance_i_NE_4\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type1_reg(9), B => 
        consumer_type1_reg(8), C => \consumer_type[9]_net_1\, D
         => \consumer_type[8]_net_1\, Y => un29_sm_advance_i_NE_4);
    
    \rx_byte_cntr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rx_byte_cntr[4]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \rx_byte_cntr_cry[3]_net_1\, S => \rx_byte_cntr_s[4]\, Y
         => OPEN, FCO => \rx_byte_cntr_cry[4]_net_1\);
    
    \rx_packet_length_ret[1]\ : SLE
      port map(D => \un56_sm_advance_i_i[10]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \un56_sm_advance_i[10]\);
    
    \rx_packet_length_13[5]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_654_mux, B => un1_ReadFIFO_WR_STATE_6_i, Y
         => \rx_packet_length_13[5]_net_1\);
    
    \rx_packet_length_13[6]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_653_mux, B => un1_ReadFIFO_WR_STATE_6_i, Y
         => \rx_packet_length_13[6]_net_1\);
    
    \ReadFIFO_WR_SM.un32_sm_advance_i_1\ : CFG2
      generic map(INIT => x"6")

      port map(A => \consumer_type[1]_net_1\, B => 
        consumer_type2_reg(1), Y => un32_sm_advance_i_1);
    
    \ReadFIFO_WR_STATE_ns[9]\ : CFG4
      generic map(INIT => x"4F44")

      port map(A => idle_line, B => \un15[0]\, C => 
        \un1_sampler_clk1x_en_0_data_tmp[7]\, D => N_315, Y => 
        \ReadFIFO_WR_STATE_ns[9]_net_1\);
    
    \rx_packet_length_ret_1[3]\ : SLE
      port map(D => \un65_sm_advance_i_i[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \un65_sm_advance_i[6]\);
    
    SM_advance_i_RNI0CAL : CFG3
      generic map(INIT => x"80")

      port map(A => \SM_advance_i\, B => sampler_clk1x_en, C => 
        \un15[7]\, Y => N_299);
    
    \rx_packet_length_ret[9]\ : SLE
      port map(D => \un56_sm_advance_i_i[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \un56_sm_advance_i[2]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \ReadFIFO_WR_STATE[7]\ : SLE
      port map(D => \ReadFIFO_WR_STATE_208\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \un15[8]\);
    
    \rx_fifo_din_d2[6]\ : SLE
      port map(D => N_20, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_sampler_clk1x_en_inv_0\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => N_21);
    
    \ReadFIFO_WR_SM.un38_sm_advance_i_NE_6\ : CFG4
      generic map(INIT => x"FFF6")

      port map(A => \consumer_type[4]_net_1\, B => 
        consumer_type4_reg(4), C => un38_sm_advance_i_NE_3, D => 
        un38_sm_advance_i_5, Y => un38_sm_advance_i_NE_6);
    
    \rx_packet_length[2]\ : SLE
      port map(D => \rx_packet_length_13[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rx_packet_length[2]_net_1\);
    
    \rx_byte_cntr_lm_0[9]\ : CFG2
      generic map(INIT => x"4")

      port map(A => un1_iRX_EarlyTerm_0_sqmuxa, B => 
        \rx_byte_cntr_s[9]\, Y => \rx_byte_cntr_lm[9]\);
    
    \rx_fifo_din_d2[0]\ : SLE
      port map(D => N_2, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_sampler_clk1x_en_inv_0\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => N_3);
    
    un56_sm_advance_i_cry_1_0 : ARI1
      generic map(INIT => x"511FF")

      port map(A => N_657_mux, B => \un15[7]\, C => \un15[8]\, D
         => GND_net_1, FCI => un56_sm_advance_i_cry_0, S => 
        \un56_sm_advance_i_i[10]\, Y => OPEN, FCO => 
        un56_sm_advance_i_cry_1);
    
    \rx_packet_length_ret_1[8]\ : SLE
      port map(D => \un65_sm_advance_i_i[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \un65_sm_advance_i[1]\);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_8\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[8]_net_1\, B => 
        \un65_sm_advance_i[4]\, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_7, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_8);
    
    \SM_advancebit_cntr[1]\ : SLE
      port map(D => N_121, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => un9_rst_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SM_advancebit_cntr[1]_net_1\);
    
    rx_byte_cntr_s_916 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rx_byte_cntr[0]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => 
        OPEN, Y => OPEN, FCO => rx_byte_cntr_s_916_FCO);
    
    \rx_packet_length_ret[3]\ : SLE
      port map(D => \un56_sm_advance_i_i[8]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \un56_sm_advance_i[8]\);
    
    \bit_cntr[1]\ : SLE
      port map(D => N_116, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => un16_rst_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \bit_cntr[1]_net_1\);
    
    \ReadFIFO_WR_STATE_ns[6]\ : CFG4
      generic map(INIT => x"0CAA")

      port map(A => \un15[3]\, B => \un15[5]\, C => 
        \un58_sm_advance_i_0_data_tmp[5]\, D => 
        \un1_sampler_clk1x_en_inv_0\, Y => 
        \ReadFIFO_WR_STATE_ns[6]_net_1\);
    
    un65_sm_advance_i_cry_1_0 : ARI1
      generic map(INIT => x"5EE00")

      port map(A => N_657_mux, B => \un15[7]\, C => \un15[8]\, D
         => GND_net_1, FCI => un65_sm_advance_i_cry_0, S => 
        \un65_sm_advance_i_i[10]\, Y => OPEN, FCO => 
        un65_sm_advance_i_cry_1);
    
    \rx_byte_cntr[9]\ : SLE
      port map(D => \rx_byte_cntr_lm[9]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => rx_byte_cntre, ALn => RESET_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \rx_byte_cntr[9]_net_1\);
    
    \ReadFIFO_WR_STATE_ns_a2[5]\ : CFG2
      generic map(INIT => x"8")

      port map(A => sampler_clk1x_en, B => \un15[1]\, Y => N_315);
    
    \un1_rx_fifo_din_d3[1]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \RX_FIFO_DIN_pipe[1]\, B => 
        \rx_crc_HighByte_en\, Y => \un1_rx_fifo_din_d3[1]_net_1\);
    
    \rx_packet_length_RNIMK731[9]\ : CFG4
      generic map(INIT => x"CCAC")

      port map(A => RX_FIFO_DIN(1), B => 
        \rx_packet_length[9]_net_1\, C => 
        \un1_sampler_clk1x_en_inv_0\, D => \un15[7]\, Y => 
        N_650_mux);
    
    \rx_packet_length_RNICKTA1[6]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => RX_FIFO_DIN(6), B => N_299, C => 
        \rx_packet_length[6]_net_1\, Y => N_653_mux);
    
    \rx_crc_data_store[13]\ : SLE
      port map(D => \RX_FIFO_DIN_pipe[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => rx_crc_data_store_151, ALn => 
        RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[13]_net_1\);
    
    \rx_crc_data_store[0]\ : SLE
      port map(D => \un1_rx_fifo_din_d3[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_sampler_clk1x_en_inv_i, 
        ALn => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[0]_net_1\);
    
    \rx_byte_cntr_s[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rx_byte_cntr[11]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \rx_byte_cntr_cry[10]_net_1\, S => 
        \rx_byte_cntr_s[11]_net_1\, Y => OPEN, FCO => OPEN);
    
    \rx_byte_cntr_lm_0[10]\ : CFG2
      generic map(INIT => x"4")

      port map(A => un1_iRX_EarlyTerm_0_sqmuxa, B => 
        \rx_byte_cntr_s[10]\, Y => \rx_byte_cntr_lm[10]\);
    
    \ReadFIFO_WR_SM.un1_sampler_clk1x_en_0_I_15\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \rx_crc_data_store[5]_net_1\, B => 
        \rx_crc_data_calc[4]\, C => \rx_crc_data_calc[5]\, D => 
        \rx_crc_data_store[4]_net_1\, FCI => 
        \un1_sampler_clk1x_en_0_data_tmp[1]\, S => OPEN, Y => 
        OPEN, FCO => \un1_sampler_clk1x_en_0_data_tmp[2]\);
    
    un65_sm_advance_i_cry_8_0 : ARI1
      generic map(INIT => x"511FF")

      port map(A => N_650_mux, B => \un15[7]\, C => \un15[8]\, D
         => GND_net_1, FCI => un65_sm_advance_i_cry_7, S => 
        \un65_sm_advance_i_i[3]\, Y => OPEN, FCO => 
        un65_sm_advance_i_cry_8);
    
    \ReadFIFO_WR_SM.un35_sm_advance_i_NE_0\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type3_reg(1), B => 
        consumer_type3_reg(0), C => \consumer_type[1]_net_1\, D
         => \consumer_type[0]_net_1\, Y => un35_sm_advance_i_NE_0);
    
    un56_sm_advance_i_cry_2_0 : ARI1
      generic map(INIT => x"511FF")

      port map(A => N_656_mux, B => \un15[7]\, C => \un15[8]\, D
         => GND_net_1, FCI => un56_sm_advance_i_cry_1, S => 
        \un56_sm_advance_i_i[9]\, Y => OPEN, FCO => 
        un56_sm_advance_i_cry_2);
    
    \rx_packet_length_ret_1[5]\ : SLE
      port map(D => \un65_sm_advance_i_i[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \un65_sm_advance_i[4]\);
    
    \consumer_type[1]\ : SLE
      port map(D => \consumer_type_12[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_12, ALn
         => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type[1]_net_1\);
    
    \bit_cntr_RNO[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => N_221, B => \bit_cntr[0]_net_1\, Y => N_44_i);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_4\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[4]_net_1\, B => 
        \un65_sm_advance_i[8]\, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_3, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_4);
    
    \rx_fifo_din_d1[4]\ : SLE
      port map(D => RX_FIFO_DIN(4), CLK => CommsFPGA_CCC_0_GL0, 
        EN => \un1_sampler_clk1x_en_inv_0\, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => N_14);
    
    rx_CRC_error_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => \un1_sampler_clk1x_en_0_data_tmp[7]\, B => 
        \un15[1]\, Y => N_676);
    
    \rx_byte_cntr_lm_0[11]\ : CFG2
      generic map(INIT => x"4")

      port map(A => un1_iRX_EarlyTerm_0_sqmuxa, B => 
        \rx_byte_cntr_s[11]_net_1\, Y => \rx_byte_cntr_lm[11]\);
    
    \rx_byte_cntr_lm_0[7]\ : CFG2
      generic map(INIT => x"4")

      port map(A => un1_iRX_EarlyTerm_0_sqmuxa, B => 
        \rx_byte_cntr_s[7]\, Y => \rx_byte_cntr_lm[7]\);
    
    \rx_fifo_din_d2[1]\ : SLE
      port map(D => N_5, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_sampler_clk1x_en_inv_0\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => N_6);
    
    \rx_byte_cntr_lm_0[3]\ : CFG2
      generic map(INIT => x"4")

      port map(A => un1_iRX_EarlyTerm_0_sqmuxa, B => 
        \rx_byte_cntr_s[3]\, Y => \rx_byte_cntr_lm[3]\);
    
    \un1_rx_fifo_din_d3[7]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \RX_FIFO_DIN_pipe[7]\, B => 
        \rx_crc_HighByte_en\, Y => \un1_rx_fifo_din_d3[7]_net_1\);
    
    \ReadFIFO_WR_STATE[0]\ : SLE
      port map(D => \ReadFIFO_WR_STATE_ns[9]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \un15[0]\);
    
    \ReadFIFO_WR_STATE[6]\ : SLE
      port map(D => \ReadFIFO_WR_STATE_ns[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \un15[7]\);
    
    un56_sm_advance_i_cry_8_0 : ARI1
      generic map(INIT => x"511FF")

      port map(A => N_650_mux, B => \un15[7]\, C => \un15[8]\, D
         => GND_net_1, FCI => un56_sm_advance_i_cry_7, S => 
        \un56_sm_advance_i_i[3]\, Y => OPEN, FCO => 
        un56_sm_advance_i_cry_8);
    
    \rx_fifo_din_d2[5]\ : SLE
      port map(D => N_17, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_sampler_clk1x_en_inv_0\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => N_18);
    
    \rx_fifo_din_d1[3]\ : SLE
      port map(D => RX_FIFO_DIN(3), CLK => CommsFPGA_CCC_0_GL0, 
        EN => \un1_sampler_clk1x_en_inv_0\, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => N_11);
    
    \un1_rx_fifo_din_d3[0]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \RX_FIFO_DIN_pipe[0]\, B => 
        \rx_crc_HighByte_en\, Y => \un1_rx_fifo_din_d3[0]_net_1\);
    
    un1_iRX_EarlyTerm_1_sqmuxa_1_0 : CFG4
      generic map(INIT => x"F0F2")

      port map(A => N_321, B => \un15[9]\, C => 
        \un1_sampler_clk1x_en_inv_0\, D => N_314, Y => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0\);
    
    \rx_byte_cntr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rx_byte_cntr[2]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \rx_byte_cntr_cry[1]_net_1\, S => \rx_byte_cntr_s[2]\, Y
         => OPEN, FCO => \rx_byte_cntr_cry[2]_net_1\);
    
    \ReadFIFO_WR_SM.un40_sm_advance_i_1\ : CFG4
      generic map(INIT => x"EEE0")

      port map(A => un35_sm_advance_i_NE_7, B => 
        un35_sm_advance_i_NE_6, C => un29_sm_advance_i_NE_7, D
         => un29_sm_advance_i_NE_6, Y => un40_sm_advance_i_1);
    
    \ReadFIFO_WRITE_PROC.un16_rst_0_RNIS9M7\ : CFG1
      generic map(INIT => "01")

      port map(A => un9_rst, Y => un9_rst_i);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_9\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[9]_net_1\, B => 
        \un65_sm_advance_i[3]\, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_8, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_9);
    
    \CoreAPB3_0_APBmslave0_PRDATA_m[5]\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        CoreAPB3_0_APBmslave0_PRDATA(5), Y => 
        CoreAPB3_0_APBmslave0_PRDATA_m(5));
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_7\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[7]_net_1\, B => 
        \un65_sm_advance_i[5]\, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_6, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_7);
    
    \ReadFIFO_WR_SM.consumer_type_12[6]\ : CFG4
      generic map(INIT => x"E4A0")

      port map(A => \un15[9]\, B => consumer_type_0_sqmuxa, C => 
        \consumer_type[6]_net_1\, D => RX_FIFO_DIN(4), Y => 
        \consumer_type_12[6]\);
    
    \rx_byte_cntr[8]\ : SLE
      port map(D => \rx_byte_cntr_lm[8]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => rx_byte_cntre, ALn => RESET_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \rx_byte_cntr[8]_net_1\);
    
    \rx_byte_cntr[2]\ : SLE
      port map(D => \rx_byte_cntr_lm[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => rx_byte_cntre, ALn => RESET_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \rx_byte_cntr[2]_net_1\);
    
    \ReadFIFO_WR_SM.un32_sm_advance_i_NE_1\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type2_reg(3), B => 
        consumer_type2_reg(2), C => \consumer_type[3]_net_1\, D
         => \consumer_type[2]_net_1\, Y => un32_sm_advance_i_NE_1);
    
    \ReadFIFO_WR_SM.un35_sm_advance_i_NE_7\ : CFG3
      generic map(INIT => x"FE")

      port map(A => un35_sm_advance_i_NE_4, B => 
        un35_sm_advance_i_NE_1, C => un35_sm_advance_i_NE_0, Y
         => un35_sm_advance_i_NE_7);
    
    \rx_packet_length[7]\ : SLE
      port map(D => \rx_packet_length_13[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rx_packet_length[7]_net_1\);
    
    \rx_byte_cntr_lm_0[2]\ : CFG2
      generic map(INIT => x"4")

      port map(A => un1_iRX_EarlyTerm_0_sqmuxa, B => 
        \rx_byte_cntr_s[2]\, Y => \rx_byte_cntr_lm[2]\);
    
    \RX_FIFO_TxColDetDis_wr_en\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \iRX_FIFO_wr_en\, B => sampler_clk1x_en, C
         => \RX_InProcess_d1\, D => tx_col_detect_en, Y => 
        RX_FIFO_TxColDetDis_wr_en);
    
    \ReadFIFO_WR_SM.consumer_type_12[0]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => RX_FIFO_DIN(6), B => \consumer_type[0]_net_1\, 
        C => consumer_type_12_sn_N_2, D => N_661, Y => 
        \consumer_type_12[0]\);
    
    \ReadFIFO_WR_SM.un58_sm_advance_i_0_I_15\ : ARI1
      generic map(INIT => x"68241")

      port map(A => \un56_sm_advance_i[10]\, B => 
        \rx_byte_cntr[2]_net_1\, C => \rx_byte_cntr[3]_net_1\, D
         => \un56_sm_advance_i[9]\, FCI => 
        \un58_sm_advance_i_0_data_tmp[0]\, S => OPEN, Y => OPEN, 
        FCO => \un58_sm_advance_i_0_data_tmp[1]\);
    
    \ReadFIFO_WR_STATE_ns_i_a3_0[0]\ : CFG4
      generic map(INIT => x"0040")

      port map(A => \un15[4]\, B => packet_avail, C => 
        \un1_sampler_clk1x_en_inv_0\, D => \un15[0]\, Y => N_294);
    
    un65_sm_advance_i_s_9 : ARI1
      generic map(INIT => x"47700")

      port map(A => VCC_net_1, B => un1_ReadFIFO_WR_STATE_6_i, C
         => N_649_mux, D => GND_net_1, FCI => 
        un65_sm_advance_i_s_9_922_FCO, S => 
        \un65_sm_advance_i_i[2]\, Y => OPEN, FCO => OPEN);
    
    RX_InProcess : SLE
      port map(D => N_314, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_InProcess\);
    
    un1_sampler_clk1x_en_inv_0 : CFG2
      generic map(INIT => x"8")

      port map(A => sampler_clk1x_en, B => \SM_advance_i\, Y => 
        \un1_sampler_clk1x_en_inv_0\);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_3\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[3]_net_1\, B => 
        \un65_sm_advance_i[9]\, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_2, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_3);
    
    \ReadFIFO_WR_SM.consumer_type_12[5]\ : CFG4
      generic map(INIT => x"E4A0")

      port map(A => \un15[9]\, B => consumer_type_0_sqmuxa, C => 
        \consumer_type[5]_net_1\, D => RX_FIFO_DIN(3), Y => 
        \consumer_type_12[5]\);
    
    \rx_fifo_din_d1[1]\ : SLE
      port map(D => RX_FIFO_DIN(1), CLK => CommsFPGA_CCC_0_GL0, 
        EN => \un1_sampler_clk1x_en_inv_0\, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => N_5);
    
    \ReadFIFO_WR_SM.un38_sm_advance_i_NE_3\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type4_reg(7), B => 
        consumer_type4_reg(6), C => \consumer_type[7]_net_1\, D
         => \consumer_type[6]_net_1\, Y => un38_sm_advance_i_NE_3);
    
    un56_sm_advance_i_s_9 : ARI1
      generic map(INIT => x"47700")

      port map(A => VCC_net_1, B => un1_ReadFIFO_WR_STATE_6_i, C
         => N_649_mux, D => GND_net_1, FCI => 
        un56_sm_advance_i_s_9_921_FCO, S => 
        \un56_sm_advance_i_i[2]\, Y => OPEN, FCO => OPEN);
    
    \rx_fifo_din_d3[5]\ : SLE
      port map(D => N_18, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_sampler_clk1x_en_inv_0\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN_pipe[5]\);
    
    rx_crc_reset : CFG2
      generic map(INIT => x"1")

      port map(A => \rx_end_rst\, B => RESET, Y => \rx_crc_reset\);
    
    rx_crc_data_store_151_0 : CFG2
      generic map(INIT => x"8")

      port map(A => \un1_sampler_clk1x_en_inv_0\, B => 
        \rx_crc_HighByte_en\, Y => rx_crc_data_store_151);
    
    un65_sm_advance_i_cry_0_0 : ARI1
      generic map(INIT => x"511FF")

      port map(A => N_658_mux, B => \un15[7]\, C => \un15[8]\, D
         => GND_net_1, FCI => GND_net_1, S => OPEN, Y => OPEN, 
        FCO => un65_sm_advance_i_cry_0);
    
    \rx_fifo_din_d2[2]\ : SLE
      port map(D => N_8, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_sampler_clk1x_en_inv_0\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => N_9);
    
    \rx_byte_cntr[0]\ : SLE
      port map(D => \rx_byte_cntr_lm[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => rx_byte_cntre, ALn => RESET_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \rx_byte_cntr[0]_net_1\);
    
    \bit_cntr_RNO[2]\ : CFG4
      generic map(INIT => x"6AAA")

      port map(A => \bit_cntr[2]_net_1\, B => \bit_cntr[1]_net_1\, 
        C => \bit_cntr[0]_net_1\, D => N_221, Y => N_117);
    
    \rx_packet_length[0]\ : SLE
      port map(D => \rx_packet_length_13[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rx_packet_length[0]_net_1\);
    
    \ReadFIFO_WR_SM.un29_sm_advance_i_NE_3\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type1_reg(7), B => 
        consumer_type1_reg(6), C => \consumer_type[7]_net_1\, D
         => \consumer_type[6]_net_1\, Y => un29_sm_advance_i_NE_3);
    
    \CoreAPB3_0_APBmslave0_PRDATA_m[0]\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        CoreAPB3_0_APBmslave0_PRDATA(0), Y => 
        CoreAPB3_0_APBmslave0_PRDATA_m(0));
    
    \un1_rx_fifo_din_d3[2]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \RX_FIFO_DIN_pipe[2]\, B => 
        \rx_crc_HighByte_en\, Y => \un1_rx_fifo_din_d3[2]_net_1\);
    
    \rx_packet_length_13[4]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_655_mux, B => un1_ReadFIFO_WR_STATE_6_i, Y
         => \rx_packet_length_13[4]_net_1\);
    
    \rx_crc_data_store[11]\ : SLE
      port map(D => \RX_FIFO_DIN_pipe[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => rx_crc_data_store_151, ALn => 
        RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[11]_net_1\);
    
    \ReadFIFO_WR_SM.consumer_type_12[2]\ : CFG4
      generic map(INIT => x"E4A0")

      port map(A => \un15[9]\, B => consumer_type_0_sqmuxa, C => 
        \consumer_type[2]_net_1\, D => RX_FIFO_DIN(0), Y => 
        \consumer_type_12[2]\);
    
    \rx_packet_length_RNIEMTA1[7]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => RX_FIFO_DIN(7), B => N_299, C => 
        \rx_packet_length[7]_net_1\, Y => N_652_mux);
    
    un1_ReadFIFO_WR_STATE_12_0 : CFG3
      generic map(INIT => x"54")

      port map(A => N_314, B => \un1_sampler_clk1x_en_inv_0\, C
         => N_321, Y => un1_ReadFIFO_WR_STATE_12);
    
    \rx_byte_cntr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rx_byte_cntr[1]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        rx_byte_cntr_s_916_FCO, S => \rx_byte_cntr_s[1]\, Y => 
        OPEN, FCO => \rx_byte_cntr_cry[1]_net_1\);
    
    \bit_cntr_RNO[1]\ : CFG3
      generic map(INIT => x"6A")

      port map(A => \bit_cntr[1]_net_1\, B => \bit_cntr[0]_net_1\, 
        C => N_221, Y => N_116);
    
    \ReadFIFO_WR_SM.consumer_type_12[1]\ : CFG4
      generic map(INIT => x"0A0C")

      port map(A => RX_FIFO_DIN(7), B => \consumer_type[1]_net_1\, 
        C => consumer_type_12_sn_N_2, D => N_661, Y => 
        \consumer_type_12[1]\);
    
    \rx_packet_length_13[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_658_mux, B => un1_ReadFIFO_WR_STATE_6_i, Y
         => \rx_packet_length_13[1]_net_1\);
    
    rx_end_rst_RNO : CFG2
      generic map(INIT => x"4")

      port map(A => N_320, B => idle_line, Y => N_279_i);
    
    \ReadFIFO_WR_SM.consumer_type_12[7]\ : CFG4
      generic map(INIT => x"E4A0")

      port map(A => \un15[9]\, B => consumer_type_0_sqmuxa, C => 
        \consumer_type[7]_net_1\, D => RX_FIFO_DIN(5), Y => 
        \consumer_type_12[7]\);
    
    un56_sm_advance_i_cry_4_0 : ARI1
      generic map(INIT => x"511FF")

      port map(A => N_654_mux, B => \un15[7]\, C => \un15[8]\, D
         => GND_net_1, FCI => un56_sm_advance_i_cry_3, S => 
        \un56_sm_advance_i_i[7]\, Y => OPEN, FCO => 
        un56_sm_advance_i_cry_4);
    
    \rx_crc_data_store[10]\ : SLE
      port map(D => \RX_FIFO_DIN_pipe[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => rx_crc_data_store_151, ALn => 
        RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[10]_net_1\);
    
    \rx_packet_length_ret[7]\ : SLE
      port map(D => \un56_sm_advance_i_i[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \un56_sm_advance_i[4]\);
    
    \rx_byte_cntr_lm_0[4]\ : CFG2
      generic map(INIT => x"4")

      port map(A => un1_iRX_EarlyTerm_0_sqmuxa, B => 
        \rx_byte_cntr_s[4]\, Y => \rx_byte_cntr_lm[4]\);
    
    \rx_byte_cntr[10]\ : SLE
      port map(D => \rx_byte_cntr_lm[10]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => rx_byte_cntre, ALn => RESET_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \rx_byte_cntr[10]_net_1\);
    
    SM_advance_i_0_sqmuxa_i : CFG2
      generic map(INIT => x"8")

      port map(A => sampler_clk1x_en, B => packet_avail, Y => 
        N_221);
    
    \rx_packet_length_ret_1[2]\ : SLE
      port map(D => \un65_sm_advance_i_i[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \un65_sm_advance_i[7]\);
    
    un65_sm_advance_i_cry_5_0 : ARI1
      generic map(INIT => x"511FF")

      port map(A => N_653_mux, B => \un15[7]\, C => \un15[8]\, D
         => GND_net_1, FCI => un65_sm_advance_i_cry_4, S => 
        \un65_sm_advance_i_i[6]\, Y => OPEN, FCO => 
        un65_sm_advance_i_cry_5);
    
    \SM_advancebit_cntr_RNO[2]\ : CFG4
      generic map(INIT => x"6AAA")

      port map(A => \SM_advancebit_cntr[2]_net_1\, B => 
        \SM_advancebit_cntr[1]_net_1\, C => 
        \SM_advancebit_cntr[0]_net_1\, D => N_221, Y => N_122);
    
    \rx_crc_data_store[7]\ : SLE
      port map(D => \un1_rx_fifo_din_d3[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_sampler_clk1x_en_inv_i, 
        ALn => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[7]_net_1\);
    
    \CoreAPB3_0_APBmslave0_PRDATA_m[6]\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        CoreAPB3_0_APBmslave0_PRDATA(6), Y => 
        CoreAPB3_0_APBmslave0_PRDATA_m(6));
    
    \ReadFIFO_WR_SM.consumer_type_12[3]\ : CFG4
      generic map(INIT => x"E4A0")

      port map(A => \un15[9]\, B => consumer_type_0_sqmuxa, C => 
        \consumer_type[3]_net_1\, D => RX_FIFO_DIN(1), Y => 
        \consumer_type_12[3]\);
    
    \ReadFIFO_WR_SM.un38_sm_advance_i_5\ : CFG2
      generic map(INIT => x"6")

      port map(A => \consumer_type[5]_net_1\, B => 
        consumer_type4_reg(5), Y => un38_sm_advance_i_5);
    
    \rx_fifo_din_d1[7]\ : SLE
      port map(D => RX_FIFO_DIN(7), CLK => CommsFPGA_CCC_0_GL0, 
        EN => \un1_sampler_clk1x_en_inv_0\, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => N_23);
    
    \ReadFIFO_WR_STATE_ns_a3_0_0[3]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \un1_sampler_clk1x_en_inv_0\, B => \un15[8]\, 
        Y => \ReadFIFO_WR_STATE_ns_a3_0_0[3]_net_1\);
    
    \CoreAPB3_0_APBmslave0_PREADY_i_m_i\ : CFG2
      generic map(INIT => x"D")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        CoreAPB3_0_APBmslave0_PREADY, Y => 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i);
    
    \rx_byte_cntr[6]\ : SLE
      port map(D => \rx_byte_cntr_lm[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => rx_byte_cntre, ALn => RESET_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \rx_byte_cntr[6]_net_1\);
    
    consumer_type_0_sqmuxa_0_a3_RNIK0S8 : CFG2
      generic map(INIT => x"1")

      port map(A => consumer_type_0_sqmuxa, B => \un15[9]\, Y => 
        consumer_type_12_sn_N_2);
    
    \rx_packet_length_RNI2ATA1[1]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => RX_FIFO_DIN(1), B => N_299, C => 
        \rx_packet_length[1]_net_1\, Y => N_658_mux);
    
    rx_crc_LowByte_en_RNIK30V : CFG3
      generic map(INIT => x"A8")

      port map(A => \un1_sampler_clk1x_en_inv_0\, B => 
        \rx_crc_HighByte_en\, C => \RX_FIFO_DIN_pipe[8]\, Y => 
        un1_sampler_clk1x_en_inv_i);
    
    \ReadFIFO_WR_STATE_ns_a3_0_1_0[3]\ : CFG4
      generic map(INIT => x"0CAC")

      port map(A => \un15[8]\, B => \un15[7]\, C => 
        \un1_sampler_clk1x_en_inv_0\, D => un40_sm_advance_i_1, Y
         => \ReadFIFO_WR_STATE_ns_a3_0_1_0[3]_net_1\);
    
    \ReadFIFO_WR_SM.un35_sm_advance_i_NE_1\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type3_reg(3), B => 
        consumer_type3_reg(2), C => \consumer_type[3]_net_1\, D
         => \consumer_type[2]_net_1\, Y => un35_sm_advance_i_NE_1);
    
    \ReadFIFO_WR_SM.un1_sampler_clk1x_en_0_I_39\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \rx_crc_data_store[13]_net_1\, B => 
        \rx_crc_data_calc[12]\, C => \rx_crc_data_calc[13]\, D
         => \rx_crc_data_store[12]_net_1\, FCI => 
        \un1_sampler_clk1x_en_0_data_tmp[5]\, S => OPEN, Y => 
        OPEN, FCO => \un1_sampler_clk1x_en_0_data_tmp[6]\);
    
    \CoreAPB3_0_APBmslave0_PRDATA_m[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        CoreAPB3_0_APBmslave0_PRDATA(1), Y => 
        CoreAPB3_0_APBmslave0_PRDATA_m(1));
    
    \rx_packet_length_ret_1[4]\ : SLE
      port map(D => \un65_sm_advance_i_i[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \un65_sm_advance_i[5]\);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_10\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[10]_net_1\, B => 
        \un65_sm_advance_i[2]\, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_9, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_10);
    
    \rx_packet_length_13[9]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_650_mux, B => un1_ReadFIFO_WR_STATE_6_i, Y
         => \rx_packet_length_13[9]_net_1\);
    
    \ReadFIFO_WR_STATE_ns_0[5]\ : CFG4
      generic map(INIT => x"F444")

      port map(A => idle_line, B => \un15[4]\, C => 
        \un1_sampler_clk1x_en_0_data_tmp[7]\, D => N_315, Y => 
        \ReadFIFO_WR_STATE_ns_0[5]_net_1\);
    
    \ReadFIFO_WR_STATE[3]\ : SLE
      port map(D => \ReadFIFO_WR_STATE_ns[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \un15[3]\);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_5\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[5]_net_1\, B => 
        \un65_sm_advance_i[7]\, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_4, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_5);
    
    \ReadFIFO_WRITE_PROC.un16_rst_0\ : CFG3
      generic map(INIT => x"EF")

      port map(A => RESET, B => \RX_EarlyTerm\, C => clk1x_enable, 
        Y => un9_rst);
    
    \ReadFIFO_WR_SM.un29_sm_advance_i_5\ : CFG2
      generic map(INIT => x"6")

      port map(A => \consumer_type[5]_net_1\, B => 
        consumer_type1_reg(5), Y => un29_sm_advance_i_5);
    
    \ReadFIFO_WR_STATE[1]\ : SLE
      port map(D => \ReadFIFO_WR_STATE_ns[8]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \un15[1]\);
    
    \ReadFIFO_WR_SM.un29_sm_advance_i_NE_0\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type1_reg(1), B => 
        consumer_type1_reg(0), C => \consumer_type[1]_net_1\, D
         => \consumer_type[0]_net_1\, Y => un29_sm_advance_i_NE_0);
    
    un1_iRX_EarlyTerm_0_sqmuxa_0 : CFG4
      generic map(INIT => x"FFEC")

      port map(A => \un15[2]\, B => N_315, C => 
        \un1_sampler_clk1x_en_inv_0\, D => N_308, Y => 
        un1_iRX_EarlyTerm_0_sqmuxa);
    
    \ReadFIFO_WR_STATE[8]\ : SLE
      port map(D => \ReadFIFO_WR_STATE_ns[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \un15[9]\);
    
    \rx_crc_data_store[9]\ : SLE
      port map(D => \RX_FIFO_DIN_pipe[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => rx_crc_data_store_151, ALn => 
        RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[9]_net_1\);
    
    \rx_packet_length_13[2]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_657_mux, B => un1_ReadFIFO_WR_STATE_6_i, Y
         => \rx_packet_length_13[2]_net_1\);
    
    \rx_packet_length_RNIAITA1[5]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => RX_FIFO_DIN(5), B => N_299, C => 
        \rx_packet_length[5]_net_1\, Y => N_654_mux);
    
    \ReadFIFO_WR_SM.un32_sm_advance_i_NE_5\ : CFG4
      generic map(INIT => x"FFF6")

      port map(A => \consumer_type[0]_net_1\, B => 
        consumer_type2_reg(0), C => un32_sm_advance_i_NE_1, D => 
        un32_sm_advance_i_1, Y => un32_sm_advance_i_NE_5);
    
    un65_sm_advance_i_cry_2_0 : ARI1
      generic map(INIT => x"511FF")

      port map(A => N_656_mux, B => \un15[7]\, C => \un15[8]\, D
         => GND_net_1, FCI => un65_sm_advance_i_cry_1, S => 
        \un65_sm_advance_i_i[9]\, Y => OPEN, FCO => 
        un65_sm_advance_i_cry_2);
    
    \un1_rx_fifo_din_d3[6]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \RX_FIFO_DIN_pipe[6]\, B => 
        \rx_crc_HighByte_en\, Y => \un1_rx_fifo_din_d3[6]_net_1\);
    
    \rx_crc_data_store[4]\ : SLE
      port map(D => \un1_rx_fifo_din_d3[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_sampler_clk1x_en_inv_i, 
        ALn => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[4]_net_1\);
    
    \rx_byte_cntr[5]\ : SLE
      port map(D => \rx_byte_cntr_lm[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => rx_byte_cntre, ALn => RESET_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \rx_byte_cntr[5]_net_1\);
    
    un56_sm_advance_i_cry_9_ma : CFG2
      generic map(INIT => x"8")

      port map(A => N_649_mux, B => un1_ReadFIFO_WR_STATE_6_i, Y
         => \un56_sm_advance_i_cry_9_ma\);
    
    \rx_fifo_din_d2[7]\ : SLE
      port map(D => N_23, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_sampler_clk1x_en_inv_0\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => N_24);
    
    \ReadFIFO_WR_SM.un35_sm_advance_i_NE_3\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type3_reg(7), B => 
        consumer_type3_reg(6), C => \consumer_type[7]_net_1\, D
         => \consumer_type[6]_net_1\, Y => un35_sm_advance_i_NE_3);
    
    \un1_rx_fifo_din_d3[3]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \RX_FIFO_DIN_pipe[3]\, B => 
        \rx_crc_HighByte_en\, Y => \un1_rx_fifo_din_d3[3]_net_1\);
    
    \ReadFIFO_WRITE_PROC.un5_packet_avail\ : CFG3
      generic map(INIT => x"80")

      port map(A => \bit_cntr[2]_net_1\, B => \bit_cntr[1]_net_1\, 
        C => \bit_cntr[0]_net_1\, Y => un5_packet_avail);
    
    rx_packet_complt_1_sqmuxa : CFG3
      generic map(INIT => x"08")

      port map(A => \un15[0]\, B => idle_line, C => 
        tx_col_detect_en, Y => \rx_packet_complt_1_sqmuxa\);
    
    \ReadFIFO_WR_SM.un32_sm_advance_i_NE_4\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type2_reg(9), B => 
        consumer_type2_reg(8), C => \consumer_type[9]_net_1\, D
         => \consumer_type[8]_net_1\, Y => un32_sm_advance_i_NE_4);
    
    \rx_packet_length_ret[10]\ : SLE
      port map(D => \un56_sm_advance_i_i[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \un56_sm_advance_i[1]\);
    
    \rx_fifo_din_d3[1]\ : SLE
      port map(D => N_6, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_sampler_clk1x_en_inv_0\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN_pipe[1]\);
    
    \ReadFIFO_WR_STATE_ns[1]\ : CFG3
      generic map(INIT => x"F2")

      port map(A => \un15[9]\, B => \un1_sampler_clk1x_en_inv_0\, 
        C => consumer_type_0_sqmuxa, Y => 
        \ReadFIFO_WR_STATE_ns[1]_net_1\);
    
    rx_crc_gen_3_sqmuxa : CFG3
      generic map(INIT => x"20")

      port map(A => \un15[5]\, B => un67_sm_advance_i, C => 
        \un58_sm_advance_i_0_data_tmp[5]\, Y => 
        \rx_crc_gen_3_sqmuxa\);
    
    \rx_crc_data_store[2]\ : SLE
      port map(D => \un1_rx_fifo_din_d3[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_sampler_clk1x_en_inv_i, 
        ALn => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[2]_net_1\);
    
    \ReadFIFO_WR_SM.un29_sm_advance_i_NE_1\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type1_reg(3), B => 
        consumer_type1_reg(2), C => \consumer_type[3]_net_1\, D
         => \consumer_type[2]_net_1\, Y => un29_sm_advance_i_NE_1);
    
    \rx_packet_length_ret_1[1]\ : SLE
      port map(D => \un65_sm_advance_i_i[8]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \un65_sm_advance_i[8]\);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_2\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[2]_net_1\, B => 
        \un65_sm_advance_i[10]\, C => GND_net_1, D => GND_net_1, 
        FCI => un67_sm_advance_i_cry_1, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_2);
    
    \rx_packet_length_ret_1[7]\ : SLE
      port map(D => \un65_sm_advance_i_i[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \un65_sm_advance_i[2]\);
    
    \rx_packet_length[4]\ : SLE
      port map(D => \rx_packet_length_13[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rx_packet_length[4]_net_1\);
    
    un65_sm_advance_i_cry_7_0 : ARI1
      generic map(INIT => x"511FF")

      port map(A => N_651_mux, B => \un15[7]\, C => \un15[8]\, D
         => GND_net_1, FCI => un65_sm_advance_i_cry_6, S => 
        \un65_sm_advance_i_i[4]\, Y => OPEN, FCO => 
        un65_sm_advance_i_cry_7);
    
    \ReadFIFO_WR_STATE_RNIDMB2[7]\ : CFG2
      generic map(INIT => x"E")

      port map(A => \un15[7]\, B => \un15[8]\, Y => 
        un1_ReadFIFO_WR_STATE_6_i);
    
    \rx_packet_length[1]\ : SLE
      port map(D => \rx_packet_length_13[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rx_packet_length[1]_net_1\);
    
    \rx_byte_cntr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rx_byte_cntr[5]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \rx_byte_cntr_cry[4]_net_1\, S => \rx_byte_cntr_s[5]\, Y
         => OPEN, FCO => \rx_byte_cntr_cry[5]_net_1\);
    
    \rx_fifo_din_d2[4]\ : SLE
      port map(D => N_14, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_sampler_clk1x_en_inv_0\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => N_15);
    
    rx_crc_reset_RNI34TD : CLKINT
      port map(A => \rx_crc_reset\, Y => rx_crc_reset_i);
    
    \rx_fifo_din_d2[3]\ : SLE
      port map(D => N_11, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_sampler_clk1x_en_inv_0\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => N_12);
    
    \consumer_type[5]\ : SLE
      port map(D => \consumer_type_12[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_12, ALn
         => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type[5]_net_1\);
    
    un1_ReadFIFO_WR_STATE_15 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \un15[10]\, B => \un15[9]\, C => 
        un1_ReadFIFO_WR_STATE_6_i, D => \rx_crc_gen_3_sqmuxa\, Y
         => \un1_ReadFIFO_WR_STATE_15\);
    
    \rx_crc_data_store[14]\ : SLE
      port map(D => \RX_FIFO_DIN_pipe[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => rx_crc_data_store_151, ALn => 
        RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[14]_net_1\);
    
    \ReadFIFO_WR_SM.consumer_type_12[8]\ : CFG4
      generic map(INIT => x"E4A0")

      port map(A => \un15[9]\, B => consumer_type_0_sqmuxa, C => 
        \consumer_type[8]_net_1\, D => RX_FIFO_DIN(6), Y => 
        \consumer_type_12[8]\);
    
    \ReadFIFO_WR_SM.un29_sm_advance_i_NE_6\ : CFG4
      generic map(INIT => x"FFF6")

      port map(A => \consumer_type[4]_net_1\, B => 
        consumer_type1_reg(4), C => un29_sm_advance_i_NE_3, D => 
        un29_sm_advance_i_5, Y => un29_sm_advance_i_NE_6);
    
    \ReadFIFO_WR_SM.un40_sm_advance_i_2\ : CFG4
      generic map(INIT => x"5400")

      port map(A => DRVR_EN_c, B => un38_sm_advance_i_NE_7, C => 
        un38_sm_advance_i_NE_6, D => un33_sm_advance_i, Y => 
        un40_sm_advance_i_2);
    
    \un1_rx_fifo_din_d3[5]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \RX_FIFO_DIN_pipe[5]\, B => 
        \rx_crc_HighByte_en\, Y => \un1_rx_fifo_din_d3[5]_net_1\);
    
    \rx_packet_length_13[8]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_651_mux, B => un1_ReadFIFO_WR_STATE_6_i, Y
         => \rx_packet_length_13[8]_net_1\);
    
    \ReadFIFO_WR_STATE[9]\ : SLE
      port map(D => N_253_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => RESET_i, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \un15[10]\);
    
    \rx_byte_cntr[4]\ : SLE
      port map(D => \rx_byte_cntr_lm[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => rx_byte_cntre, ALn => RESET_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \rx_byte_cntr[4]_net_1\);
    
    \SM_advancebit_cntr[2]\ : SLE
      port map(D => N_122, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => un9_rst_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SM_advancebit_cntr[2]_net_1\);
    
    irx_packet_end_RNO : CFG3
      generic map(INIT => x"FE")

      port map(A => \un15[2]\, B => \un15[1]\, C => \un15[0]\, Y
         => N_689_i);
    
    \consumer_type[0]\ : SLE
      port map(D => \consumer_type_12[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_12, ALn
         => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type[0]_net_1\);
    
    RX_CRC_GEN_INST : CRC16_Generator_1
      port map(RX_FIFO_DIN(7) => RX_FIFO_DIN(7), RX_FIFO_DIN(6)
         => RX_FIFO_DIN(6), RX_FIFO_DIN(5) => RX_FIFO_DIN(5), 
        RX_FIFO_DIN(4) => RX_FIFO_DIN(4), RX_FIFO_DIN(3) => 
        RX_FIFO_DIN(3), RX_FIFO_DIN(2) => RX_FIFO_DIN(2), 
        RX_FIFO_DIN(1) => RX_FIFO_DIN(1), RX_FIFO_DIN(0) => 
        RX_FIFO_DIN(0), rx_crc_data_calc(15) => 
        \rx_crc_data_calc[15]\, rx_crc_data_calc(14) => 
        \rx_crc_data_calc[14]\, rx_crc_data_calc(13) => 
        \rx_crc_data_calc[13]\, rx_crc_data_calc(12) => 
        \rx_crc_data_calc[12]\, rx_crc_data_calc(11) => 
        \rx_crc_data_calc[11]\, rx_crc_data_calc(10) => 
        \rx_crc_data_calc[10]\, rx_crc_data_calc(9) => 
        \rx_crc_data_calc[9]\, rx_crc_data_calc(8) => 
        \rx_crc_data_calc[8]\, rx_crc_data_calc(7) => 
        \rx_crc_data_calc[7]\, rx_crc_data_calc(6) => 
        \rx_crc_data_calc[6]\, rx_crc_data_calc(5) => 
        \rx_crc_data_calc[5]\, rx_crc_data_calc(4) => 
        \rx_crc_data_calc[4]\, rx_crc_data_calc(3) => 
        \rx_crc_data_calc[3]\, rx_crc_data_calc(2) => 
        \rx_crc_data_calc[2]\, rx_crc_data_calc(1) => 
        \rx_crc_data_calc[1]\, rx_crc_data_calc(0) => 
        \rx_crc_data_calc[0]\, rx_crc_gen => \rx_crc_gen\, 
        sampler_clk1x_en => sampler_clk1x_en, iRX_FIFO_wr_en => 
        \iRX_FIFO_wr_en\, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, rx_crc_reset_i => rx_crc_reset_i);
    
    \ReadFIFO_WR_SM.un67_sm_advance_i_cry_0\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \rx_byte_cntr[0]_net_1\, B => 
        \rx_packet_length[0]_net_1\, C => GND_net_1, D => 
        GND_net_1, FCI => GND_net_1, S => OPEN, Y => OPEN, FCO
         => un67_sm_advance_i_cry_0);
    
    \rx_fifo_din_d3[7]\ : SLE
      port map(D => N_24, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_sampler_clk1x_en_inv_0\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN_pipe[7]\);
    
    \rx_packet_length[9]\ : SLE
      port map(D => \rx_packet_length_13[9]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rx_packet_length[9]_net_1\);
    
    \rx_byte_cntr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rx_byte_cntr[6]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \rx_byte_cntr_cry[5]_net_1\, S => \rx_byte_cntr_s[6]\, Y
         => OPEN, FCO => \rx_byte_cntr_cry[6]_net_1\);
    
    un1_ReadFIFO_WR_STATE_14_0_o2_RNIGH1Q : CFG4
      generic map(INIT => x"EEEC")

      port map(A => \un1_sampler_clk1x_en_inv_0\, B => 
        un1_iRX_EarlyTerm_0_sqmuxa, C => \un15[7]\, D => N_276, Y
         => rx_byte_cntre);
    
    un1_ReadFIFO_WR_STATE_14_0 : CFG4
      generic map(INIT => x"00CE")

      port map(A => N_321, B => \un1_sampler_clk1x_en_inv_0\, C
         => \un15[9]\, D => N_276, Y => un1_ReadFIFO_WR_STATE_14);
    
    \rx_packet_length_RNI6ETA1[3]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => RX_FIFO_DIN(3), B => N_299, C => 
        \rx_packet_length[3]_net_1\, Y => N_656_mux);
    
    rx_packet_length_ret_0 : SLE
      port map(D => \un65_sm_advance_i_i[10]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \un65_sm_advance_i[10]\);
    
    \rx_fifo_din_d3[6]\ : SLE
      port map(D => N_21, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_sampler_clk1x_en_inv_0\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN_pipe[6]\);
    
    \consumer_type[9]\ : SLE
      port map(D => \consumer_type_12[9]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_12, ALn
         => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type[9]_net_1\);
    
    \ReadFIFO_WR_SM.un35_sm_advance_i_NE_6\ : CFG4
      generic map(INIT => x"FFF6")

      port map(A => \consumer_type[4]_net_1\, B => 
        consumer_type3_reg(4), C => un35_sm_advance_i_NE_3, D => 
        un35_sm_advance_i_5, Y => un35_sm_advance_i_NE_6);
    
    \ReadFIFO_WR_SM.un1_sampler_clk1x_en_0_I_33\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \rx_crc_data_store[11]_net_1\, B => 
        \rx_crc_data_calc[10]\, C => \rx_crc_data_calc[11]\, D
         => \rx_crc_data_store[10]_net_1\, FCI => 
        \un1_sampler_clk1x_en_0_data_tmp[4]\, S => OPEN, Y => 
        OPEN, FCO => \un1_sampler_clk1x_en_0_data_tmp[5]\);
    
    \rx_crc_data_store[6]\ : SLE
      port map(D => \un1_rx_fifo_din_d3[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_sampler_clk1x_en_inv_i, 
        ALn => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[6]_net_1\);
    
    SM_advance_i : SLE
      port map(D => un2_packet_avail, CLK => CommsFPGA_CCC_0_GL0, 
        EN => N_221, ALn => un9_rst_i, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \SM_advance_i\);
    
    rx_crc_HighByte_en_RNO : CFG2
      generic map(INIT => x"4")

      port map(A => \un58_sm_advance_i_0_data_tmp[5]\, B => 
        \un15[5]\, Y => N_225_i);
    
    \consumer_type[3]\ : SLE
      port map(D => \consumer_type_12[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_12, ALn
         => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type[3]_net_1\);
    
    un1_ReadFIFO_WR_STATE_14_0_o2 : CFG2
      generic map(INIT => x"E")

      port map(A => \un15[5]\, B => \un15[3]\, Y => N_276);
    
    \rx_byte_cntr[3]\ : SLE
      port map(D => \rx_byte_cntr_lm[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => rx_byte_cntre, ALn => RESET_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \rx_byte_cntr[3]_net_1\);
    
    \rx_crc_data_store[3]\ : SLE
      port map(D => \un1_rx_fifo_din_d3[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_sampler_clk1x_en_inv_i, 
        ALn => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[3]_net_1\);
    
    \rx_byte_cntr[7]\ : SLE
      port map(D => \rx_byte_cntr_lm[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => rx_byte_cntre, ALn => RESET_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \rx_byte_cntr[7]_net_1\);
    
    RX_InProcess_d1 : SLE
      port map(D => \RX_InProcess\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => RESET_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RX_InProcess_d1\);
    
    \consumer_type[8]\ : SLE
      port map(D => \consumer_type_12[8]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_12, ALn
         => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type[8]_net_1\);
    
    \rx_packet_length[3]\ : SLE
      port map(D => \rx_packet_length_13[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rx_packet_length[3]_net_1\);
    
    \SM_advancebit_cntr_RNO[1]\ : CFG3
      generic map(INIT => x"6A")

      port map(A => \SM_advancebit_cntr[1]_net_1\, B => 
        \SM_advancebit_cntr[0]_net_1\, C => N_221, Y => N_121);
    
    \rx_packet_length_ret[6]\ : SLE
      port map(D => \un56_sm_advance_i_i[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_14, ALn
         => RESET_i, ADn => GND_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \un56_sm_advance_i[5]\);
    
    irx_packet_end : SLE
      port map(D => N_689_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => rx_packet_end);
    
    rx_crc_gen : SLE
      port map(D => \un1_ReadFIFO_WR_STATE_15\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => 
        \un1_iRX_EarlyTerm_1_sqmuxa_1_0\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_crc_gen\);
    
    \rx_fifo_din_d1[6]\ : SLE
      port map(D => RX_FIFO_DIN(6), CLK => CommsFPGA_CCC_0_GL0, 
        EN => \un1_sampler_clk1x_en_inv_0\, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => N_20);
    
    \rx_packet_length_13[7]\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_652_mux, B => un1_ReadFIFO_WR_STATE_6_i, Y
         => \rx_packet_length_13[7]_net_1\);
    
    \rx_fifo_din_d3[3]\ : SLE
      port map(D => N_12, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_sampler_clk1x_en_inv_0\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN_pipe[3]\);
    
    un56_sm_advance_i_cry_7_0 : ARI1
      generic map(INIT => x"511FF")

      port map(A => N_651_mux, B => \un15[7]\, C => \un15[8]\, D
         => GND_net_1, FCI => un56_sm_advance_i_cry_6, S => 
        \un56_sm_advance_i_i[4]\, Y => OPEN, FCO => 
        un56_sm_advance_i_cry_7);
    
    \rx_fifo_din_d3[0]\ : SLE
      port map(D => N_3, CLK => CommsFPGA_CCC_0_GL0, EN => 
        \un1_sampler_clk1x_en_inv_0\, ALn => RESET_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_DIN_pipe[0]\);
    
    \ReadFIFO_WR_STATE[5]\ : SLE
      port map(D => \ReadFIFO_WR_STATE_ns[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \un15[5]\);
    
    \ReadFIFO_WR_SM.un1_sampler_clk1x_en_0_I_1\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \rx_crc_data_store[1]_net_1\, B => 
        \rx_crc_data_calc[0]\, C => \rx_crc_data_calc[1]\, D => 
        \rx_crc_data_store[0]_net_1\, FCI => GND_net_1, S => OPEN, 
        Y => OPEN, FCO => \un1_sampler_clk1x_en_0_data_tmp[0]\);
    
    un65_sm_advance_i_cry_6_0 : ARI1
      generic map(INIT => x"511FF")

      port map(A => N_652_mux, B => \un15[7]\, C => \un15[8]\, D
         => GND_net_1, FCI => un65_sm_advance_i_cry_5, S => 
        \un65_sm_advance_i_i[5]\, Y => OPEN, FCO => 
        un65_sm_advance_i_cry_6);
    
    un65_sm_advance_i_s_10 : CFG3
      generic map(INIT => x"27")

      port map(A => N_4706_i, B => un65_sm_advance_i_cry_8, C => 
        \un65_sm_advance_i_cry_9_ma\, Y => 
        \un65_sm_advance_i_i[1]\);
    
    un1_ReadFIFO_WR_STATE_14_0_a2 : CFG3
      generic map(INIT => x"51")

      port map(A => \un15[2]\, B => \un15[1]\, C => 
        sampler_clk1x_en, Y => N_321);
    
    \ReadFIFO_WR_SM.un1_sampler_clk1x_en_0_I_27\ : ARI1
      generic map(INIT => x"68421")

      port map(A => \rx_crc_data_store[7]_net_1\, B => 
        \rx_crc_data_calc[6]\, C => \rx_crc_data_calc[7]\, D => 
        \rx_crc_data_store[6]_net_1\, FCI => 
        \un1_sampler_clk1x_en_0_data_tmp[2]\, S => OPEN, Y => 
        OPEN, FCO => \un1_sampler_clk1x_en_0_data_tmp[3]\);
    
    \consumer_type[2]\ : SLE
      port map(D => \consumer_type_12[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => un1_ReadFIFO_WR_STATE_12, ALn
         => RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type[2]_net_1\);
    
    \rx_crc_data_store[15]\ : SLE
      port map(D => \RX_FIFO_DIN_pipe[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => rx_crc_data_store_151, ALn => 
        RESET_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \rx_crc_data_store[15]_net_1\);
    
    rx_CRC_error_RNIASV4 : CFG1
      generic map(INIT => "01")

      port map(A => rx_CRC_error_net_1, Y => rx_CRC_error_i);
    
    \ReadFIFO_WR_SM.un32_sm_advance_i_NE_3\ : CFG4
      generic map(INIT => x"7BDE")

      port map(A => consumer_type2_reg(7), B => 
        consumer_type2_reg(6), C => \consumer_type[7]_net_1\, D
         => \consumer_type[6]_net_1\, Y => un32_sm_advance_i_NE_3);
    
    \CoreAPB3_0_APBmslave0_PRDATA_m[4]\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        CoreAPB3_0_APBmslave0_PRDATA(4), Y => 
        CoreAPB3_0_APBmslave0_PRDATA_m(4));
    
    \rx_byte_cntr_lm_0[8]\ : CFG2
      generic map(INIT => x"4")

      port map(A => un1_iRX_EarlyTerm_0_sqmuxa, B => 
        \rx_byte_cntr_s[8]\, Y => \rx_byte_cntr_lm[8]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity AFE_RX_SM is

    port( RX_FIFO_DIN         : in    std_logic_vector(7 downto 0);
          manches_in_dly      : in    std_logic_vector(1 downto 0);
          un6                 : out   std_logic_vector(5 downto 0);
          irx_center_sample   : in    std_logic;
          idle_line           : in    std_logic;
          RX_EarlyTerm        : in    std_logic;
          RESET               : in    std_logic;
          clk1x_enable        : out   std_logic;
          packet_avail        : out   std_logic;
          RESET_i             : in    std_logic;
          rx_packet_end_all   : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic
        );

end AFE_RX_SM;

architecture DEF_ARCH of AFE_RX_SM is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \RX_EarlyTerm_s\, VCC_net_1, \RX_EarlyTerm_s_0\, 
        GND_net_1, \rx_packet_end_all\, irx_packet_end_all_5, 
        packet_avail_6, clk1x_enable_1, \start_bit_mask\, 
        start_bit_cntre, \start_bit_maskce\, \un6[5]\, N_88_i, 
        \un6[4]\, \AFE_RX_STATE_ns[1]\, \un6[3]\, 
        \AFE_RX_STATE_ns[2]_net_1\, \un6[2]\, 
        \AFE_RX_STATE_ns[3]_net_1\, \un6[0]\, 
        \AFE_RX_STATE_ns[4]_net_1\, \start_bit_cntr[0]_net_1\, 
        \start_bit_cntr_s[0]\, \start_bit_cntr[1]_net_1\, 
        \start_bit_cntr_s[1]\, \start_bit_cntr[2]_net_1\, 
        \start_bit_cntr_s[2]\, \start_bit_cntr[3]_net_1\, 
        \start_bit_cntr_s[3]\, \start_bit_cntr[4]_net_1\, 
        \start_bit_cntr_s[4]\, \start_bit_cntr[5]_net_1\, 
        \start_bit_cntr_s[5]\, \start_bit_cntr[6]_net_1\, 
        \start_bit_cntr_s[6]\, \start_bit_cntr[7]_net_1\, 
        \start_bit_cntr_s[7]_net_1\, start_bit_cntr_cry_cy, 
        un5_reset, \start_bit_cntr_cry[0]_net_1\, 
        \start_bit_cntr_cry[1]_net_1\, 
        \start_bit_cntr_cry[2]_net_1\, 
        \start_bit_cntr_cry[3]_net_1\, 
        \start_bit_cntr_cry[4]_net_1\, 
        \start_bit_cntr_cry[5]_net_1\, 
        \start_bit_cntr_cry[6]_net_1\, un1_rx_fifo_din_5, 
        un1_rx_fifo_din_4, un2_sample_5, un2_sample_4, 
        un1_rx_fifo_din, N_93 : std_logic;

begin 

    un6(5) <= \un6[5]\;
    un6(4) <= \un6[4]\;
    un6(3) <= \un6[3]\;
    un6(2) <= \un6[2]\;
    un6(0) <= \un6[0]\;
    rx_packet_end_all <= \rx_packet_end_all\;

    \start_bit_cntr[2]\ : SLE
      port map(D => \start_bit_cntr_s[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => start_bit_cntre, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \start_bit_cntr[2]_net_1\);
    
    RX_EarlyTerm_s_0 : CFG2
      generic map(INIT => x"4")

      port map(A => RESET, B => RX_EarlyTerm, Y => 
        \RX_EarlyTerm_s_0\);
    
    \AFE_RX_STATE[3]\ : SLE
      port map(D => \AFE_RX_STATE_ns[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \un6[4]\);
    
    \AFE_RX_SM.irx_packet_end_all_5_0_a3\ : CFG3
      generic map(INIT => x"04")

      port map(A => \un6[5]\, B => idle_line, C => \un6[2]\, Y
         => irx_packet_end_all_5);
    
    \AFE_RX_STATE_ns[2]\ : CFG4
      generic map(INIT => x"0A0E")

      port map(A => \un6[4]\, B => \un6[3]\, C => idle_line, D
         => un1_rx_fifo_din, Y => \AFE_RX_STATE_ns[2]_net_1\);
    
    \start_bit_cntr[5]\ : SLE
      port map(D => \start_bit_cntr_s[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => start_bit_cntre, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \start_bit_cntr[5]_net_1\);
    
    \AFE_RX_SM.un1_rx_fifo_din_4\ : CFG3
      generic map(INIT => x"02")

      port map(A => RX_FIFO_DIN(2), B => \start_bit_mask\, C => 
        RX_FIFO_DIN(3), Y => un1_rx_fifo_din_4);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \start_bit_cntr_cry_cy[0]\ : ARI1
      generic map(INIT => x"45500")

      port map(A => VCC_net_1, B => un5_reset, C => GND_net_1, D
         => GND_net_1, FCI => VCC_net_1, S => OPEN, Y => OPEN, 
        FCO => start_bit_cntr_cry_cy);
    
    start_bit_maskce : CFG2
      generic map(INIT => x"E")

      port map(A => un5_reset, B => irx_center_sample, Y => 
        \start_bit_maskce\);
    
    \start_bit_cntr[3]\ : SLE
      port map(D => \start_bit_cntr_s[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => start_bit_cntre, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \start_bit_cntr[3]_net_1\);
    
    \start_bit_cntr_cry[5]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => un5_reset, C => 
        \start_bit_cntr[5]_net_1\, D => GND_net_1, FCI => 
        \start_bit_cntr_cry[4]_net_1\, S => \start_bit_cntr_s[5]\, 
        Y => OPEN, FCO => \start_bit_cntr_cry[5]_net_1\);
    
    \AFE_RX_STATE_ns_a3[3]\ : CFG3
      generic map(INIT => x"20")

      port map(A => \un6[3]\, B => idle_line, C => 
        un1_rx_fifo_din, Y => N_93);
    
    \AFE_RX_STATE_ns_a3[1]\ : CFG3
      generic map(INIT => x"40")

      port map(A => manches_in_dly(1), B => manches_in_dly(0), C
         => \un6[5]\, Y => \AFE_RX_STATE_ns[1]\);
    
    \start_bit_cntr_cry[0]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => un5_reset, C => 
        \start_bit_cntr[0]_net_1\, D => GND_net_1, FCI => 
        start_bit_cntr_cry_cy, S => \start_bit_cntr_s[0]\, Y => 
        OPEN, FCO => \start_bit_cntr_cry[0]_net_1\);
    
    \AFE_RX_STATE[1]\ : SLE
      port map(D => \AFE_RX_STATE_ns[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \un6[2]\);
    
    clk1x_enable_1_0 : CFG4
      generic map(INIT => x"3337")

      port map(A => \un6[5]\, B => N_88_i, C => \un6[4]\, D => 
        \un6[3]\, Y => clk1x_enable_1);
    
    \AFE_RX_STATE[4]\ : SLE
      port map(D => N_88_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => RESET_i, ADn => GND_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \un6[5]\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \start_bit_cntr[0]\ : SLE
      port map(D => \start_bit_cntr_s[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => start_bit_cntre, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \start_bit_cntr[0]_net_1\);
    
    RX_EarlyTerm_s : SLE
      port map(D => \RX_EarlyTerm_s_0\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => VCC_net_1, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RX_EarlyTerm_s\);
    
    \start_bit_cntr[1]\ : SLE
      port map(D => \start_bit_cntr_s[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => start_bit_cntre, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \start_bit_cntr[1]_net_1\);
    
    \AFE_RX_STATE[0]\ : SLE
      port map(D => \AFE_RX_STATE_ns[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \un6[0]\);
    
    \START_BIT_COUNTER_PROC.un2_sample_4_RNIC6DG1\ : CFG4
      generic map(INIT => x"FF2A")

      port map(A => irx_center_sample, B => un2_sample_5, C => 
        un2_sample_4, D => un5_reset, Y => start_bit_cntre);
    
    \start_bit_cntr[4]\ : SLE
      port map(D => \start_bit_cntr_s[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => start_bit_cntre, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \start_bit_cntr[4]_net_1\);
    
    \start_bit_cntr_s[7]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => un5_reset, C => 
        \start_bit_cntr[7]_net_1\, D => GND_net_1, FCI => 
        \start_bit_cntr_cry[6]_net_1\, S => 
        \start_bit_cntr_s[7]_net_1\, Y => OPEN, FCO => OPEN);
    
    \AFE_RX_SM.un1_rx_fifo_din\ : CFG4
      generic map(INIT => x"4000")

      port map(A => RX_FIFO_DIN(1), B => RX_FIFO_DIN(6), C => 
        un1_rx_fifo_din_5, D => un1_rx_fifo_din_4, Y => 
        un1_rx_fifo_din);
    
    packet_avail_6_0 : CFG4
      generic map(INIT => x"FAF2")

      port map(A => \un6[2]\, B => \RX_EarlyTerm_s\, C => N_93, D
         => idle_line, Y => packet_avail_6);
    
    \AFE_RX_SM.un1_rx_fifo_din_5\ : CFG4
      generic map(INIT => x"2000")

      port map(A => RX_FIFO_DIN(7), B => RX_FIFO_DIN(5), C => 
        RX_FIFO_DIN(4), D => RX_FIFO_DIN(0), Y => 
        un1_rx_fifo_din_5);
    
    \START_BIT_COUNTER_PROC.un2_sample_5\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \start_bit_cntr[4]_net_1\, B => 
        \start_bit_cntr[3]_net_1\, C => \start_bit_cntr[1]_net_1\, 
        D => \start_bit_cntr[0]_net_1\, Y => un2_sample_5);
    
    \start_bit_cntr_cry[6]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => un5_reset, C => 
        \start_bit_cntr[6]_net_1\, D => GND_net_1, FCI => 
        \start_bit_cntr_cry[5]_net_1\, S => \start_bit_cntr_s[6]\, 
        Y => OPEN, FCO => \start_bit_cntr_cry[6]_net_1\);
    
    \AFE_RX_STATE_ns[3]\ : CFG4
      generic map(INIT => x"F0F2")

      port map(A => \un6[2]\, B => \RX_EarlyTerm_s\, C => N_93, D
         => idle_line, Y => \AFE_RX_STATE_ns[3]_net_1\);
    
    \AFE_RX_STATE_ns[4]\ : CFG4
      generic map(INIT => x"0E0A")

      port map(A => \un6[0]\, B => \RX_EarlyTerm_s\, C => 
        idle_line, D => \un6[2]\, Y => \AFE_RX_STATE_ns[4]_net_1\);
    
    \start_bit_cntr[6]\ : SLE
      port map(D => \start_bit_cntr_s[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => start_bit_cntre, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \start_bit_cntr[6]_net_1\);
    
    \AFE_RX_STATE_ns_i_o3[0]\ : CFG3
      generic map(INIT => x"0E")

      port map(A => \un6[5]\, B => idle_line, C => 
        \AFE_RX_STATE_ns[1]\, Y => N_88_i);
    
    \packet_avail\ : SLE
      port map(D => packet_avail_6, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => RESET_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        packet_avail);
    
    irx_packet_end_all : SLE
      port map(D => irx_packet_end_all_5, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_packet_end_all\);
    
    \start_bit_cntr_cry[3]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => un5_reset, C => 
        \start_bit_cntr[3]_net_1\, D => GND_net_1, FCI => 
        \start_bit_cntr_cry[2]_net_1\, S => \start_bit_cntr_s[3]\, 
        Y => OPEN, FCO => \start_bit_cntr_cry[3]_net_1\);
    
    \AFE_RX_STATE[2]\ : SLE
      port map(D => \AFE_RX_STATE_ns[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \un6[3]\);
    
    \start_bit_cntr_cry[2]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => un5_reset, C => 
        \start_bit_cntr[2]_net_1\, D => GND_net_1, FCI => 
        \start_bit_cntr_cry[1]_net_1\, S => \start_bit_cntr_s[2]\, 
        Y => OPEN, FCO => \start_bit_cntr_cry[2]_net_1\);
    
    \start_bit_cntr[7]\ : SLE
      port map(D => \start_bit_cntr_s[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => start_bit_cntre, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        \start_bit_cntr[7]_net_1\);
    
    start_bit_mask : SLE
      port map(D => start_bit_cntre, CLK => CommsFPGA_CCC_0_GL0, 
        EN => \start_bit_maskce\, ALn => VCC_net_1, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \start_bit_mask\);
    
    \start_bit_cntr_cry[4]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => un5_reset, C => 
        \start_bit_cntr[4]_net_1\, D => GND_net_1, FCI => 
        \start_bit_cntr_cry[3]_net_1\, S => \start_bit_cntr_s[4]\, 
        Y => OPEN, FCO => \start_bit_cntr_cry[4]_net_1\);
    
    \start_bit_cntr_cry[1]\ : ARI1
      generic map(INIT => x"44400")

      port map(A => VCC_net_1, B => un5_reset, C => 
        \start_bit_cntr[1]_net_1\, D => GND_net_1, FCI => 
        \start_bit_cntr_cry[0]_net_1\, S => \start_bit_cntr_s[1]\, 
        Y => OPEN, FCO => \start_bit_cntr_cry[1]_net_1\);
    
    \START_BIT_COUNTER_PROC.un5_reset\ : CFG3
      generic map(INIT => x"FE")

      port map(A => RESET, B => \rx_packet_end_all\, C => 
        \un6[5]\, Y => un5_reset);
    
    \clk1x_enable\ : SLE
      port map(D => clk1x_enable_1, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => RESET_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        clk1x_enable);
    
    \START_BIT_COUNTER_PROC.un2_sample_4\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \start_bit_cntr[7]_net_1\, B => 
        \start_bit_cntr[6]_net_1\, C => \start_bit_cntr[5]_net_1\, 
        D => \start_bit_cntr[2]_net_1\, Y => un2_sample_4);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity ManchesDecoder is

    port( un6                                : out   std_logic_vector(5 downto 0);
          manches_in_dly                     : out   std_logic_vector(1 downto 0);
          clkdiv                             : out   std_logic_vector(3 downto 0);
          RX_FIFO_DIN_pipe                   : out   std_logic_vector(8 downto 0);
          RX_FIFO_DIN                        : out   std_logic_vector(7 downto 0);
          un15                               : out   std_logic_vector(10 downto 0);
          CoreAPB3_0_APBmslave0_PRDATA       : in    std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PRDATA_m     : out   std_logic_vector(7 downto 0);
          consumer_type2_reg                 : in    std_logic_vector(9 downto 0);
          consumer_type1_reg                 : in    std_logic_vector(9 downto 0);
          consumer_type3_reg                 : in    std_logic_vector(9 downto 0);
          consumer_type4_reg                 : in    std_logic_vector(9 downto 0);
          iNRZ_data                          : out   std_logic;
          irx_center_sample                  : out   std_logic;
          internal_loopback                  : in    std_logic;
          MANCH_OUT_P_c                      : in    std_logic;
          MANCHESTER_IN_c                    : in    std_logic;
          idle_line5                         : in    std_logic;
          rx_CRC_error                       : out   std_logic;
          rx_CRC_error_i                     : out   std_logic;
          CommsFPGA_CCC_0_GL0                : in    std_logic;
          RESET_i                            : in    std_logic;
          RX_EarlyTerm                       : out   std_logic;
          rx_packet_complt                   : out   std_logic;
          CoreAPB3_0_APBmslave0_PSELx        : in    std_logic;
          tx_col_detect_en                   : in    std_logic;
          RX_FIFO_TxColDetDis_wr_en          : out   std_logic;
          RESET                              : in    std_logic;
          CoreAPB3_0_APBmslave0_PREADY       : in    std_logic;
          CoreAPB3_0_APBmslave0_PREADY_i_m_i : out   std_logic;
          DRVR_EN_c                          : in    std_logic
        );

end ManchesDecoder;

architecture DEF_ARCH of ManchesDecoder is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component ManchesDecoder_Adapter
    port( clkdiv              : out   std_logic_vector(3 downto 0);
          RX_FIFO_DIN         : out   std_logic_vector(7 downto 0);
          manches_in_dly      : out   std_logic_vector(1 downto 0);
          idle_line5          : in    std_logic := 'U';
          RESET               : in    std_logic := 'U';
          MANCHESTER_IN_c     : in    std_logic := 'U';
          MANCH_OUT_P_c       : in    std_logic := 'U';
          internal_loopback   : in    std_logic := 'U';
          rx_packet_end_all   : in    std_logic := 'U';
          idle_line           : out   std_logic;
          irx_center_sample   : out   std_logic;
          sampler_clk1x_en    : out   std_logic;
          iNRZ_data           : out   std_logic;
          clk1x_enable        : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          RESET_i             : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component ReadFIFO_Write_SM
    port( consumer_type4_reg                 : in    std_logic_vector(9 downto 0) := (others => 'U');
          consumer_type3_reg                 : in    std_logic_vector(9 downto 0) := (others => 'U');
          consumer_type1_reg                 : in    std_logic_vector(9 downto 0) := (others => 'U');
          consumer_type2_reg                 : in    std_logic_vector(9 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PRDATA_m     : out   std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PRDATA       : in    std_logic_vector(7 downto 0) := (others => 'U');
          un15                               : out   std_logic_vector(10 downto 0);
          RX_FIFO_DIN                        : in    std_logic_vector(7 downto 0) := (others => 'U');
          RX_FIFO_DIN_pipe                   : out   std_logic_vector(8 downto 0);
          DRVR_EN_c                          : in    std_logic := 'U';
          clk1x_enable                       : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PREADY_i_m_i : out   std_logic;
          CoreAPB3_0_APBmslave0_PREADY       : in    std_logic := 'U';
          RESET                              : in    std_logic := 'U';
          RX_FIFO_TxColDetDis_wr_en          : out   std_logic;
          tx_col_detect_en                   : in    std_logic := 'U';
          idle_line                          : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PSELx        : in    std_logic := 'U';
          sampler_clk1x_en                   : in    std_logic := 'U';
          packet_avail                       : in    std_logic := 'U';
          rx_packet_complt                   : out   std_logic;
          RX_EarlyTerm                       : out   std_logic;
          RESET_i                            : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0                : in    std_logic := 'U';
          rx_CRC_error_i                     : out   std_logic;
          rx_CRC_error                       : out   std_logic
        );
  end component;

  component AFE_RX_SM
    port( RX_FIFO_DIN         : in    std_logic_vector(7 downto 0) := (others => 'U');
          manches_in_dly      : in    std_logic_vector(1 downto 0) := (others => 'U');
          un6                 : out   std_logic_vector(5 downto 0);
          irx_center_sample   : in    std_logic := 'U';
          idle_line           : in    std_logic := 'U';
          RX_EarlyTerm        : in    std_logic := 'U';
          RESET               : in    std_logic := 'U';
          clk1x_enable        : out   std_logic;
          packet_avail        : out   std_logic;
          RESET_i             : in    std_logic := 'U';
          rx_packet_end_all   : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U'
        );
  end component;

    signal \RX_FIFO_DIN[0]\, \RX_FIFO_DIN[1]\, \RX_FIFO_DIN[2]\, 
        \RX_FIFO_DIN[3]\, \RX_FIFO_DIN[4]\, \RX_FIFO_DIN[5]\, 
        \RX_FIFO_DIN[6]\, \RX_FIFO_DIN[7]\, clk1x_enable, 
        idle_line, sampler_clk1x_en, packet_avail, \RX_EarlyTerm\, 
        \manches_in_dly[0]\, \manches_in_dly[1]\, 
        rx_packet_end_all, \irx_center_sample\, GND_net_1, 
        VCC_net_1 : std_logic;
    signal nc2, nc1 : std_logic;

    for all : ManchesDecoder_Adapter
	Use entity work.ManchesDecoder_Adapter(DEF_ARCH);
    for all : ReadFIFO_Write_SM
	Use entity work.ReadFIFO_Write_SM(DEF_ARCH);
    for all : AFE_RX_SM
	Use entity work.AFE_RX_SM(DEF_ARCH);
begin 

    manches_in_dly(1) <= \manches_in_dly[1]\;
    manches_in_dly(0) <= \manches_in_dly[0]\;
    RX_FIFO_DIN(7) <= \RX_FIFO_DIN[7]\;
    RX_FIFO_DIN(6) <= \RX_FIFO_DIN[6]\;
    RX_FIFO_DIN(5) <= \RX_FIFO_DIN[5]\;
    RX_FIFO_DIN(4) <= \RX_FIFO_DIN[4]\;
    RX_FIFO_DIN(3) <= \RX_FIFO_DIN[3]\;
    RX_FIFO_DIN(2) <= \RX_FIFO_DIN[2]\;
    RX_FIFO_DIN(1) <= \RX_FIFO_DIN[1]\;
    RX_FIFO_DIN(0) <= \RX_FIFO_DIN[0]\;
    irx_center_sample <= \irx_center_sample\;
    RX_EarlyTerm <= \RX_EarlyTerm\;

    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    MANCHESTER_DECODER_ADAPTER_INST : ManchesDecoder_Adapter
      port map(clkdiv(3) => clkdiv(3), clkdiv(2) => clkdiv(2), 
        clkdiv(1) => clkdiv(1), clkdiv(0) => clkdiv(0), 
        RX_FIFO_DIN(7) => \RX_FIFO_DIN[7]\, RX_FIFO_DIN(6) => 
        \RX_FIFO_DIN[6]\, RX_FIFO_DIN(5) => \RX_FIFO_DIN[5]\, 
        RX_FIFO_DIN(4) => \RX_FIFO_DIN[4]\, RX_FIFO_DIN(3) => 
        \RX_FIFO_DIN[3]\, RX_FIFO_DIN(2) => \RX_FIFO_DIN[2]\, 
        RX_FIFO_DIN(1) => \RX_FIFO_DIN[1]\, RX_FIFO_DIN(0) => 
        \RX_FIFO_DIN[0]\, manches_in_dly(1) => 
        \manches_in_dly[1]\, manches_in_dly(0) => 
        \manches_in_dly[0]\, idle_line5 => idle_line5, RESET => 
        RESET, MANCHESTER_IN_c => MANCHESTER_IN_c, MANCH_OUT_P_c
         => MANCH_OUT_P_c, internal_loopback => internal_loopback, 
        rx_packet_end_all => rx_packet_end_all, idle_line => 
        idle_line, irx_center_sample => \irx_center_sample\, 
        sampler_clk1x_en => sampler_clk1x_en, iNRZ_data => 
        iNRZ_data, clk1x_enable => clk1x_enable, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, RESET_i => 
        RESET_i);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    ReadFIFO_Write_SM_PROC : ReadFIFO_Write_SM
      port map(consumer_type4_reg(9) => consumer_type4_reg(9), 
        consumer_type4_reg(8) => consumer_type4_reg(8), 
        consumer_type4_reg(7) => consumer_type4_reg(7), 
        consumer_type4_reg(6) => consumer_type4_reg(6), 
        consumer_type4_reg(5) => consumer_type4_reg(5), 
        consumer_type4_reg(4) => consumer_type4_reg(4), 
        consumer_type4_reg(3) => consumer_type4_reg(3), 
        consumer_type4_reg(2) => consumer_type4_reg(2), 
        consumer_type4_reg(1) => consumer_type4_reg(1), 
        consumer_type4_reg(0) => consumer_type4_reg(0), 
        consumer_type3_reg(9) => consumer_type3_reg(9), 
        consumer_type3_reg(8) => consumer_type3_reg(8), 
        consumer_type3_reg(7) => consumer_type3_reg(7), 
        consumer_type3_reg(6) => consumer_type3_reg(6), 
        consumer_type3_reg(5) => consumer_type3_reg(5), 
        consumer_type3_reg(4) => consumer_type3_reg(4), 
        consumer_type3_reg(3) => consumer_type3_reg(3), 
        consumer_type3_reg(2) => consumer_type3_reg(2), 
        consumer_type3_reg(1) => consumer_type3_reg(1), 
        consumer_type3_reg(0) => consumer_type3_reg(0), 
        consumer_type1_reg(9) => consumer_type1_reg(9), 
        consumer_type1_reg(8) => consumer_type1_reg(8), 
        consumer_type1_reg(7) => consumer_type1_reg(7), 
        consumer_type1_reg(6) => consumer_type1_reg(6), 
        consumer_type1_reg(5) => consumer_type1_reg(5), 
        consumer_type1_reg(4) => consumer_type1_reg(4), 
        consumer_type1_reg(3) => consumer_type1_reg(3), 
        consumer_type1_reg(2) => consumer_type1_reg(2), 
        consumer_type1_reg(1) => consumer_type1_reg(1), 
        consumer_type1_reg(0) => consumer_type1_reg(0), 
        consumer_type2_reg(9) => consumer_type2_reg(9), 
        consumer_type2_reg(8) => consumer_type2_reg(8), 
        consumer_type2_reg(7) => consumer_type2_reg(7), 
        consumer_type2_reg(6) => consumer_type2_reg(6), 
        consumer_type2_reg(5) => consumer_type2_reg(5), 
        consumer_type2_reg(4) => consumer_type2_reg(4), 
        consumer_type2_reg(3) => consumer_type2_reg(3), 
        consumer_type2_reg(2) => consumer_type2_reg(2), 
        consumer_type2_reg(1) => consumer_type2_reg(1), 
        consumer_type2_reg(0) => consumer_type2_reg(0), 
        CoreAPB3_0_APBmslave0_PRDATA_m(7) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(7), 
        CoreAPB3_0_APBmslave0_PRDATA_m(6) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(6), 
        CoreAPB3_0_APBmslave0_PRDATA_m(5) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(5), 
        CoreAPB3_0_APBmslave0_PRDATA_m(4) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(4), 
        CoreAPB3_0_APBmslave0_PRDATA_m(3) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(3), 
        CoreAPB3_0_APBmslave0_PRDATA_m(2) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(2), 
        CoreAPB3_0_APBmslave0_PRDATA_m(1) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(1), 
        CoreAPB3_0_APBmslave0_PRDATA_m(0) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(0), 
        CoreAPB3_0_APBmslave0_PRDATA(7) => 
        CoreAPB3_0_APBmslave0_PRDATA(7), 
        CoreAPB3_0_APBmslave0_PRDATA(6) => 
        CoreAPB3_0_APBmslave0_PRDATA(6), 
        CoreAPB3_0_APBmslave0_PRDATA(5) => 
        CoreAPB3_0_APBmslave0_PRDATA(5), 
        CoreAPB3_0_APBmslave0_PRDATA(4) => 
        CoreAPB3_0_APBmslave0_PRDATA(4), 
        CoreAPB3_0_APBmslave0_PRDATA(3) => 
        CoreAPB3_0_APBmslave0_PRDATA(3), 
        CoreAPB3_0_APBmslave0_PRDATA(2) => 
        CoreAPB3_0_APBmslave0_PRDATA(2), 
        CoreAPB3_0_APBmslave0_PRDATA(1) => 
        CoreAPB3_0_APBmslave0_PRDATA(1), 
        CoreAPB3_0_APBmslave0_PRDATA(0) => 
        CoreAPB3_0_APBmslave0_PRDATA(0), un15(10) => un15(10), 
        un15(9) => un15(9), un15(8) => un15(8), un15(7) => 
        un15(7), un15(6) => nc2, un15(5) => un15(5), un15(4) => 
        un15(4), un15(3) => un15(3), un15(2) => un15(2), un15(1)
         => un15(1), un15(0) => un15(0), RX_FIFO_DIN(7) => 
        \RX_FIFO_DIN[7]\, RX_FIFO_DIN(6) => \RX_FIFO_DIN[6]\, 
        RX_FIFO_DIN(5) => \RX_FIFO_DIN[5]\, RX_FIFO_DIN(4) => 
        \RX_FIFO_DIN[4]\, RX_FIFO_DIN(3) => \RX_FIFO_DIN[3]\, 
        RX_FIFO_DIN(2) => \RX_FIFO_DIN[2]\, RX_FIFO_DIN(1) => 
        \RX_FIFO_DIN[1]\, RX_FIFO_DIN(0) => \RX_FIFO_DIN[0]\, 
        RX_FIFO_DIN_pipe(8) => RX_FIFO_DIN_pipe(8), 
        RX_FIFO_DIN_pipe(7) => RX_FIFO_DIN_pipe(7), 
        RX_FIFO_DIN_pipe(6) => RX_FIFO_DIN_pipe(6), 
        RX_FIFO_DIN_pipe(5) => RX_FIFO_DIN_pipe(5), 
        RX_FIFO_DIN_pipe(4) => RX_FIFO_DIN_pipe(4), 
        RX_FIFO_DIN_pipe(3) => RX_FIFO_DIN_pipe(3), 
        RX_FIFO_DIN_pipe(2) => RX_FIFO_DIN_pipe(2), 
        RX_FIFO_DIN_pipe(1) => RX_FIFO_DIN_pipe(1), 
        RX_FIFO_DIN_pipe(0) => RX_FIFO_DIN_pipe(0), DRVR_EN_c => 
        DRVR_EN_c, clk1x_enable => clk1x_enable, 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i => 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i, 
        CoreAPB3_0_APBmslave0_PREADY => 
        CoreAPB3_0_APBmslave0_PREADY, RESET => RESET, 
        RX_FIFO_TxColDetDis_wr_en => RX_FIFO_TxColDetDis_wr_en, 
        tx_col_detect_en => tx_col_detect_en, idle_line => 
        idle_line, CoreAPB3_0_APBmslave0_PSELx => 
        CoreAPB3_0_APBmslave0_PSELx, sampler_clk1x_en => 
        sampler_clk1x_en, packet_avail => packet_avail, 
        rx_packet_complt => rx_packet_complt, RX_EarlyTerm => 
        \RX_EarlyTerm\, RESET_i => RESET_i, CommsFPGA_CCC_0_GL0
         => CommsFPGA_CCC_0_GL0, rx_CRC_error_i => rx_CRC_error_i, 
        rx_CRC_error => rx_CRC_error);
    
    AFE_RX_STATE_MACHINE : AFE_RX_SM
      port map(RX_FIFO_DIN(7) => \RX_FIFO_DIN[7]\, RX_FIFO_DIN(6)
         => \RX_FIFO_DIN[6]\, RX_FIFO_DIN(5) => \RX_FIFO_DIN[5]\, 
        RX_FIFO_DIN(4) => \RX_FIFO_DIN[4]\, RX_FIFO_DIN(3) => 
        \RX_FIFO_DIN[3]\, RX_FIFO_DIN(2) => \RX_FIFO_DIN[2]\, 
        RX_FIFO_DIN(1) => \RX_FIFO_DIN[1]\, RX_FIFO_DIN(0) => 
        \RX_FIFO_DIN[0]\, manches_in_dly(1) => 
        \manches_in_dly[1]\, manches_in_dly(0) => 
        \manches_in_dly[0]\, un6(5) => un6(5), un6(4) => un6(4), 
        un6(3) => un6(3), un6(2) => un6(2), un6(1) => nc1, un6(0)
         => un6(0), irx_center_sample => \irx_center_sample\, 
        idle_line => idle_line, RX_EarlyTerm => \RX_EarlyTerm\, 
        RESET => RESET, clk1x_enable => clk1x_enable, 
        packet_avail => packet_avail, RESET_i => RESET_i, 
        rx_packet_end_all => rx_packet_end_all, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_2Kx8_FIFO_2Kx8_0_LSRAM_top is

    port( fifo_MEMWADDR                : in    std_logic_vector(10 downto 0);
          CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0);
          fifo_MEMRADDR                : in    std_logic_vector(10 downto 0);
          RDATA_int                    : out   std_logic_vector(7 downto 0);
          fifo_MEMWE                   : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic;
          N_19_i                       : in    std_logic;
          BIT_CLK                      : in    std_logic
        );

end FIFO_2Kx8_FIFO_2Kx8_0_LSRAM_top;

architecture DEF_ARCH of FIFO_2Kx8_FIFO_2Kx8_0_LSRAM_top is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component RAM1K18
    generic (MEMORYFILE:string := "");

    port( A_DOUT        : out   std_logic_vector(17 downto 0);
          B_DOUT        : out   std_logic_vector(17 downto 0);
          BUSY          : out   std_logic;
          A_CLK         : in    std_logic := 'U';
          A_DOUT_CLK    : in    std_logic := 'U';
          A_ARST_N      : in    std_logic := 'U';
          A_DOUT_EN     : in    std_logic := 'U';
          A_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_DOUT_ARST_N : in    std_logic := 'U';
          A_DOUT_SRST_N : in    std_logic := 'U';
          A_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          A_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          A_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          B_CLK         : in    std_logic := 'U';
          B_DOUT_CLK    : in    std_logic := 'U';
          B_ARST_N      : in    std_logic := 'U';
          B_DOUT_EN     : in    std_logic := 'U';
          B_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_DOUT_ARST_N : in    std_logic := 'U';
          B_DOUT_SRST_N : in    std_logic := 'U';
          B_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          B_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          B_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          A_EN          : in    std_logic := 'U';
          A_DOUT_LAT    : in    std_logic := 'U';
          A_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_WMODE       : in    std_logic := 'U';
          B_EN          : in    std_logic := 'U';
          B_DOUT_LAT    : in    std_logic := 'U';
          B_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_WMODE       : in    std_logic := 'U';
          SII_LOCK      : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;
    signal nc24, nc1, nc8, nc13, nc16, nc19, nc25, nc20, nc27, 
        nc9, nc22, nc28, nc14, nc5, nc21, nc15, nc3, nc10, nc7, 
        nc17, nc4, nc12, nc2, nc23, nc18, nc26, nc6, nc11
         : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    FIFO_2Kx8_FIFO_2Kx8_0_LSRAM_top_R0C0 : RAM1K18
      port map(A_DOUT(17) => nc24, A_DOUT(16) => nc1, A_DOUT(15)
         => nc8, A_DOUT(14) => nc13, A_DOUT(13) => nc16, 
        A_DOUT(12) => nc19, A_DOUT(11) => nc25, A_DOUT(10) => 
        nc20, A_DOUT(9) => nc27, A_DOUT(8) => nc9, A_DOUT(7) => 
        RDATA_int(7), A_DOUT(6) => RDATA_int(6), A_DOUT(5) => 
        RDATA_int(5), A_DOUT(4) => RDATA_int(4), A_DOUT(3) => 
        RDATA_int(3), A_DOUT(2) => RDATA_int(2), A_DOUT(1) => 
        RDATA_int(1), A_DOUT(0) => RDATA_int(0), B_DOUT(17) => 
        nc22, B_DOUT(16) => nc28, B_DOUT(15) => nc14, B_DOUT(14)
         => nc5, B_DOUT(13) => nc21, B_DOUT(12) => nc15, 
        B_DOUT(11) => nc3, B_DOUT(10) => nc10, B_DOUT(9) => nc7, 
        B_DOUT(8) => nc17, B_DOUT(7) => nc4, B_DOUT(6) => nc12, 
        B_DOUT(5) => nc2, B_DOUT(4) => nc23, B_DOUT(3) => nc18, 
        B_DOUT(2) => nc26, B_DOUT(1) => nc6, B_DOUT(0) => nc11, 
        BUSY => OPEN, A_CLK => BIT_CLK, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => N_19_i, A_BLK(1) => VCC_net_1, A_BLK(0) => VCC_net_1, 
        A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => VCC_net_1, 
        A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, A_DIN(15)
         => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13) => 
        GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => GND_net_1, 
        A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, A_DIN(8)
         => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6) => 
        GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => GND_net_1, 
        A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, A_DIN(1)
         => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13) => 
        fifo_MEMRADDR(10), A_ADDR(12) => fifo_MEMRADDR(9), 
        A_ADDR(11) => fifo_MEMRADDR(8), A_ADDR(10) => 
        fifo_MEMRADDR(7), A_ADDR(9) => fifo_MEMRADDR(6), 
        A_ADDR(8) => fifo_MEMRADDR(5), A_ADDR(7) => 
        fifo_MEMRADDR(4), A_ADDR(6) => fifo_MEMRADDR(3), 
        A_ADDR(5) => fifo_MEMRADDR(2), A_ADDR(4) => 
        fifo_MEMRADDR(1), A_ADDR(3) => fifo_MEMRADDR(0), 
        A_ADDR(2) => GND_net_1, A_ADDR(1) => GND_net_1, A_ADDR(0)
         => GND_net_1, A_WEN(1) => GND_net_1, A_WEN(0) => 
        GND_net_1, B_CLK => m2s010_som_sb_0_CCC_71MHz, B_DOUT_CLK
         => VCC_net_1, B_ARST_N => VCC_net_1, B_DOUT_EN => 
        VCC_net_1, B_BLK(2) => fifo_MEMWE, B_BLK(1) => VCC_net_1, 
        B_BLK(0) => VCC_net_1, B_DOUT_ARST_N => GND_net_1, 
        B_DOUT_SRST_N => VCC_net_1, B_DIN(17) => GND_net_1, 
        B_DIN(16) => GND_net_1, B_DIN(15) => GND_net_1, B_DIN(14)
         => GND_net_1, B_DIN(13) => GND_net_1, B_DIN(12) => 
        GND_net_1, B_DIN(11) => GND_net_1, B_DIN(10) => GND_net_1, 
        B_DIN(9) => GND_net_1, B_DIN(8) => GND_net_1, B_DIN(7)
         => CoreAPB3_0_APBmslave0_PWDATA(7), B_DIN(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), B_DIN(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), B_DIN(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), B_DIN(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), B_DIN(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), B_DIN(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), B_DIN(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), B_ADDR(13) => 
        fifo_MEMWADDR(10), B_ADDR(12) => fifo_MEMWADDR(9), 
        B_ADDR(11) => fifo_MEMWADDR(8), B_ADDR(10) => 
        fifo_MEMWADDR(7), B_ADDR(9) => fifo_MEMWADDR(6), 
        B_ADDR(8) => fifo_MEMWADDR(5), B_ADDR(7) => 
        fifo_MEMWADDR(4), B_ADDR(6) => fifo_MEMWADDR(3), 
        B_ADDR(5) => fifo_MEMWADDR(2), B_ADDR(4) => 
        fifo_MEMWADDR(1), B_ADDR(3) => fifo_MEMWADDR(0), 
        B_ADDR(2) => GND_net_1, B_ADDR(1) => GND_net_1, B_ADDR(0)
         => GND_net_1, B_WEN(1) => GND_net_1, B_WEN(0) => 
        VCC_net_1, A_EN => VCC_net_1, A_DOUT_LAT => VCC_net_1, 
        A_WIDTH(2) => GND_net_1, A_WIDTH(1) => VCC_net_1, 
        A_WIDTH(0) => VCC_net_1, A_WMODE => GND_net_1, B_EN => 
        VCC_net_1, B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => 
        GND_net_1, B_WIDTH(1) => VCC_net_1, B_WIDTH(0) => 
        VCC_net_1, B_WMODE => GND_net_1, SII_LOCK => GND_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_2Kx8_FIFO_2Kx8_0_ram_wrapper is

    port( RDATA_int                    : out   std_logic_vector(7 downto 0);
          fifo_MEMRADDR                : in    std_logic_vector(10 downto 0);
          CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0);
          fifo_MEMWADDR                : in    std_logic_vector(10 downto 0);
          BIT_CLK                      : in    std_logic;
          N_19_i                       : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic;
          fifo_MEMWE                   : in    std_logic
        );

end FIFO_2Kx8_FIFO_2Kx8_0_ram_wrapper;

architecture DEF_ARCH of FIFO_2Kx8_FIFO_2Kx8_0_ram_wrapper is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component FIFO_2Kx8_FIFO_2Kx8_0_LSRAM_top
    port( fifo_MEMWADDR                : in    std_logic_vector(10 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0) := (others => 'U');
          fifo_MEMRADDR                : in    std_logic_vector(10 downto 0) := (others => 'U');
          RDATA_int                    : out   std_logic_vector(7 downto 0);
          fifo_MEMWE                   : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic := 'U';
          N_19_i                       : in    std_logic := 'U';
          BIT_CLK                      : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : FIFO_2Kx8_FIFO_2Kx8_0_LSRAM_top
	Use entity work.FIFO_2Kx8_FIFO_2Kx8_0_LSRAM_top(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    L1_asyncnonpipe : FIFO_2Kx8_FIFO_2Kx8_0_LSRAM_top
      port map(fifo_MEMWADDR(10) => fifo_MEMWADDR(10), 
        fifo_MEMWADDR(9) => fifo_MEMWADDR(9), fifo_MEMWADDR(8)
         => fifo_MEMWADDR(8), fifo_MEMWADDR(7) => 
        fifo_MEMWADDR(7), fifo_MEMWADDR(6) => fifo_MEMWADDR(6), 
        fifo_MEMWADDR(5) => fifo_MEMWADDR(5), fifo_MEMWADDR(4)
         => fifo_MEMWADDR(4), fifo_MEMWADDR(3) => 
        fifo_MEMWADDR(3), fifo_MEMWADDR(2) => fifo_MEMWADDR(2), 
        fifo_MEMWADDR(1) => fifo_MEMWADDR(1), fifo_MEMWADDR(0)
         => fifo_MEMWADDR(0), CoreAPB3_0_APBmslave0_PWDATA(7) => 
        CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), fifo_MEMRADDR(10) => 
        fifo_MEMRADDR(10), fifo_MEMRADDR(9) => fifo_MEMRADDR(9), 
        fifo_MEMRADDR(8) => fifo_MEMRADDR(8), fifo_MEMRADDR(7)
         => fifo_MEMRADDR(7), fifo_MEMRADDR(6) => 
        fifo_MEMRADDR(6), fifo_MEMRADDR(5) => fifo_MEMRADDR(5), 
        fifo_MEMRADDR(4) => fifo_MEMRADDR(4), fifo_MEMRADDR(3)
         => fifo_MEMRADDR(3), fifo_MEMRADDR(2) => 
        fifo_MEMRADDR(2), fifo_MEMRADDR(1) => fifo_MEMRADDR(1), 
        fifo_MEMRADDR(0) => fifo_MEMRADDR(0), RDATA_int(7) => 
        RDATA_int(7), RDATA_int(6) => RDATA_int(6), RDATA_int(5)
         => RDATA_int(5), RDATA_int(4) => RDATA_int(4), 
        RDATA_int(3) => RDATA_int(3), RDATA_int(2) => 
        RDATA_int(2), RDATA_int(1) => RDATA_int(1), RDATA_int(0)
         => RDATA_int(0), fifo_MEMWE => fifo_MEMWE, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz, 
        N_19_i => N_19_i, BIT_CLK => BIT_CLK);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv_0 is

    port( wptr_bin_sync  : inout std_logic_vector(11 downto 0) := (others => 'Z');
          wptr_gray_sync : in    std_logic_vector(10 downto 0);
          bin_N_4_0_i    : out   std_logic
        );

end FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv_0;

architecture DEF_ARCH of 
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv_0 is 

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \bin_m3_0_3\, \bin_m3_0_2\, GND_net_1, VCC_net_1
         : std_logic;

begin 


    \bin_out_xhdl1_i_o2_RNIS01B2[10]\ : CFG3
      generic map(INIT => x"69")

      port map(A => \bin_m3_0_3\, B => \bin_m3_0_2\, C => 
        wptr_bin_sync(10), Y => bin_N_4_0_i);
    
    \bin_out_xhdl1_0_a2[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => wptr_bin_sync(2), B => wptr_gray_sync(1), Y
         => wptr_bin_sync(1));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \bin_out_xhdl1_0_a2[5]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(7), B => wptr_bin_sync(8), C
         => wptr_gray_sync(6), D => wptr_gray_sync(5), Y => 
        wptr_bin_sync(5));
    
    \bin_out_xhdl1_0_a2[2]\ : CFG4
      generic map(INIT => x"9669")

      port map(A => wptr_bin_sync(10), B => \bin_m3_0_3\, C => 
        wptr_gray_sync(2), D => \bin_m3_0_2\, Y => 
        wptr_bin_sync(2));
    
    \bin_out_xhdl1_0_a2[0]\ : CFG3
      generic map(INIT => x"96")

      port map(A => wptr_gray_sync(1), B => wptr_bin_sync(2), C
         => wptr_gray_sync(0), Y => wptr_bin_sync(0));
    
    \bin_out_xhdl1_i_o2[9]\ : CFG3
      generic map(INIT => x"96")

      port map(A => wptr_gray_sync(9), B => wptr_bin_sync(11), C
         => wptr_gray_sync(10), Y => wptr_bin_sync(9));
    
    \bin_out_xhdl1_i_o2[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => wptr_bin_sync(11), B => wptr_gray_sync(10), Y
         => wptr_bin_sync(10));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \bin_out_xhdl1_0_a2[6]\ : CFG3
      generic map(INIT => x"96")

      port map(A => wptr_gray_sync(6), B => wptr_gray_sync(7), C
         => wptr_bin_sync(8), Y => wptr_bin_sync(6));
    
    \bin_out_xhdl1_0_a2[4]\ : CFG3
      generic map(INIT => x"96")

      port map(A => wptr_gray_sync(5), B => wptr_bin_sync(6), C
         => wptr_gray_sync(4), Y => wptr_bin_sync(4));
    
    bin_m3_0_2 : CFG3
      generic map(INIT => x"96")

      port map(A => wptr_gray_sync(3), B => wptr_gray_sync(6), C
         => wptr_gray_sync(7), Y => \bin_m3_0_2\);
    
    \bin_out_xhdl1_0_a2[8]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(10), B => wptr_bin_sync(11), C
         => wptr_gray_sync(8), D => wptr_gray_sync(9), Y => 
        wptr_bin_sync(8));
    
    bin_m3_0_3 : CFG4
      generic map(INIT => x"9669")

      port map(A => wptr_gray_sync(8), B => wptr_gray_sync(4), C
         => wptr_gray_sync(9), D => wptr_gray_sync(5), Y => 
        \bin_m3_0_3\);
    
    \bin_out_xhdl1_0_a2[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => wptr_bin_sync(8), B => wptr_gray_sync(7), Y
         => wptr_bin_sync(7));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_1 is

    port( wptr_gray       : in    std_logic_vector(11 downto 0);
          wptr_gray_sync  : out   std_logic_vector(10 downto 0);
          wptr_bin_sync_0 : out   std_logic;
          BIT_CLK         : in    std_logic;
          itx_fifo_rst_i  : in    std_logic
        );

end FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_1;

architecture DEF_ARCH of 
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_1 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \sync_int[7]_net_1\, GND_net_1, 
        \sync_int[8]_net_1\, \sync_int[9]_net_1\, 
        \sync_int[10]_net_1\, \sync_int[11]_net_1\, 
        \sync_int[4]_net_1\, \sync_int[5]_net_1\, 
        \sync_int[6]_net_1\, \sync_int[0]_net_1\, 
        \sync_int[1]_net_1\, \sync_int[2]_net_1\, 
        \sync_int[3]_net_1\ : std_logic;

begin 


    \sync_int[9]\ : SLE
      port map(D => wptr_gray(9), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[9]_net_1\);
    
    \sync_int[4]\ : SLE
      port map(D => wptr_gray(4), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[4]_net_1\);
    
    \sync_out_xhdl1[10]\ : SLE
      port map(D => \sync_int[10]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(10));
    
    \sync_int[1]\ : SLE
      port map(D => wptr_gray(1), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[1]_net_1\);
    
    \sync_int[11]\ : SLE
      port map(D => wptr_gray(11), CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[11]_net_1\);
    
    \sync_out_xhdl1[6]\ : SLE
      port map(D => \sync_int[6]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(6));
    
    \sync_out_xhdl1[3]\ : SLE
      port map(D => \sync_int[3]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(3));
    
    \sync_int[6]\ : SLE
      port map(D => wptr_gray(6), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[6]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \sync_out_xhdl1[11]\ : SLE
      port map(D => \sync_int[11]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_bin_sync_0);
    
    \sync_int[3]\ : SLE
      port map(D => wptr_gray(3), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[3]_net_1\);
    
    \sync_out_xhdl1[4]\ : SLE
      port map(D => \sync_int[4]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(4));
    
    \sync_int[0]\ : SLE
      port map(D => wptr_gray(0), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[0]_net_1\);
    
    \sync_out_xhdl1[1]\ : SLE
      port map(D => \sync_int[1]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(1));
    
    \sync_int[5]\ : SLE
      port map(D => wptr_gray(5), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[5]_net_1\);
    
    \sync_int[2]\ : SLE
      port map(D => wptr_gray(2), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[2]_net_1\);
    
    \sync_out_xhdl1[9]\ : SLE
      port map(D => \sync_int[9]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(9));
    
    \sync_out_xhdl1[2]\ : SLE
      port map(D => \sync_int[2]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(2));
    
    \sync_int[8]\ : SLE
      port map(D => wptr_gray(8), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[8]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sync_out_xhdl1[7]\ : SLE
      port map(D => \sync_int[7]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(7));
    
    \sync_out_xhdl1[5]\ : SLE
      port map(D => \sync_int[5]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(5));
    
    \sync_out_xhdl1[0]\ : SLE
      port map(D => \sync_int[0]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(0));
    
    \sync_out_xhdl1[8]\ : SLE
      port map(D => \sync_int[8]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        wptr_gray_sync(8));
    
    \sync_int[7]\ : SLE
      port map(D => wptr_gray(7), CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[7]_net_1\);
    
    \sync_int[10]\ : SLE
      port map(D => wptr_gray(10), CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_0 is

    port( rptr_gray                 : in    std_logic_vector(11 downto 0);
          rptr_gray_sync            : out   std_logic_vector(10 downto 0);
          rptr_bin_sync_0           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          itx_fifo_rst_i            : in    std_logic
        );

end FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_0;

architecture DEF_ARCH of 
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_0 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \sync_int[10]_net_1\, VCC_net_1, GND_net_1, 
        \sync_int[11]_net_1\, \sync_int[0]_net_1\, 
        \sync_int[1]_net_1\, \sync_int[2]_net_1\, 
        \sync_int[3]_net_1\, \sync_int[4]_net_1\, 
        \sync_int[5]_net_1\, \sync_int[6]_net_1\, 
        \sync_int[7]_net_1\, \sync_int[8]_net_1\, 
        \sync_int[9]_net_1\ : std_logic;

begin 


    \sync_int[9]\ : SLE
      port map(D => rptr_gray(9), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[9]_net_1\);
    
    \sync_int[4]\ : SLE
      port map(D => rptr_gray(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[4]_net_1\);
    
    \sync_out_xhdl1[10]\ : SLE
      port map(D => \sync_int[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(10));
    
    \sync_int[1]\ : SLE
      port map(D => rptr_gray(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[1]_net_1\);
    
    \sync_int[11]\ : SLE
      port map(D => rptr_gray(11), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[11]_net_1\);
    
    \sync_out_xhdl1[6]\ : SLE
      port map(D => \sync_int[6]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(6));
    
    \sync_out_xhdl1[3]\ : SLE
      port map(D => \sync_int[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(3));
    
    \sync_int[6]\ : SLE
      port map(D => rptr_gray(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[6]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \sync_out_xhdl1[11]\ : SLE
      port map(D => \sync_int[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_bin_sync_0);
    
    \sync_int[3]\ : SLE
      port map(D => rptr_gray(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[3]_net_1\);
    
    \sync_out_xhdl1[4]\ : SLE
      port map(D => \sync_int[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(4));
    
    \sync_int[0]\ : SLE
      port map(D => rptr_gray(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[0]_net_1\);
    
    \sync_out_xhdl1[1]\ : SLE
      port map(D => \sync_int[1]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(1));
    
    \sync_int[5]\ : SLE
      port map(D => rptr_gray(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[5]_net_1\);
    
    \sync_int[2]\ : SLE
      port map(D => rptr_gray(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[2]_net_1\);
    
    \sync_out_xhdl1[9]\ : SLE
      port map(D => \sync_int[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(9));
    
    \sync_out_xhdl1[2]\ : SLE
      port map(D => \sync_int[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(2));
    
    \sync_int[8]\ : SLE
      port map(D => rptr_gray(8), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[8]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sync_out_xhdl1[7]\ : SLE
      port map(D => \sync_int[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(7));
    
    \sync_out_xhdl1[5]\ : SLE
      port map(D => \sync_int[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(5));
    
    \sync_out_xhdl1[0]\ : SLE
      port map(D => \sync_int[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(0));
    
    \sync_out_xhdl1[8]\ : SLE
      port map(D => \sync_int[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(8));
    
    \sync_int[7]\ : SLE
      port map(D => rptr_gray(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[7]_net_1\);
    
    \sync_int[10]\ : SLE
      port map(D => rptr_gray(10), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[10]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv is

    port( rptr_bin_sync  : inout std_logic_vector(11 downto 0) := (others => 'Z');
          rptr_gray_sync : in    std_logic_vector(10 downto 0)
        );

end FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv;

architecture DEF_ARCH of 
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    \bin_out_xhdl1_0_a2[1]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(3), B => rptr_gray_sync(1), C
         => rptr_bin_sync(4), D => rptr_gray_sync(2), Y => 
        rptr_bin_sync(1));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \bin_out_xhdl1_0_a2[5]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(7), B => rptr_gray_sync(6), C
         => rptr_gray_sync(5), D => rptr_bin_sync(8), Y => 
        rptr_bin_sync(5));
    
    \bin_out_xhdl1_0_a2[2]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(4), B => rptr_gray_sync(3), C
         => rptr_gray_sync(2), D => rptr_bin_sync(5), Y => 
        rptr_bin_sync(2));
    
    \bin_out_xhdl1_0_a2[0]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(2), B => rptr_bin_sync(3), C
         => rptr_gray_sync(0), D => rptr_gray_sync(1), Y => 
        rptr_bin_sync(0));
    
    \bin_out_xhdl1_i_o2[9]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(10), B => rptr_gray_sync(9), C
         => rptr_bin_sync(11), Y => rptr_bin_sync(9));
    
    \bin_out_xhdl1_i_o2[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(11), B => rptr_gray_sync(10), Y
         => rptr_bin_sync(10));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \bin_out_xhdl1_0_a2[6]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(8), B => rptr_gray_sync(7), C
         => rptr_gray_sync(6), D => rptr_bin_sync(9), Y => 
        rptr_bin_sync(6));
    
    \bin_out_xhdl1_0_a2[4]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(6), B => rptr_gray_sync(5), C
         => rptr_gray_sync(4), D => rptr_bin_sync(7), Y => 
        rptr_bin_sync(4));
    
    \bin_out_xhdl1_0_a2[8]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(10), B => rptr_gray_sync(9), C
         => rptr_gray_sync(8), D => rptr_bin_sync(11), Y => 
        rptr_bin_sync(8));
    
    \bin_out_xhdl1_0_a2[7]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(9), B => rptr_gray_sync(8), C
         => rptr_gray_sync(7), D => rptr_bin_sync(10), Y => 
        rptr_bin_sync(7));
    
    \bin_out_xhdl1_0_a2[3]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(5), B => rptr_gray_sync(4), C
         => rptr_gray_sync(3), D => rptr_bin_sync(6), Y => 
        rptr_bin_sync(3));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_2Kx8_FIFO_2Kx8_0_corefifo_async is

    port( fifo_MEMWADDR             : out   std_logic_vector(10 downto 0);
          fifo_MEMRADDR             : out   std_logic_vector(10 downto 0);
          N_114                     : in    std_logic;
          TX_FIFO_wr_en             : in    std_logic;
          fifo_MEMWE                : out   std_logic;
          N_19_i                    : out   std_logic;
          TX_FIFO_Full              : out   std_logic;
          TX_FIFO_Empty             : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          BIT_CLK                   : in    std_logic;
          itx_fifo_rst_i            : in    std_logic;
          TX_FIFO_OVERFLOW_i        : out   std_logic;
          TX_FIFO_OVERFLOW          : out   std_logic;
          TX_FIFO_UNDERRUN_i        : out   std_logic;
          TX_FIFO_UNDERRUN          : out   std_logic
        );

end FIFO_2Kx8_FIFO_2Kx8_0_corefifo_async;

architecture DEF_ARCH of FIFO_2Kx8_FIFO_2Kx8_0_corefifo_async is 

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv_0
    port( wptr_bin_sync  : inout   std_logic_vector(11 downto 0);
          wptr_gray_sync : in    std_logic_vector(10 downto 0) := (others => 'U');
          bin_N_4_0_i    : out   std_logic
        );
  end component;

  component FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_1
    port( wptr_gray       : in    std_logic_vector(11 downto 0) := (others => 'U');
          wptr_gray_sync  : out   std_logic_vector(10 downto 0);
          wptr_bin_sync_0 : out   std_logic;
          BIT_CLK         : in    std_logic := 'U';
          itx_fifo_rst_i  : in    std_logic := 'U'
        );
  end component;

  component FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_0
    port( rptr_gray                 : in    std_logic_vector(11 downto 0) := (others => 'U');
          rptr_gray_sync            : out   std_logic_vector(10 downto 0);
          rptr_bin_sync_0           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          itx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv
    port( rptr_bin_sync  : inout   std_logic_vector(11 downto 0);
          rptr_gray_sync : in    std_logic_vector(10 downto 0) := (others => 'U')
        );
  end component;

    signal \wptr[0]_net_1\, \wptr_s[0]\, \fifo_MEMWADDR[0]\, 
        \memwaddr_r_s[0]\, \fifo_MEMRADDR[0]\, \memraddr_r_s[0]\, 
        \rptr[0]_net_1\, \rptr_s[0]\, \TX_FIFO_UNDERRUN\, 
        \TX_FIFO_OVERFLOW\, \rptr_gray[7]_net_1\, VCC_net_1, 
        \rptr_gray_1[7]_net_1\, GND_net_1, \rptr_gray[8]_net_1\, 
        \rptr_gray_1[8]_net_1\, \rptr_gray[9]_net_1\, 
        \rptr_gray_1[9]_net_1\, \rptr_gray[10]_net_1\, 
        \rptr_gray_1[10]_net_1\, \rptr_gray[11]_net_1\, 
        \rptr[11]_net_1\, \wptr_gray[4]_net_1\, 
        \wptr_gray_1[4]_net_1\, \wptr_gray[5]_net_1\, 
        \wptr_gray_1[5]_net_1\, \wptr_gray[6]_net_1\, 
        \wptr_gray_1[6]_net_1\, \wptr_gray[7]_net_1\, 
        \wptr_gray_1[7]_net_1\, \wptr_gray[8]_net_1\, 
        \wptr_gray_1[8]_net_1\, \wptr_gray[9]_net_1\, 
        \wptr_gray_1[9]_net_1\, \wptr_gray[10]_net_1\, 
        \wptr_gray_1[10]_net_1\, \wptr_gray[11]_net_1\, 
        \wptr[11]_net_1\, \rptr_gray[0]_net_1\, 
        \rptr_gray_1[0]_net_1\, \rptr_gray[1]_net_1\, 
        \rptr_gray_1[1]_net_1\, \rptr_gray[2]_net_1\, 
        \rptr_gray_1[2]_net_1\, \rptr_gray[3]_net_1\, 
        \rptr_gray_1[3]_net_1\, \rptr_gray[4]_net_1\, 
        \rptr_gray_1[4]_net_1\, \rptr_gray[5]_net_1\, 
        \rptr_gray_1[5]_net_1\, \rptr_gray[6]_net_1\, 
        \rptr_gray_1[6]_net_1\, \rptr_bin_sync2[1]_net_1\, 
        \rptr_bin_sync[1]\, \rptr_bin_sync2[2]_net_1\, 
        \rptr_bin_sync[2]\, \rptr_bin_sync2[3]_net_1\, 
        \rptr_bin_sync[3]\, \rptr_bin_sync2[4]_net_1\, 
        \rptr_bin_sync[4]\, \rptr_bin_sync2[5]_net_1\, 
        \rptr_bin_sync[5]\, \rptr_bin_sync2[6]_net_1\, 
        \rptr_bin_sync[6]\, \rptr_bin_sync2[7]_net_1\, 
        \rptr_bin_sync[7]\, \rptr_bin_sync2[8]_net_1\, 
        \rptr_bin_sync[8]\, \rptr_bin_sync2[9]_net_1\, 
        \rptr_bin_sync[9]\, \rptr_bin_sync2[10]_net_1\, 
        \rptr_bin_sync[10]\, \rptr_bin_sync2[11]_net_1\, 
        \rptr_bin_sync[11]\, \wptr_gray[0]_net_1\, 
        \wptr_gray_1[0]_net_1\, \wptr_gray[1]_net_1\, 
        \wptr_gray_1[1]_net_1\, \wptr_gray[2]_net_1\, 
        \wptr_gray_1[2]_net_1\, \wptr_gray[3]_net_1\, 
        \wptr_gray_1[3]_net_1\, \rptr_bin_sync2[0]_net_1\, 
        \rptr_bin_sync[0]\, \wptr_bin_sync2[1]_net_1\, 
        \wptr_bin_sync[1]\, \wptr_bin_sync2[2]_net_1\, 
        \wptr_bin_sync[2]\, \wptr_bin_sync2[3]_net_1\, 
        bin_N_4_0_i, \wptr_bin_sync2[4]_net_1\, 
        \wptr_bin_sync[4]\, \wptr_bin_sync2[5]_net_1\, 
        \wptr_bin_sync[5]\, \wptr_bin_sync2[6]_net_1\, 
        \wptr_bin_sync[6]\, \wptr_bin_sync2[7]_net_1\, 
        \wptr_bin_sync[7]\, \wptr_bin_sync2[8]_net_1\, 
        \wptr_bin_sync[8]\, \wptr_bin_sync2[9]_net_1\, 
        \wptr_bin_sync[9]\, \wptr_bin_sync2[10]_net_1\, 
        \wptr_bin_sync[10]\, \wptr_bin_sync2[11]_net_1\, 
        \wptr_bin_sync[11]\, rdiff_bus, \wptr_bin_sync[0]\, 
        N_12_i, N_7_i, \TX_FIFO_Empty\, empty_r_3, \TX_FIFO_Full\, 
        fulli, \N_19_i\, \rptr[1]_net_1\, \rptr_s[1]\, 
        \rptr[2]_net_1\, \rptr_s[2]\, \rptr[3]_net_1\, 
        \rptr_s[3]\, \rptr[4]_net_1\, \rptr_s[4]\, 
        \rptr[5]_net_1\, \rptr_s[5]\, \rptr[6]_net_1\, 
        \rptr_s[6]\, \rptr[7]_net_1\, \rptr_s[7]\, 
        \rptr[8]_net_1\, \rptr_s[8]\, \rptr[9]_net_1\, 
        \rptr_s[9]\, \rptr[10]_net_1\, \rptr_s[10]\, 
        \rptr_s[11]_net_1\, \fifo_MEMRADDR[1]\, \memraddr_r_s[1]\, 
        \fifo_MEMRADDR[2]\, \memraddr_r_s[2]\, \fifo_MEMRADDR[3]\, 
        \memraddr_r_s[3]\, \fifo_MEMRADDR[4]\, \memraddr_r_s[4]\, 
        \fifo_MEMRADDR[5]\, \memraddr_r_s[5]\, \fifo_MEMRADDR[6]\, 
        \memraddr_r_s[6]\, \fifo_MEMRADDR[7]\, \memraddr_r_s[7]\, 
        \fifo_MEMRADDR[8]\, \memraddr_r_s[8]\, \fifo_MEMRADDR[9]\, 
        \memraddr_r_s[9]\, \fifo_MEMRADDR[10]\, 
        \memraddr_r_s[10]_net_1\, \fifo_MEMWE\, 
        \fifo_MEMWADDR[1]\, \memwaddr_r_s[1]\, \fifo_MEMWADDR[2]\, 
        \memwaddr_r_s[2]\, \fifo_MEMWADDR[3]\, \memwaddr_r_s[3]\, 
        \fifo_MEMWADDR[4]\, \memwaddr_r_s[4]\, \fifo_MEMWADDR[5]\, 
        \memwaddr_r_s[5]\, \fifo_MEMWADDR[6]\, \memwaddr_r_s[6]\, 
        \fifo_MEMWADDR[7]\, \memwaddr_r_s[7]\, \fifo_MEMWADDR[8]\, 
        \memwaddr_r_s[8]\, \fifo_MEMWADDR[9]\, \memwaddr_r_s[9]\, 
        \fifo_MEMWADDR[10]\, \memwaddr_r_s[10]_net_1\, 
        \wptr[1]_net_1\, \wptr_s[1]\, \wptr[2]_net_1\, 
        \wptr_s[2]\, \wptr[3]_net_1\, \wptr_s[3]\, 
        \wptr[4]_net_1\, \wptr_s[4]\, \wptr[5]_net_1\, 
        \wptr_s[5]\, \wptr[6]_net_1\, \wptr_s[6]\, 
        \wptr[7]_net_1\, \wptr_s[7]\, \wptr[8]_net_1\, 
        \wptr_s[8]\, \wptr[9]_net_1\, \wptr_s[9]\, 
        \wptr[10]_net_1\, \wptr_s[10]\, \wptr_s[11]_net_1\, 
        \wdiff_bus_cry_0\, wdiff_bus_cry_0_Y, \wdiff_bus_cry_1\, 
        \wdiff_bus[1]\, \wdiff_bus_cry_2\, \wdiff_bus[2]\, 
        \wdiff_bus_cry_3\, \wdiff_bus[3]\, \wdiff_bus_cry_4\, 
        \wdiff_bus[4]\, \wdiff_bus_cry_5\, \wdiff_bus[5]\, 
        \wdiff_bus_cry_6\, \wdiff_bus[6]\, \wdiff_bus_cry_7\, 
        \wdiff_bus[7]\, \wdiff_bus_cry_8\, \wdiff_bus[8]\, 
        \wdiff_bus_cry_9\, \wdiff_bus[9]\, \wdiff_bus[11]\, 
        \wdiff_bus_cry_10\, \wdiff_bus[10]\, \rdiff_bus_cry_0\, 
        rdiff_bus_cry_0_Y, \rdiff_bus_cry_1\, \rdiff_bus[1]\, 
        \rdiff_bus_cry_2\, \rdiff_bus[2]\, \rdiff_bus_cry_3\, 
        \rdiff_bus[3]\, \rdiff_bus_cry_4\, \rdiff_bus[4]\, 
        \rdiff_bus_cry_5\, \rdiff_bus[5]\, \rdiff_bus_cry_6\, 
        \rdiff_bus[6]\, \rdiff_bus_cry_7\, \rdiff_bus[7]\, 
        \rdiff_bus_cry_8\, \rdiff_bus[8]\, \rdiff_bus_cry_9\, 
        \rdiff_bus[9]\, \rdiff_bus[11]\, \rdiff_bus_cry_10\, 
        \rdiff_bus[10]\, wptr_s_910_FCO, \wptr_cry[1]_net_1\, 
        \wptr_cry[2]_net_1\, \wptr_cry[3]_net_1\, 
        \wptr_cry[4]_net_1\, \wptr_cry[5]_net_1\, 
        \wptr_cry[6]_net_1\, \wptr_cry[7]_net_1\, 
        \wptr_cry[8]_net_1\, \wptr_cry[9]_net_1\, 
        \wptr_cry[10]_net_1\, memwaddr_r_s_911_FCO, 
        \memwaddr_r_cry[1]_net_1\, \memwaddr_r_cry[2]_net_1\, 
        \memwaddr_r_cry[3]_net_1\, \memwaddr_r_cry[4]_net_1\, 
        \memwaddr_r_cry[5]_net_1\, \memwaddr_r_cry[6]_net_1\, 
        \memwaddr_r_cry[7]_net_1\, \memwaddr_r_cry[8]_net_1\, 
        \memwaddr_r_cry[9]_net_1\, memraddr_r_s_912_FCO, 
        \memraddr_r_cry[1]_net_1\, \memraddr_r_cry[2]_net_1\, 
        \memraddr_r_cry[3]_net_1\, \memraddr_r_cry[4]_net_1\, 
        \memraddr_r_cry[5]_net_1\, \memraddr_r_cry[6]_net_1\, 
        \memraddr_r_cry[7]_net_1\, \memraddr_r_cry[8]_net_1\, 
        \memraddr_r_cry[9]_net_1\, rptr_s_913_FCO, 
        \rptr_cry[1]_net_1\, \rptr_cry[2]_net_1\, 
        \rptr_cry[3]_net_1\, \rptr_cry[4]_net_1\, 
        \rptr_cry[5]_net_1\, \rptr_cry[6]_net_1\, 
        \rptr_cry[7]_net_1\, \rptr_cry[8]_net_1\, 
        \rptr_cry[9]_net_1\, \rptr_cry[10]_net_1\, 
        empty_r_3_0_a3_2, empty_r_3_0_a3_7, empty_r_3_0_a3_5, 
        \fulli_0_a3_8\, \fulli_0_a3_7\, empty_r_3_0_a3_9, 
        \fulli_0_a3_6\, \wptr_gray_sync[0]\, \wptr_gray_sync[1]\, 
        \wptr_gray_sync[2]\, \wptr_gray_sync[3]\, 
        \wptr_gray_sync[4]\, \wptr_gray_sync[5]\, 
        \wptr_gray_sync[6]\, \wptr_gray_sync[7]\, 
        \wptr_gray_sync[8]\, \wptr_gray_sync[9]\, 
        \wptr_gray_sync[10]\, \rptr_gray_sync[0]\, 
        \rptr_gray_sync[1]\, \rptr_gray_sync[2]\, 
        \rptr_gray_sync[3]\, \rptr_gray_sync[4]\, 
        \rptr_gray_sync[5]\, \rptr_gray_sync[6]\, 
        \rptr_gray_sync[7]\, \rptr_gray_sync[8]\, 
        \rptr_gray_sync[9]\, \rptr_gray_sync[10]\ : std_logic;
    signal nc1 : std_logic;

    for all : FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv_0
	Use entity work.
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv_0(DEF_ARCH);
    for all : FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_1
	Use entity work.
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_1(DEF_ARCH);
    for all : FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_0
	Use entity work.
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_0(DEF_ARCH);
    for all : FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv
	Use entity work.
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv(DEF_ARCH);
begin 

    fifo_MEMWADDR(10) <= \fifo_MEMWADDR[10]\;
    fifo_MEMWADDR(9) <= \fifo_MEMWADDR[9]\;
    fifo_MEMWADDR(8) <= \fifo_MEMWADDR[8]\;
    fifo_MEMWADDR(7) <= \fifo_MEMWADDR[7]\;
    fifo_MEMWADDR(6) <= \fifo_MEMWADDR[6]\;
    fifo_MEMWADDR(5) <= \fifo_MEMWADDR[5]\;
    fifo_MEMWADDR(4) <= \fifo_MEMWADDR[4]\;
    fifo_MEMWADDR(3) <= \fifo_MEMWADDR[3]\;
    fifo_MEMWADDR(2) <= \fifo_MEMWADDR[2]\;
    fifo_MEMWADDR(1) <= \fifo_MEMWADDR[1]\;
    fifo_MEMWADDR(0) <= \fifo_MEMWADDR[0]\;
    fifo_MEMRADDR(10) <= \fifo_MEMRADDR[10]\;
    fifo_MEMRADDR(9) <= \fifo_MEMRADDR[9]\;
    fifo_MEMRADDR(8) <= \fifo_MEMRADDR[8]\;
    fifo_MEMRADDR(7) <= \fifo_MEMRADDR[7]\;
    fifo_MEMRADDR(6) <= \fifo_MEMRADDR[6]\;
    fifo_MEMRADDR(5) <= \fifo_MEMRADDR[5]\;
    fifo_MEMRADDR(4) <= \fifo_MEMRADDR[4]\;
    fifo_MEMRADDR(3) <= \fifo_MEMRADDR[3]\;
    fifo_MEMRADDR(2) <= \fifo_MEMRADDR[2]\;
    fifo_MEMRADDR(1) <= \fifo_MEMRADDR[1]\;
    fifo_MEMRADDR(0) <= \fifo_MEMRADDR[0]\;
    fifo_MEMWE <= \fifo_MEMWE\;
    N_19_i <= \N_19_i\;
    TX_FIFO_Full <= \TX_FIFO_Full\;
    TX_FIFO_Empty <= \TX_FIFO_Empty\;
    TX_FIFO_OVERFLOW <= \TX_FIFO_OVERFLOW\;
    TX_FIFO_UNDERRUN <= \TX_FIFO_UNDERRUN\;

    \rptr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[4]_net_1\, S
         => \rptr_s[5]\, Y => OPEN, FCO => \rptr_cry[5]_net_1\);
    
    \L1.empty_r_3_0_a3_9\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \rdiff_bus[3]\, B => \rdiff_bus[4]\, C => 
        empty_r_3_0_a3_2, D => empty_r_3_0_a3_7, Y => 
        empty_r_3_0_a3_9);
    
    underflow_r_RNIFFTA : CFG1
      generic map(INIT => "01")

      port map(A => \TX_FIFO_UNDERRUN\, Y => TX_FIFO_UNDERRUN_i);
    
    wdiff_bus_cry_8 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[8]_net_1\, B => 
        \rptr_bin_sync2[8]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_7\, S => \wdiff_bus[8]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_8\);
    
    \wptr_gray[4]\ : SLE
      port map(D => \wptr_gray_1[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[4]_net_1\);
    
    \rptr_gray_1[3]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[3]_net_1\, B => \rptr[4]_net_1\, Y => 
        \rptr_gray_1[3]_net_1\);
    
    \rptr_bin_sync2[6]\ : SLE
      port map(D => \rptr_bin_sync[6]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[6]_net_1\);
    
    \rptr[1]\ : SLE
      port map(D => \rptr_s[1]\, CLK => BIT_CLK, EN => \N_19_i\, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[1]_net_1\);
    
    \wptr_gray_1[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[9]_net_1\, B => \wptr[10]_net_1\, Y => 
        \wptr_gray_1[9]_net_1\);
    
    \rptr_gray_1[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[5]_net_1\, B => \rptr[6]_net_1\, Y => 
        \rptr_gray_1[5]_net_1\);
    
    \rptr_gray[9]\ : SLE
      port map(D => \rptr_gray_1[9]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[9]_net_1\);
    
    \rptr_gray[8]\ : SLE
      port map(D => \rptr_gray_1[8]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[8]_net_1\);
    
    \rptr_gray_1[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[2]_net_1\, B => \rptr[3]_net_1\, Y => 
        \rptr_gray_1[2]_net_1\);
    
    \rptr_bin_sync2[7]\ : SLE
      port map(D => \rptr_bin_sync[7]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[7]_net_1\);
    
    \memwaddr_r[1]\ : SLE
      port map(D => \memwaddr_r_s[1]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[1]\);
    
    \memwaddr_r_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[5]_net_1\, S => \memwaddr_r_s[6]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[6]_net_1\);
    
    \memwaddr_r_s[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[9]_net_1\, S => \memwaddr_r_s[10]_net_1\, 
        Y => OPEN, FCO => OPEN);
    
    \wptr_gray_1[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[7]_net_1\, B => \wptr[8]_net_1\, Y => 
        \wptr_gray_1[7]_net_1\);
    
    \memraddr_r[0]\ : SLE
      port map(D => \memraddr_r_s[0]\, CLK => BIT_CLK, EN => 
        \N_19_i\, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[0]\);
    
    \wptr[0]\ : SLE
      port map(D => \wptr_s[0]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[0]_net_1\);
    
    \rptr_bin_sync2[8]\ : SLE
      port map(D => \rptr_bin_sync[8]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[8]_net_1\);
    
    \rptr_gray_1[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[1]_net_1\, B => \rptr[2]_net_1\, Y => 
        \rptr_gray_1[1]_net_1\);
    
    \rptr_gray[10]\ : SLE
      port map(D => \rptr_gray_1[10]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[10]_net_1\);
    
    \wptr_gray_1[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[0]_net_1\, B => \wptr[1]_net_1\, Y => 
        \wptr_gray_1[0]_net_1\);
    
    wdiff_bus_cry_9 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[9]_net_1\, B => 
        \rptr_bin_sync2[9]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_8\, S => \wdiff_bus[9]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_9\);
    
    \rptr[5]\ : SLE
      port map(D => \rptr_s[5]\, CLK => BIT_CLK, EN => \N_19_i\, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[5]_net_1\);
    
    \rptr_gray[3]\ : SLE
      port map(D => \rptr_gray_1[3]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[3]_net_1\);
    
    \rptr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[5]_net_1\, S
         => \rptr_s[6]\, Y => OPEN, FCO => \rptr_cry[6]_net_1\);
    
    \memwaddr_r_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[1]\, C => 
        GND_net_1, D => GND_net_1, FCI => memwaddr_r_s_911_FCO, S
         => \memwaddr_r_s[1]\, Y => OPEN, FCO => 
        \memwaddr_r_cry[1]_net_1\);
    
    \L1.empty_r_3_0_a3\ : CFG4
      generic map(INIT => x"E000")

      port map(A => rdiff_bus_cry_0_Y, B => N_114, C => 
        empty_r_3_0_a3_5, D => empty_r_3_0_a3_9, Y => empty_r_3);
    
    \wptr_gray[3]\ : SLE
      port map(D => \wptr_gray_1[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[3]_net_1\);
    
    \rptr_gray_1[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[11]_net_1\, B => \rptr[10]_net_1\, Y
         => \rptr_gray_1[10]_net_1\);
    
    wdiff_bus_s_11 : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \rptr_bin_sync2[11]_net_1\, C
         => \wptr[11]_net_1\, D => GND_net_1, FCI => 
        \wdiff_bus_cry_10\, S => \wdiff_bus[11]\, Y => OPEN, FCO
         => OPEN);
    
    \rptr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[7]_net_1\, S
         => \rptr_s[8]\, Y => OPEN, FCO => \rptr_cry[8]_net_1\);
    
    \rptr[7]\ : SLE
      port map(D => \rptr_s[7]\, CLK => BIT_CLK, EN => \N_19_i\, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[7]_net_1\);
    
    rdiff_bus_cry_4 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[4]_net_1\, B => 
        \rptr[4]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_3\, S => \rdiff_bus[4]\, Y => OPEN, FCO
         => \rdiff_bus_cry_4\);
    
    \rptr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[9]_net_1\, S
         => \rptr_s[10]\, Y => OPEN, FCO => \rptr_cry[10]_net_1\);
    
    memwe_0_a3 : CFG2
      generic map(INIT => x"4")

      port map(A => \TX_FIFO_Full\, B => TX_FIFO_wr_en, Y => 
        \fifo_MEMWE\);
    
    \rptr_bin_sync2[0]\ : SLE
      port map(D => \rptr_bin_sync[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[0]_net_1\);
    
    \wptr[11]\ : SLE
      port map(D => \wptr_s[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \wptr[11]_net_1\);
    
    rdiff_bus_cry_1 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[1]_net_1\, B => 
        \rptr[1]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_0\, S => \rdiff_bus[1]\, Y => OPEN, FCO
         => \rdiff_bus_cry_1\);
    
    \memraddr_r[1]\ : SLE
      port map(D => \memraddr_r_s[1]\, CLK => BIT_CLK, EN => 
        \N_19_i\, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[1]\);
    
    \rptr_bin_sync2[2]\ : SLE
      port map(D => \rptr_bin_sync[2]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[2]_net_1\);
    
    rdiff_bus_cry_6 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[6]_net_1\, B => 
        \rptr[6]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_5\, S => \rdiff_bus[6]\, Y => OPEN, FCO
         => \rdiff_bus_cry_6\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \memwaddr_r_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[3]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[2]_net_1\, S => \memwaddr_r_s[3]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[3]_net_1\);
    
    \rptr_gray[1]\ : SLE
      port map(D => \rptr_gray_1[1]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[1]_net_1\);
    
    \memwaddr_r[7]\ : SLE
      port map(D => \memwaddr_r_s[7]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[7]\);
    
    \memraddr_r_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[2]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[1]_net_1\, S => \memraddr_r_s[2]\, Y => 
        OPEN, FCO => \memraddr_r_cry[2]_net_1\);
    
    \wptr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[3]_net_1\, S
         => \wptr_s[4]\, Y => OPEN, FCO => \wptr_cry[4]_net_1\);
    
    \L1.empty_r_3_0_a3_7\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \rdiff_bus[7]\, B => \rdiff_bus[8]\, C => 
        \rdiff_bus[9]\, D => \rdiff_bus[10]\, Y => 
        empty_r_3_0_a3_7);
    
    \memraddr_r_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[8]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[7]_net_1\, S => \memraddr_r_s[8]\, Y => 
        OPEN, FCO => \memraddr_r_cry[8]_net_1\);
    
    \wptr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[9]_net_1\, S
         => \wptr_s[10]\, Y => OPEN, FCO => \wptr_cry[10]_net_1\);
    
    wdiff_bus_cry_5 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[5]_net_1\, B => 
        \rptr_bin_sync2[5]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_4\, S => \wdiff_bus[5]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_5\);
    
    \memwaddr_r[4]\ : SLE
      port map(D => \memwaddr_r_s[4]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[4]\);
    
    \wptr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[1]_net_1\, S
         => \wptr_s[2]\, Y => OPEN, FCO => \wptr_cry[2]_net_1\);
    
    memraddr_r_s_912 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[0]\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => memraddr_r_s_912_FCO);
    
    wdiff_bus_cry_0 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[0]_net_1\, B => 
        \rptr_bin_sync2[0]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => VCC_net_1, S => OPEN, Y => wdiff_bus_cry_0_Y, FCO
         => \wdiff_bus_cry_0\);
    
    \wptr[1]\ : SLE
      port map(D => \wptr_s[1]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[1]_net_1\);
    
    \rptr_bin_sync2[4]\ : SLE
      port map(D => \rptr_bin_sync[4]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[4]_net_1\);
    
    \wptr_bin_sync2[6]\ : SLE
      port map(D => \wptr_bin_sync[6]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[6]_net_1\);
    
    \rptr[3]\ : SLE
      port map(D => \rptr_s[3]\, CLK => BIT_CLK, EN => \N_19_i\, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[3]_net_1\);
    
    \wptr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[2]_net_1\, S
         => \wptr_s[3]\, Y => OPEN, FCO => \wptr_cry[3]_net_1\);
    
    \rptr[6]\ : SLE
      port map(D => \rptr_s[6]\, CLK => BIT_CLK, EN => \N_19_i\, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[6]_net_1\);
    
    rdiff_bus_cry_8 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[8]_net_1\, B => 
        \rptr[8]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_7\, S => \rdiff_bus[8]\, Y => OPEN, FCO
         => \rdiff_bus_cry_8\);
    
    \wptr_gray[10]\ : SLE
      port map(D => \wptr_gray_1[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[10]_net_1\);
    
    rdiff_bus_cry_7 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[7]_net_1\, B => 
        \rptr[7]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_6\, S => \rdiff_bus[7]\, Y => OPEN, FCO
         => \rdiff_bus_cry_7\);
    
    \wptr_bin_sync2[7]\ : SLE
      port map(D => \wptr_bin_sync[7]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[7]_net_1\);
    
    overflow_r_RNIDBD3 : CFG1
      generic map(INIT => "01")

      port map(A => \TX_FIFO_OVERFLOW\, Y => TX_FIFO_OVERFLOW_i);
    
    \rptr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[8]_net_1\, S
         => \rptr_s[9]\, Y => OPEN, FCO => \rptr_cry[9]_net_1\);
    
    wptr_s_910 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => wptr_s_910_FCO);
    
    \rptr_gray[5]\ : SLE
      port map(D => \rptr_gray_1[5]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[5]_net_1\);
    
    \wptr_gray_1[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[2]_net_1\, B => \wptr[3]_net_1\, Y => 
        \wptr_gray_1[2]_net_1\);
    
    \wptr[5]\ : SLE
      port map(D => \wptr_s[5]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[5]_net_1\);
    
    rdiff_bus_cry_5 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[5]_net_1\, B => 
        \rptr[5]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_4\, S => \rdiff_bus[5]\, Y => OPEN, FCO
         => \rdiff_bus_cry_5\);
    
    \wptr_bin_sync2[8]\ : SLE
      port map(D => \wptr_bin_sync[8]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[8]_net_1\);
    
    \wptr[7]\ : SLE
      port map(D => \wptr_s[7]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[7]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \wptr_gray[1]\ : SLE
      port map(D => \wptr_gray_1[1]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[1]_net_1\);
    
    rptr_s_913 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => rptr_s_913_FCO);
    
    \rptr_gray_1[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[9]_net_1\, B => \rptr[10]_net_1\, Y => 
        \rptr_gray_1[9]_net_1\);
    
    \rptr_bin_sync2[5]\ : SLE
      port map(D => \rptr_bin_sync[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[5]_net_1\);
    
    \rptr_bin_sync2[1]\ : SLE
      port map(D => \rptr_bin_sync[1]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[1]_net_1\);
    
    \memwaddr_r[10]\ : SLE
      port map(D => \memwaddr_r_s[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[10]\);
    
    wdiff_bus_cry_7 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[7]_net_1\, B => 
        \rptr_bin_sync2[7]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_6\, S => \wdiff_bus[7]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_7\);
    
    \wptr_bin_sync2[0]\ : SLE
      port map(D => \wptr_bin_sync[0]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        rdiff_bus);
    
    rdiff_bus_s_11 : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \rptr[11]_net_1\, C => 
        \wptr_bin_sync2[11]_net_1\, D => GND_net_1, FCI => 
        \rdiff_bus_cry_10\, S => \rdiff_bus[11]\, Y => OPEN, FCO
         => OPEN);
    
    \memwaddr_r_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[8]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[7]_net_1\, S => \memwaddr_r_s[8]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[8]_net_1\);
    
    \wptr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => wptr_s_910_FCO, S => 
        \wptr_s[1]\, Y => OPEN, FCO => \wptr_cry[1]_net_1\);
    
    \memraddr_r[8]\ : SLE
      port map(D => \memraddr_r_s[8]\, CLK => BIT_CLK, EN => 
        \N_19_i\, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[8]\);
    
    \rptr[9]\ : SLE
      port map(D => \rptr_s[9]\, CLK => BIT_CLK, EN => \N_19_i\, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[9]_net_1\);
    
    \wptr_gray_1[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[6]_net_1\, B => \wptr[7]_net_1\, Y => 
        \wptr_gray_1[6]_net_1\);
    
    \wptr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[6]_net_1\, S
         => \wptr_s[7]\, Y => OPEN, FCO => \wptr_cry[7]_net_1\);
    
    \wptr_bin_sync2[2]\ : SLE
      port map(D => \wptr_bin_sync[2]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[2]_net_1\);
    
    \rptr_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \rptr[0]_net_1\, Y => \rptr_s[0]\);
    
    \rptr[4]\ : SLE
      port map(D => \rptr_s[4]\, CLK => BIT_CLK, EN => \N_19_i\, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[4]_net_1\);
    
    \memwaddr_r_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[4]_net_1\, S => \memwaddr_r_s[5]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[5]_net_1\);
    
    \memraddr_r_s[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[9]_net_1\, S => \memraddr_r_s[10]_net_1\, 
        Y => OPEN, FCO => OPEN);
    
    \wptr_gray[6]\ : SLE
      port map(D => \wptr_gray_1[6]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[6]_net_1\);
    
    \wptr_gray_1[3]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[3]_net_1\, B => \wptr[4]_net_1\, Y => 
        \wptr_gray_1[3]_net_1\);
    
    \wptr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[4]_net_1\, S
         => \wptr_s[5]\, Y => OPEN, FCO => \wptr_cry[5]_net_1\);
    
    \memraddr_r_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[4]_net_1\, S => \memraddr_r_s[5]\, Y => 
        OPEN, FCO => \memraddr_r_cry[5]_net_1\);
    
    \memraddr_r_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[1]\, C => 
        GND_net_1, D => GND_net_1, FCI => memraddr_r_s_912_FCO, S
         => \memraddr_r_s[1]\, Y => OPEN, FCO => 
        \memraddr_r_cry[1]_net_1\);
    
    \rptr_gray[4]\ : SLE
      port map(D => \rptr_gray_1[4]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[4]_net_1\);
    
    \wptr_bin_sync2[4]\ : SLE
      port map(D => \wptr_bin_sync[4]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[4]_net_1\);
    
    \wptr[3]\ : SLE
      port map(D => \wptr_s[3]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[3]_net_1\);
    
    \memwaddr_r[6]\ : SLE
      port map(D => \memwaddr_r_s[6]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[6]\);
    
    \wptr_s[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[10]_net_1\, S
         => \wptr_s[11]_net_1\, Y => OPEN, FCO => OPEN);
    
    \wptr[6]\ : SLE
      port map(D => \wptr_s[6]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[6]_net_1\);
    
    \memwaddr_r[9]\ : SLE
      port map(D => \memwaddr_r_s[9]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[9]\);
    
    \memraddr_r_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[3]_net_1\, S => \memraddr_r_s[4]\, Y => 
        OPEN, FCO => \memraddr_r_cry[4]_net_1\);
    
    \memraddr_r[10]\ : SLE
      port map(D => \memraddr_r_s[10]_net_1\, CLK => BIT_CLK, EN
         => \N_19_i\, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \fifo_MEMRADDR[10]\);
    
    \memwaddr_r[3]\ : SLE
      port map(D => \memwaddr_r_s[3]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[3]\);
    
    empty_r_RNI5ING : CFG2
      generic map(INIT => x"2")

      port map(A => N_114, B => \TX_FIFO_Empty\, Y => \N_19_i\);
    
    full_r : SLE
      port map(D => fulli, CLK => m2s010_som_sb_0_CCC_71MHz, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \TX_FIFO_Full\);
    
    \rptr_bin_sync2[3]\ : SLE
      port map(D => \rptr_bin_sync[3]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[3]_net_1\);
    
    \wptr_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \wptr[0]_net_1\, Y => \wptr_s[0]\);
    
    \rptr[2]\ : SLE
      port map(D => \rptr_s[2]\, CLK => BIT_CLK, EN => \N_19_i\, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[2]_net_1\);
    
    \memraddr_r[3]\ : SLE
      port map(D => \memraddr_r_s[3]\, CLK => BIT_CLK, EN => 
        \N_19_i\, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[3]\);
    
    \rptr_bin_sync2[9]\ : SLE
      port map(D => \rptr_bin_sync[9]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[9]_net_1\);
    
    \L1.empty_r_3_0_a3_2\ : CFG2
      generic map(INIT => x"1")

      port map(A => \rdiff_bus[6]\, B => \rdiff_bus[5]\, Y => 
        empty_r_3_0_a3_2);
    
    \rptr[11]\ : SLE
      port map(D => \rptr_s[11]_net_1\, CLK => BIT_CLK, EN => 
        \N_19_i\, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rptr[11]_net_1\);
    
    \wptr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[5]_net_1\, S
         => \wptr_s[6]\, Y => OPEN, FCO => \wptr_cry[6]_net_1\);
    
    \rptr_bin_sync2[11]\ : SLE
      port map(D => \rptr_bin_sync[11]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[11]_net_1\);
    
    \wptr_bin_sync2[5]\ : SLE
      port map(D => \wptr_bin_sync[5]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[5]_net_1\);
    
    \wptr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[7]_net_1\, S
         => \wptr_s[8]\, Y => OPEN, FCO => \wptr_cry[8]_net_1\);
    
    \wptr_bin_sync2[1]\ : SLE
      port map(D => \wptr_bin_sync[1]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[1]_net_1\);
    
    Wr_corefifo_grayToBinConv : 
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv_0
      port map(wptr_bin_sync(11) => \wptr_bin_sync[11]\, 
        wptr_bin_sync(10) => \wptr_bin_sync[10]\, 
        wptr_bin_sync(9) => \wptr_bin_sync[9]\, wptr_bin_sync(8)
         => \wptr_bin_sync[8]\, wptr_bin_sync(7) => 
        \wptr_bin_sync[7]\, wptr_bin_sync(6) => 
        \wptr_bin_sync[6]\, wptr_bin_sync(5) => 
        \wptr_bin_sync[5]\, wptr_bin_sync(4) => 
        \wptr_bin_sync[4]\, wptr_bin_sync(3) => nc1, 
        wptr_bin_sync(2) => \wptr_bin_sync[2]\, wptr_bin_sync(1)
         => \wptr_bin_sync[1]\, wptr_bin_sync(0) => 
        \wptr_bin_sync[0]\, wptr_gray_sync(10) => 
        \wptr_gray_sync[10]\, wptr_gray_sync(9) => 
        \wptr_gray_sync[9]\, wptr_gray_sync(8) => 
        \wptr_gray_sync[8]\, wptr_gray_sync(7) => 
        \wptr_gray_sync[7]\, wptr_gray_sync(6) => 
        \wptr_gray_sync[6]\, wptr_gray_sync(5) => 
        \wptr_gray_sync[5]\, wptr_gray_sync(4) => 
        \wptr_gray_sync[4]\, wptr_gray_sync(3) => 
        \wptr_gray_sync[3]\, wptr_gray_sync(2) => 
        \wptr_gray_sync[2]\, wptr_gray_sync(1) => 
        \wptr_gray_sync[1]\, wptr_gray_sync(0) => 
        \wptr_gray_sync[0]\, bin_N_4_0_i => bin_N_4_0_i);
    
    \wptr_gray_1[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[4]_net_1\, B => \wptr[5]_net_1\, Y => 
        \wptr_gray_1[4]_net_1\);
    
    overflow_r : SLE
      port map(D => N_7_i, CLK => m2s010_som_sb_0_CCC_71MHz, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \TX_FIFO_OVERFLOW\);
    
    fulli_0 : CFG4
      generic map(INIT => x"ECCC")

      port map(A => \fulli_0_a3_7\, B => \wdiff_bus[11]\, C => 
        \fulli_0_a3_8\, D => \fulli_0_a3_6\, Y => fulli);
    
    \memraddr_r_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \fifo_MEMRADDR[0]\, Y => \memraddr_r_s[0]\);
    
    \rptr_gray[11]\ : SLE
      port map(D => \rptr[11]_net_1\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[11]_net_1\);
    
    \wptr_bin_sync2[10]\ : SLE
      port map(D => \wptr_bin_sync[10]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[10]_net_1\);
    
    \rptr[10]\ : SLE
      port map(D => \rptr_s[10]\, CLK => BIT_CLK, EN => \N_19_i\, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[10]_net_1\);
    
    \wptr[9]\ : SLE
      port map(D => \wptr_s[9]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[9]_net_1\);
    
    Wr_corefifo_doubleSync : 
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_1
      port map(wptr_gray(11) => \wptr_gray[11]_net_1\, 
        wptr_gray(10) => \wptr_gray[10]_net_1\, wptr_gray(9) => 
        \wptr_gray[9]_net_1\, wptr_gray(8) => 
        \wptr_gray[8]_net_1\, wptr_gray(7) => 
        \wptr_gray[7]_net_1\, wptr_gray(6) => 
        \wptr_gray[6]_net_1\, wptr_gray(5) => 
        \wptr_gray[5]_net_1\, wptr_gray(4) => 
        \wptr_gray[4]_net_1\, wptr_gray(3) => 
        \wptr_gray[3]_net_1\, wptr_gray(2) => 
        \wptr_gray[2]_net_1\, wptr_gray(1) => 
        \wptr_gray[1]_net_1\, wptr_gray(0) => 
        \wptr_gray[0]_net_1\, wptr_gray_sync(10) => 
        \wptr_gray_sync[10]\, wptr_gray_sync(9) => 
        \wptr_gray_sync[9]\, wptr_gray_sync(8) => 
        \wptr_gray_sync[8]\, wptr_gray_sync(7) => 
        \wptr_gray_sync[7]\, wptr_gray_sync(6) => 
        \wptr_gray_sync[6]\, wptr_gray_sync(5) => 
        \wptr_gray_sync[5]\, wptr_gray_sync(4) => 
        \wptr_gray_sync[4]\, wptr_gray_sync(3) => 
        \wptr_gray_sync[3]\, wptr_gray_sync(2) => 
        \wptr_gray_sync[2]\, wptr_gray_sync(1) => 
        \wptr_gray_sync[1]\, wptr_gray_sync(0) => 
        \wptr_gray_sync[0]\, wptr_bin_sync_0 => 
        \wptr_bin_sync[11]\, BIT_CLK => BIT_CLK, itx_fifo_rst_i
         => itx_fifo_rst_i);
    
    \rptr_gray[0]\ : SLE
      port map(D => \rptr_gray_1[0]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[0]_net_1\);
    
    empty_r : SLE
      port map(D => empty_r_3, CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => GND_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \TX_FIFO_Empty\);
    
    \memwaddr_r_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \fifo_MEMWADDR[0]\, Y => \memwaddr_r_s[0]\);
    
    \rptr_gray_1[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[7]_net_1\, B => \rptr[8]_net_1\, Y => 
        \rptr_gray_1[7]_net_1\);
    
    \wptr[4]\ : SLE
      port map(D => \wptr_s[4]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[4]_net_1\);
    
    \memwaddr_r[8]\ : SLE
      port map(D => \memwaddr_r_s[8]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[8]\);
    
    \memwaddr_r[2]\ : SLE
      port map(D => \memwaddr_r_s[2]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[2]\);
    
    \wptr_bin_sync2[11]\ : SLE
      port map(D => \wptr_bin_sync[11]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[11]_net_1\);
    
    memwaddr_r_s_911 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[0]\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => memwaddr_r_s_911_FCO);
    
    \wptr_gray_1[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[1]_net_1\, B => \wptr[2]_net_1\, Y => 
        \wptr_gray_1[1]_net_1\);
    
    underflow_r : SLE
      port map(D => N_12_i, CLK => BIT_CLK, EN => VCC_net_1, ALn
         => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \TX_FIFO_UNDERRUN\);
    
    fulli_0_a3_7 : CFG4
      generic map(INIT => x"8000")

      port map(A => \wdiff_bus[2]\, B => \wdiff_bus[3]\, C => 
        \wdiff_bus[5]\, D => \wdiff_bus[4]\, Y => \fulli_0_a3_7\);
    
    \memwaddr_r_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[6]_net_1\, S => \memwaddr_r_s[7]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[7]_net_1\);
    
    \wptr_gray[5]\ : SLE
      port map(D => \wptr_gray_1[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[5]_net_1\);
    
    overflow_r_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => \TX_FIFO_Full\, B => TX_FIFO_wr_en, Y => 
        N_7_i);
    
    \memraddr_r[7]\ : SLE
      port map(D => \memraddr_r_s[7]\, CLK => BIT_CLK, EN => 
        \N_19_i\, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[7]\);
    
    \rptr_bin_sync2[10]\ : SLE
      port map(D => \rptr_bin_sync[10]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[10]_net_1\);
    
    wdiff_bus_cry_10 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[10]_net_1\, B => 
        \rptr_bin_sync2[10]_net_1\, C => GND_net_1, D => 
        GND_net_1, FCI => \wdiff_bus_cry_9\, S => \wdiff_bus[10]\, 
        Y => OPEN, FCO => \wdiff_bus_cry_10\);
    
    \memwaddr_r_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[9]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[8]_net_1\, S => \memwaddr_r_s[9]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[9]_net_1\);
    
    \wptr_gray[8]\ : SLE
      port map(D => \wptr_gray_1[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[8]_net_1\);
    
    \wptr_gray[7]\ : SLE
      port map(D => \wptr_gray_1[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[7]_net_1\);
    
    \wptr_gray_1[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[5]_net_1\, B => \wptr[6]_net_1\, Y => 
        \wptr_gray_1[5]_net_1\);
    
    \memwaddr_r[5]\ : SLE
      port map(D => \memwaddr_r_s[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[5]\);
    
    \rptr[8]\ : SLE
      port map(D => \rptr_s[8]\, CLK => BIT_CLK, EN => \N_19_i\, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[8]_net_1\);
    
    Rd_corefifo_doubleSync : 
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_doubleSync_0
      port map(rptr_gray(11) => \rptr_gray[11]_net_1\, 
        rptr_gray(10) => \rptr_gray[10]_net_1\, rptr_gray(9) => 
        \rptr_gray[9]_net_1\, rptr_gray(8) => 
        \rptr_gray[8]_net_1\, rptr_gray(7) => 
        \rptr_gray[7]_net_1\, rptr_gray(6) => 
        \rptr_gray[6]_net_1\, rptr_gray(5) => 
        \rptr_gray[5]_net_1\, rptr_gray(4) => 
        \rptr_gray[4]_net_1\, rptr_gray(3) => 
        \rptr_gray[3]_net_1\, rptr_gray(2) => 
        \rptr_gray[2]_net_1\, rptr_gray(1) => 
        \rptr_gray[1]_net_1\, rptr_gray(0) => 
        \rptr_gray[0]_net_1\, rptr_gray_sync(10) => 
        \rptr_gray_sync[10]\, rptr_gray_sync(9) => 
        \rptr_gray_sync[9]\, rptr_gray_sync(8) => 
        \rptr_gray_sync[8]\, rptr_gray_sync(7) => 
        \rptr_gray_sync[7]\, rptr_gray_sync(6) => 
        \rptr_gray_sync[6]\, rptr_gray_sync(5) => 
        \rptr_gray_sync[5]\, rptr_gray_sync(4) => 
        \rptr_gray_sync[4]\, rptr_gray_sync(3) => 
        \rptr_gray_sync[3]\, rptr_gray_sync(2) => 
        \rptr_gray_sync[2]\, rptr_gray_sync(1) => 
        \rptr_gray_sync[1]\, rptr_gray_sync(0) => 
        \rptr_gray_sync[0]\, rptr_bin_sync_0 => 
        \rptr_bin_sync[11]\, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, itx_fifo_rst_i => 
        itx_fifo_rst_i);
    
    underflow_r_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => N_114, B => \TX_FIFO_Empty\, Y => N_12_i);
    
    \rptr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[3]_net_1\, S
         => \rptr_s[4]\, Y => OPEN, FCO => \rptr_cry[4]_net_1\);
    
    wdiff_bus_cry_2 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[2]_net_1\, B => 
        \rptr_bin_sync2[2]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_1\, S => \wdiff_bus[2]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_2\);
    
    \rptr_gray[2]\ : SLE
      port map(D => \rptr_gray_1[2]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[2]_net_1\);
    
    \wptr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[8]_net_1\, S
         => \wptr_s[9]\, Y => OPEN, FCO => \wptr_cry[9]_net_1\);
    
    \wptr_bin_sync2[3]\ : SLE
      port map(D => bin_N_4_0_i, CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[3]_net_1\);
    
    \wptr[2]\ : SLE
      port map(D => \wptr_s[2]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[2]_net_1\);
    
    \rptr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[1]_net_1\, S
         => \rptr_s[2]\, Y => OPEN, FCO => \rptr_cry[2]_net_1\);
    
    rdiff_bus_cry_9 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[9]_net_1\, B => 
        \rptr[9]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_8\, S => \rdiff_bus[9]\, Y => OPEN, FCO
         => \rdiff_bus_cry_9\);
    
    \memwaddr_r[0]\ : SLE
      port map(D => \memwaddr_r_s[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[0]\);
    
    \wptr_gray[2]\ : SLE
      port map(D => \wptr_gray_1[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[2]_net_1\);
    
    wdiff_bus_cry_4 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[4]_net_1\, B => 
        \rptr_bin_sync2[4]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_3\, S => \wdiff_bus[4]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_4\);
    
    \memwaddr_r_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[2]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[1]_net_1\, S => \memwaddr_r_s[2]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[2]_net_1\);
    
    \wptr_gray[11]\ : SLE
      port map(D => \wptr[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[11]_net_1\);
    
    \wptr_bin_sync2[9]\ : SLE
      port map(D => \wptr_bin_sync[9]\, CLK => BIT_CLK, EN => 
        VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[9]_net_1\);
    
    \rptr_gray_1[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[6]_net_1\, B => \rptr[7]_net_1\, Y => 
        \rptr_gray_1[6]_net_1\);
    
    \wptr_gray_1[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[11]_net_1\, B => \wptr[10]_net_1\, Y
         => \wptr_gray_1[10]_net_1\);
    
    wdiff_bus_cry_6 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[6]_net_1\, B => 
        \rptr_bin_sync2[6]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_5\, S => \wdiff_bus[6]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_6\);
    
    \rptr_s[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[10]_net_1\, S
         => \rptr_s[11]_net_1\, Y => OPEN, FCO => OPEN);
    
    \rptr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[2]_net_1\, S
         => \rptr_s[3]\, Y => OPEN, FCO => \rptr_cry[3]_net_1\);
    
    \memraddr_r[4]\ : SLE
      port map(D => \memraddr_r_s[4]\, CLK => BIT_CLK, EN => 
        \N_19_i\, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[4]\);
    
    \memraddr_r_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[6]_net_1\, S => \memraddr_r_s[7]\, Y => 
        OPEN, FCO => \memraddr_r_cry[7]_net_1\);
    
    \L1.empty_r_3_0_a3_5\ : CFG3
      generic map(INIT => x"01")

      port map(A => \rdiff_bus[1]\, B => \rdiff_bus[11]\, C => 
        \rdiff_bus[2]\, Y => empty_r_3_0_a3_5);
    
    \memraddr_r_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[9]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[8]_net_1\, S => \memraddr_r_s[9]\, Y => 
        OPEN, FCO => \memraddr_r_cry[9]_net_1\);
    
    \memraddr_r[5]\ : SLE
      port map(D => \memraddr_r_s[5]\, CLK => BIT_CLK, EN => 
        \N_19_i\, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[5]\);
    
    \rptr_gray[6]\ : SLE
      port map(D => \rptr_gray_1[6]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[6]_net_1\);
    
    \memraddr_r[9]\ : SLE
      port map(D => \memraddr_r_s[9]\, CLK => BIT_CLK, EN => 
        \N_19_i\, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[9]\);
    
    \rptr[0]\ : SLE
      port map(D => \rptr_s[0]\, CLK => BIT_CLK, EN => \N_19_i\, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \rptr[0]_net_1\);
    
    fulli_0_a3_6 : CFG4
      generic map(INIT => x"4000")

      port map(A => wdiff_bus_cry_0_Y, B => TX_FIFO_wr_en, C => 
        \wdiff_bus[10]\, D => \wdiff_bus[1]\, Y => \fulli_0_a3_6\);
    
    \wptr[10]\ : SLE
      port map(D => \wptr_s[10]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMWE\, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \wptr[10]_net_1\);
    
    \memwaddr_r_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memwaddr_r_cry[3]_net_1\, S => \memwaddr_r_s[4]\, Y => 
        OPEN, FCO => \memwaddr_r_cry[4]_net_1\);
    
    \memraddr_r_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[3]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[2]_net_1\, S => \memraddr_r_s[3]\, Y => 
        OPEN, FCO => \memraddr_r_cry[3]_net_1\);
    
    wdiff_bus_cry_1 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[1]_net_1\, B => 
        \rptr_bin_sync2[1]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_0\, S => \wdiff_bus[1]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_1\);
    
    rdiff_bus_cry_2 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[2]_net_1\, B => 
        \rptr[2]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_1\, S => \rdiff_bus[2]\, Y => OPEN, FCO
         => \rdiff_bus_cry_2\);
    
    \wptr_gray[9]\ : SLE
      port map(D => \wptr_gray_1[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[9]_net_1\);
    
    \rptr_gray_1[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[4]_net_1\, B => \rptr[5]_net_1\, Y => 
        \rptr_gray_1[4]_net_1\);
    
    \wptr_gray_1[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[8]_net_1\, B => \wptr[9]_net_1\, Y => 
        \wptr_gray_1[8]_net_1\);
    
    Rd_corefifo_grayToBinConv : 
        FIFO_2Kx8_FIFO_2Kx8_0_corefifo_grayToBinConv
      port map(rptr_bin_sync(11) => \rptr_bin_sync[11]\, 
        rptr_bin_sync(10) => \rptr_bin_sync[10]\, 
        rptr_bin_sync(9) => \rptr_bin_sync[9]\, rptr_bin_sync(8)
         => \rptr_bin_sync[8]\, rptr_bin_sync(7) => 
        \rptr_bin_sync[7]\, rptr_bin_sync(6) => 
        \rptr_bin_sync[6]\, rptr_bin_sync(5) => 
        \rptr_bin_sync[5]\, rptr_bin_sync(4) => 
        \rptr_bin_sync[4]\, rptr_bin_sync(3) => 
        \rptr_bin_sync[3]\, rptr_bin_sync(2) => 
        \rptr_bin_sync[2]\, rptr_bin_sync(1) => 
        \rptr_bin_sync[1]\, rptr_bin_sync(0) => 
        \rptr_bin_sync[0]\, rptr_gray_sync(10) => 
        \rptr_gray_sync[10]\, rptr_gray_sync(9) => 
        \rptr_gray_sync[9]\, rptr_gray_sync(8) => 
        \rptr_gray_sync[8]\, rptr_gray_sync(7) => 
        \rptr_gray_sync[7]\, rptr_gray_sync(6) => 
        \rptr_gray_sync[6]\, rptr_gray_sync(5) => 
        \rptr_gray_sync[5]\, rptr_gray_sync(4) => 
        \rptr_gray_sync[4]\, rptr_gray_sync(3) => 
        \rptr_gray_sync[3]\, rptr_gray_sync(2) => 
        \rptr_gray_sync[2]\, rptr_gray_sync(1) => 
        \rptr_gray_sync[1]\, rptr_gray_sync(0) => 
        \rptr_gray_sync[0]\);
    
    \rptr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => rptr_s_913_FCO, S => 
        \rptr_s[1]\, Y => OPEN, FCO => \rptr_cry[1]_net_1\);
    
    rdiff_bus_cry_3 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[3]_net_1\, B => 
        \rptr[3]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_2\, S => \rdiff_bus[3]\, Y => OPEN, FCO
         => \rdiff_bus_cry_3\);
    
    rdiff_bus_cry_10 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[10]_net_1\, B => 
        \rptr[10]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_9\, S => \rdiff_bus[10]\, Y => OPEN, FCO
         => \rdiff_bus_cry_10\);
    
    \memraddr_r_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        \memraddr_r_cry[5]_net_1\, S => \memraddr_r_s[6]\, Y => 
        OPEN, FCO => \memraddr_r_cry[6]_net_1\);
    
    \memraddr_r[6]\ : SLE
      port map(D => \memraddr_r_s[6]\, CLK => BIT_CLK, EN => 
        \N_19_i\, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[6]\);
    
    \rptr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[6]_net_1\, S
         => \rptr_s[7]\, Y => OPEN, FCO => \rptr_cry[7]_net_1\);
    
    rdiff_bus_cry_0 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => rdiff_bus, B => \rptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => rdiff_bus_cry_0_Y, FCO => \rdiff_bus_cry_0\);
    
    \memraddr_r[2]\ : SLE
      port map(D => \memraddr_r_s[2]\, CLK => BIT_CLK, EN => 
        \N_19_i\, ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \fifo_MEMRADDR[2]\);
    
    \wptr[8]\ : SLE
      port map(D => \wptr_s[8]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMWE\, ALn => itx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \wptr[8]_net_1\);
    
    wdiff_bus_cry_3 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[3]_net_1\, B => 
        \rptr_bin_sync2[3]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_2\, S => \wdiff_bus[3]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_3\);
    
    fulli_0_a3_8 : CFG4
      generic map(INIT => x"8000")

      port map(A => \wdiff_bus[6]\, B => \wdiff_bus[7]\, C => 
        \wdiff_bus[8]\, D => \wdiff_bus[9]\, Y => \fulli_0_a3_8\);
    
    \rptr_gray[7]\ : SLE
      port map(D => \rptr_gray_1[7]_net_1\, CLK => BIT_CLK, EN
         => VCC_net_1, ALn => itx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_gray[7]_net_1\);
    
    \wptr_gray[0]\ : SLE
      port map(D => \wptr_gray_1[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[0]_net_1\);
    
    \rptr_gray_1[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[0]_net_1\, B => \rptr[1]_net_1\, Y => 
        \rptr_gray_1[0]_net_1\);
    
    \rptr_gray_1[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[8]_net_1\, B => \rptr[9]_net_1\, Y => 
        \rptr_gray_1[8]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_2Kx8_FIFO_2Kx8_0_COREFIFO is

    port( CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0);
          TX_FIFO_DOUT                 : out   std_logic_vector(7 downto 0);
          TX_FIFO_UNDERRUN             : out   std_logic;
          TX_FIFO_UNDERRUN_i           : out   std_logic;
          TX_FIFO_OVERFLOW             : out   std_logic;
          TX_FIFO_OVERFLOW_i           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic;
          TX_FIFO_Full                 : out   std_logic;
          TX_FIFO_wr_en                : in    std_logic;
          TX_FIFO_Empty                : out   std_logic;
          N_114                        : in    std_logic;
          BIT_CLK                      : in    std_logic;
          itx_fifo_rst_i               : in    std_logic
        );

end FIFO_2Kx8_FIFO_2Kx8_0_COREFIFO;

architecture DEF_ARCH of FIFO_2Kx8_FIFO_2Kx8_0_COREFIFO is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component FIFO_2Kx8_FIFO_2Kx8_0_ram_wrapper
    port( RDATA_int                    : out   std_logic_vector(7 downto 0);
          fifo_MEMRADDR                : in    std_logic_vector(10 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0) := (others => 'U');
          fifo_MEMWADDR                : in    std_logic_vector(10 downto 0) := (others => 'U');
          BIT_CLK                      : in    std_logic := 'U';
          N_19_i                       : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic := 'U';
          fifo_MEMWE                   : in    std_logic := 'U'
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component FIFO_2Kx8_FIFO_2Kx8_0_corefifo_async
    port( fifo_MEMWADDR             : out   std_logic_vector(10 downto 0);
          fifo_MEMRADDR             : out   std_logic_vector(10 downto 0);
          N_114                     : in    std_logic := 'U';
          TX_FIFO_wr_en             : in    std_logic := 'U';
          fifo_MEMWE                : out   std_logic;
          N_19_i                    : out   std_logic;
          TX_FIFO_Full              : out   std_logic;
          TX_FIFO_Empty             : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          BIT_CLK                   : in    std_logic := 'U';
          itx_fifo_rst_i            : in    std_logic := 'U';
          TX_FIFO_OVERFLOW_i        : out   std_logic;
          TX_FIFO_OVERFLOW          : out   std_logic;
          TX_FIFO_UNDERRUN_i        : out   std_logic;
          TX_FIFO_UNDERRUN          : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \RDATA_r[5]_net_1\, VCC_net_1, \RDATA_int[5]\, N_8_i, 
        GND_net_1, \RDATA_r[6]_net_1\, \RDATA_int[6]\, 
        \RDATA_r[7]_net_1\, \RDATA_int[7]\, \re_set\, \REN_d1\, 
        N_24_i_i, \RDATA_r[0]_net_1\, \RDATA_int[0]\, 
        \RDATA_r[1]_net_1\, \RDATA_int[1]\, \RDATA_r[2]_net_1\, 
        \RDATA_int[2]\, \RDATA_r[3]_net_1\, \RDATA_int[3]\, 
        \RDATA_r[4]_net_1\, \RDATA_int[4]\, N_19_i, \RE_d1\, 
        \re_pulse_d1\, \re_pulse\, \TX_FIFO_Empty\, 
        \fifo_MEMWADDR[0]\, \fifo_MEMWADDR[1]\, 
        \fifo_MEMWADDR[2]\, \fifo_MEMWADDR[3]\, 
        \fifo_MEMWADDR[4]\, \fifo_MEMWADDR[5]\, 
        \fifo_MEMWADDR[6]\, \fifo_MEMWADDR[7]\, 
        \fifo_MEMWADDR[8]\, \fifo_MEMWADDR[9]\, 
        \fifo_MEMWADDR[10]\, \fifo_MEMRADDR[0]\, 
        \fifo_MEMRADDR[1]\, \fifo_MEMRADDR[2]\, 
        \fifo_MEMRADDR[3]\, \fifo_MEMRADDR[4]\, 
        \fifo_MEMRADDR[5]\, \fifo_MEMRADDR[6]\, 
        \fifo_MEMRADDR[7]\, \fifo_MEMRADDR[8]\, 
        \fifo_MEMRADDR[9]\, \fifo_MEMRADDR[10]\, fifo_MEMWE
         : std_logic;

    for all : FIFO_2Kx8_FIFO_2Kx8_0_ram_wrapper
	Use entity work.FIFO_2Kx8_FIFO_2Kx8_0_ram_wrapper(DEF_ARCH);
    for all : FIFO_2Kx8_FIFO_2Kx8_0_corefifo_async
	Use entity work.FIFO_2Kx8_FIFO_2Kx8_0_corefifo_async(DEF_ARCH);
begin 

    TX_FIFO_Empty <= \TX_FIFO_Empty\;

    re_pulse : CFG4
      generic map(INIT => x"EAEE")

      port map(A => \re_set\, B => \REN_d1\, C => \TX_FIFO_Empty\, 
        D => N_114, Y => \re_pulse\);
    
    \RDATA_r[3]\ : SLE
      port map(D => \RDATA_int[3]\, CLK => BIT_CLK, EN => N_8_i, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[3]_net_1\);
    
    \Q[6]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[6]_net_1\, C => 
        \RDATA_int[6]\, D => \RE_d1\, Y => TX_FIFO_DOUT(6));
    
    re_pulse_d1 : SLE
      port map(D => \re_pulse\, CLK => BIT_CLK, EN => VCC_net_1, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \re_pulse_d1\);
    
    \RDATA_r[5]\ : SLE
      port map(D => \RDATA_int[5]\, CLK => BIT_CLK, EN => N_8_i, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[5]_net_1\);
    
    \Q[2]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[2]_net_1\, C => 
        \RDATA_int[2]\, D => \RE_d1\, Y => TX_FIFO_DOUT(2));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \RW1.UI_ram_wrapper_1\ : FIFO_2Kx8_FIFO_2Kx8_0_ram_wrapper
      port map(RDATA_int(7) => \RDATA_int[7]\, RDATA_int(6) => 
        \RDATA_int[6]\, RDATA_int(5) => \RDATA_int[5]\, 
        RDATA_int(4) => \RDATA_int[4]\, RDATA_int(3) => 
        \RDATA_int[3]\, RDATA_int(2) => \RDATA_int[2]\, 
        RDATA_int(1) => \RDATA_int[1]\, RDATA_int(0) => 
        \RDATA_int[0]\, fifo_MEMRADDR(10) => \fifo_MEMRADDR[10]\, 
        fifo_MEMRADDR(9) => \fifo_MEMRADDR[9]\, fifo_MEMRADDR(8)
         => \fifo_MEMRADDR[8]\, fifo_MEMRADDR(7) => 
        \fifo_MEMRADDR[7]\, fifo_MEMRADDR(6) => 
        \fifo_MEMRADDR[6]\, fifo_MEMRADDR(5) => 
        \fifo_MEMRADDR[5]\, fifo_MEMRADDR(4) => 
        \fifo_MEMRADDR[4]\, fifo_MEMRADDR(3) => 
        \fifo_MEMRADDR[3]\, fifo_MEMRADDR(2) => 
        \fifo_MEMRADDR[2]\, fifo_MEMRADDR(1) => 
        \fifo_MEMRADDR[1]\, fifo_MEMRADDR(0) => 
        \fifo_MEMRADDR[0]\, CoreAPB3_0_APBmslave0_PWDATA(7) => 
        CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), fifo_MEMWADDR(10) => 
        \fifo_MEMWADDR[10]\, fifo_MEMWADDR(9) => 
        \fifo_MEMWADDR[9]\, fifo_MEMWADDR(8) => 
        \fifo_MEMWADDR[8]\, fifo_MEMWADDR(7) => 
        \fifo_MEMWADDR[7]\, fifo_MEMWADDR(6) => 
        \fifo_MEMWADDR[6]\, fifo_MEMWADDR(5) => 
        \fifo_MEMWADDR[5]\, fifo_MEMWADDR(4) => 
        \fifo_MEMWADDR[4]\, fifo_MEMWADDR(3) => 
        \fifo_MEMWADDR[3]\, fifo_MEMWADDR(2) => 
        \fifo_MEMWADDR[2]\, fifo_MEMWADDR(1) => 
        \fifo_MEMWADDR[1]\, fifo_MEMWADDR(0) => 
        \fifo_MEMWADDR[0]\, BIT_CLK => BIT_CLK, N_19_i => N_19_i, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz, 
        fifo_MEMWE => fifo_MEMWE);
    
    \RDATA_r[0]\ : SLE
      port map(D => \RDATA_int[0]\, CLK => BIT_CLK, EN => N_8_i, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[0]_net_1\);
    
    \Q[4]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[4]_net_1\, C => 
        \RDATA_int[4]\, D => \RE_d1\, Y => TX_FIFO_DOUT(4));
    
    \RDATA_r[2]\ : SLE
      port map(D => \RDATA_int[2]\, CLK => BIT_CLK, EN => N_8_i, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[2]_net_1\);
    
    \RDATA_r[6]\ : SLE
      port map(D => \RDATA_int[6]\, CLK => BIT_CLK, EN => N_8_i, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[6]_net_1\);
    
    REN_d1_RNISQRI : CFG3
      generic map(INIT => x"C4")

      port map(A => N_114, B => \REN_d1\, C => \TX_FIFO_Empty\, Y
         => N_8_i);
    
    \L31.U_corefifo_async\ : FIFO_2Kx8_FIFO_2Kx8_0_corefifo_async
      port map(fifo_MEMWADDR(10) => \fifo_MEMWADDR[10]\, 
        fifo_MEMWADDR(9) => \fifo_MEMWADDR[9]\, fifo_MEMWADDR(8)
         => \fifo_MEMWADDR[8]\, fifo_MEMWADDR(7) => 
        \fifo_MEMWADDR[7]\, fifo_MEMWADDR(6) => 
        \fifo_MEMWADDR[6]\, fifo_MEMWADDR(5) => 
        \fifo_MEMWADDR[5]\, fifo_MEMWADDR(4) => 
        \fifo_MEMWADDR[4]\, fifo_MEMWADDR(3) => 
        \fifo_MEMWADDR[3]\, fifo_MEMWADDR(2) => 
        \fifo_MEMWADDR[2]\, fifo_MEMWADDR(1) => 
        \fifo_MEMWADDR[1]\, fifo_MEMWADDR(0) => 
        \fifo_MEMWADDR[0]\, fifo_MEMRADDR(10) => 
        \fifo_MEMRADDR[10]\, fifo_MEMRADDR(9) => 
        \fifo_MEMRADDR[9]\, fifo_MEMRADDR(8) => 
        \fifo_MEMRADDR[8]\, fifo_MEMRADDR(7) => 
        \fifo_MEMRADDR[7]\, fifo_MEMRADDR(6) => 
        \fifo_MEMRADDR[6]\, fifo_MEMRADDR(5) => 
        \fifo_MEMRADDR[5]\, fifo_MEMRADDR(4) => 
        \fifo_MEMRADDR[4]\, fifo_MEMRADDR(3) => 
        \fifo_MEMRADDR[3]\, fifo_MEMRADDR(2) => 
        \fifo_MEMRADDR[2]\, fifo_MEMRADDR(1) => 
        \fifo_MEMRADDR[1]\, fifo_MEMRADDR(0) => 
        \fifo_MEMRADDR[0]\, N_114 => N_114, TX_FIFO_wr_en => 
        TX_FIFO_wr_en, fifo_MEMWE => fifo_MEMWE, N_19_i => N_19_i, 
        TX_FIFO_Full => TX_FIFO_Full, TX_FIFO_Empty => 
        \TX_FIFO_Empty\, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, BIT_CLK => BIT_CLK, 
        itx_fifo_rst_i => itx_fifo_rst_i, TX_FIFO_OVERFLOW_i => 
        TX_FIFO_OVERFLOW_i, TX_FIFO_OVERFLOW => TX_FIFO_OVERFLOW, 
        TX_FIFO_UNDERRUN_i => TX_FIFO_UNDERRUN_i, 
        TX_FIFO_UNDERRUN => TX_FIFO_UNDERRUN);
    
    re_set : SLE
      port map(D => \REN_d1\, CLK => BIT_CLK, EN => N_24_i_i, ALn
         => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \re_set\);
    
    \Q[3]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[3]_net_1\, C => 
        \RDATA_int[3]\, D => \RE_d1\, Y => TX_FIFO_DOUT(3));
    
    \Q[7]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[7]_net_1\, C => 
        \RDATA_int[7]\, D => \RE_d1\, Y => TX_FIFO_DOUT(7));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    RE_d1 : SLE
      port map(D => N_114, CLK => BIT_CLK, EN => VCC_net_1, ALn
         => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \RE_d1\);
    
    \RDATA_r[7]\ : SLE
      port map(D => \RDATA_int[7]\, CLK => BIT_CLK, EN => N_8_i, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[7]_net_1\);
    
    \RDATA_r[4]\ : SLE
      port map(D => \RDATA_int[4]\, CLK => BIT_CLK, EN => N_8_i, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[4]_net_1\);
    
    \Q[1]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[1]_net_1\, C => 
        \RDATA_int[1]\, D => \RE_d1\, Y => TX_FIFO_DOUT(1));
    
    \Q[0]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[0]_net_1\, C => 
        \RDATA_int[0]\, D => \RE_d1\, Y => TX_FIFO_DOUT(0));
    
    REN_d1 : SLE
      port map(D => N_19_i, CLK => BIT_CLK, EN => VCC_net_1, ALn
         => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => \REN_d1\);
    
    \Q[5]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[5]_net_1\, C => 
        \RDATA_int[5]\, D => \RE_d1\, Y => TX_FIFO_DOUT(5));
    
    re_set_RNO : CFG3
      generic map(INIT => x"C6")

      port map(A => N_114, B => \REN_d1\, C => \TX_FIFO_Empty\, Y
         => N_24_i_i);
    
    \RDATA_r[1]\ : SLE
      port map(D => \RDATA_int[1]\, CLK => BIT_CLK, EN => N_8_i, 
        ALn => itx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[1]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_2Kx8 is

    port( TX_FIFO_DOUT                 : out   std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0);
          itx_fifo_rst_i               : in    std_logic;
          BIT_CLK                      : in    std_logic;
          N_114                        : in    std_logic;
          TX_FIFO_Empty                : out   std_logic;
          TX_FIFO_wr_en                : in    std_logic;
          TX_FIFO_Full                 : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic;
          TX_FIFO_OVERFLOW_i           : out   std_logic;
          TX_FIFO_OVERFLOW             : out   std_logic;
          TX_FIFO_UNDERRUN_i           : out   std_logic;
          TX_FIFO_UNDERRUN             : out   std_logic
        );

end FIFO_2Kx8;

architecture DEF_ARCH of FIFO_2Kx8 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component FIFO_2Kx8_FIFO_2Kx8_0_COREFIFO
    port( CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0) := (others => 'U');
          TX_FIFO_DOUT                 : out   std_logic_vector(7 downto 0);
          TX_FIFO_UNDERRUN             : out   std_logic;
          TX_FIFO_UNDERRUN_i           : out   std_logic;
          TX_FIFO_OVERFLOW             : out   std_logic;
          TX_FIFO_OVERFLOW_i           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic := 'U';
          TX_FIFO_Full                 : out   std_logic;
          TX_FIFO_wr_en                : in    std_logic := 'U';
          TX_FIFO_Empty                : out   std_logic;
          N_114                        : in    std_logic := 'U';
          BIT_CLK                      : in    std_logic := 'U';
          itx_fifo_rst_i               : in    std_logic := 'U'
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : FIFO_2Kx8_FIFO_2Kx8_0_COREFIFO
	Use entity work.FIFO_2Kx8_FIFO_2Kx8_0_COREFIFO(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    FIFO_2Kx8_0 : FIFO_2Kx8_FIFO_2Kx8_0_COREFIFO
      port map(CoreAPB3_0_APBmslave0_PWDATA(7) => 
        CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), TX_FIFO_DOUT(7) => 
        TX_FIFO_DOUT(7), TX_FIFO_DOUT(6) => TX_FIFO_DOUT(6), 
        TX_FIFO_DOUT(5) => TX_FIFO_DOUT(5), TX_FIFO_DOUT(4) => 
        TX_FIFO_DOUT(4), TX_FIFO_DOUT(3) => TX_FIFO_DOUT(3), 
        TX_FIFO_DOUT(2) => TX_FIFO_DOUT(2), TX_FIFO_DOUT(1) => 
        TX_FIFO_DOUT(1), TX_FIFO_DOUT(0) => TX_FIFO_DOUT(0), 
        TX_FIFO_UNDERRUN => TX_FIFO_UNDERRUN, TX_FIFO_UNDERRUN_i
         => TX_FIFO_UNDERRUN_i, TX_FIFO_OVERFLOW => 
        TX_FIFO_OVERFLOW, TX_FIFO_OVERFLOW_i => 
        TX_FIFO_OVERFLOW_i, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, TX_FIFO_Full => TX_FIFO_Full, 
        TX_FIFO_wr_en => TX_FIFO_wr_en, TX_FIFO_Empty => 
        TX_FIFO_Empty, N_114 => N_114, BIT_CLK => BIT_CLK, 
        itx_fifo_rst_i => itx_fifo_rst_i);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_0 is

    port( RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          RDATA_int                 : out   std_logic_vector(8 downto 0);
          fifo_MEMWADDR             : in    std_logic_vector(12 downto 0);
          fifo_MEMRADDR             : in    std_logic_vector(12 downto 0);
          fifo_MEMWE                : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          fifo_MEMRE                : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_0;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component RAM1K18
    generic (MEMORYFILE:string := "");

    port( A_DOUT        : out   std_logic_vector(17 downto 0);
          B_DOUT        : out   std_logic_vector(17 downto 0);
          BUSY          : out   std_logic;
          A_CLK         : in    std_logic := 'U';
          A_DOUT_CLK    : in    std_logic := 'U';
          A_ARST_N      : in    std_logic := 'U';
          A_DOUT_EN     : in    std_logic := 'U';
          A_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_DOUT_ARST_N : in    std_logic := 'U';
          A_DOUT_SRST_N : in    std_logic := 'U';
          A_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          A_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          A_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          B_CLK         : in    std_logic := 'U';
          B_DOUT_CLK    : in    std_logic := 'U';
          B_ARST_N      : in    std_logic := 'U';
          B_DOUT_EN     : in    std_logic := 'U';
          B_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_DOUT_ARST_N : in    std_logic := 'U';
          B_DOUT_SRST_N : in    std_logic := 'U';
          B_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          B_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          B_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          A_EN          : in    std_logic := 'U';
          A_DOUT_LAT    : in    std_logic := 'U';
          A_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_WMODE       : in    std_logic := 'U';
          B_EN          : in    std_logic := 'U';
          B_DOUT_LAT    : in    std_logic := 'U';
          B_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_WMODE       : in    std_logic := 'U';
          SII_LOCK      : in    std_logic := 'U'
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;
    signal nc151, nc23, nc58, nc116, nc74, nc133, nc167, nc84, 
        nc39, nc72, nc82, nc145, nc160, nc57, nc156, nc125, nc73, 
        nc107, nc66, nc83, nc9, nc171, nc54, nc135, nc41, nc100, 
        nc52, nc29, nc118, nc60, nc141, nc45, nc53, nc121, nc158, 
        nc162, nc11, nc131, nc96, nc79, nc146, nc89, nc119, nc48, 
        nc126, nc15, nc102, nc3, nc47, nc90, nc159, nc136, nc59, 
        nc18, nc44, nc117, nc164, nc148, nc42, nc17, nc2, nc110, 
        nc128, nc43, nc157, nc36, nc61, nc104, nc138, nc14, nc150, 
        nc149, nc12, nc30, nc65, nc7, nc129, nc8, nc13, nc26, 
        nc139, nc163, nc112, nc68, nc49, nc170, nc91, nc5, nc20, 
        nc147, nc67, nc152, nc127, nc103, nc76, nc140, nc86, nc95, 
        nc120, nc165, nc137, nc64, nc19, nc70, nc62, nc80, nc130, 
        nc98, nc114, nc56, nc105, nc63, nc97, nc161, nc31, nc154, 
        nc50, nc142, nc94, nc122, nc35, nc4, nc92, nc101, nc166, 
        nc132, nc21, nc93, nc69, nc38, nc113, nc106, nc25, nc1, 
        nc37, nc144, nc153, nc46, nc71, nc124, nc81, nc168, nc34, 
        nc28, nc115, nc134, nc32, nc40, nc99, nc75, nc85, nc27, 
        nc108, nc16, nc155, nc51, nc33, nc169, nc78, nc24, nc88, 
        nc111, nc55, nc10, nc22, nc143, nc77, nc6, nc109, nc87, 
        nc123 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C2 : RAM1K18
      port map(A_DOUT(17) => nc151, A_DOUT(16) => nc23, 
        A_DOUT(15) => nc58, A_DOUT(14) => nc116, A_DOUT(13) => 
        nc74, A_DOUT(12) => nc133, A_DOUT(11) => nc167, 
        A_DOUT(10) => nc84, A_DOUT(9) => nc39, A_DOUT(8) => nc72, 
        A_DOUT(7) => nc82, A_DOUT(6) => nc145, A_DOUT(5) => nc160, 
        A_DOUT(4) => nc57, A_DOUT(3) => nc156, A_DOUT(2) => nc125, 
        A_DOUT(1) => RDATA_int(5), A_DOUT(0) => RDATA_int(4), 
        B_DOUT(17) => nc73, B_DOUT(16) => nc107, B_DOUT(15) => 
        nc66, B_DOUT(14) => nc83, B_DOUT(13) => nc9, B_DOUT(12)
         => nc171, B_DOUT(11) => nc54, B_DOUT(10) => nc135, 
        B_DOUT(9) => nc41, B_DOUT(8) => nc100, B_DOUT(7) => nc52, 
        B_DOUT(6) => nc29, B_DOUT(5) => nc118, B_DOUT(4) => nc60, 
        B_DOUT(3) => nc141, B_DOUT(2) => nc45, B_DOUT(1) => nc53, 
        B_DOUT(0) => nc121, BUSY => OPEN, A_CLK => 
        m2s010_som_sb_0_CCC_71MHz, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => fifo_MEMRE, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => fifo_MEMRADDR(12), A_ADDR(12) => fifo_MEMRADDR(11), 
        A_ADDR(11) => fifo_MEMRADDR(10), A_ADDR(10) => 
        fifo_MEMRADDR(9), A_ADDR(9) => fifo_MEMRADDR(8), 
        A_ADDR(8) => fifo_MEMRADDR(7), A_ADDR(7) => 
        fifo_MEMRADDR(6), A_ADDR(6) => fifo_MEMRADDR(5), 
        A_ADDR(5) => fifo_MEMRADDR(4), A_ADDR(4) => 
        fifo_MEMRADDR(3), A_ADDR(3) => fifo_MEMRADDR(2), 
        A_ADDR(2) => fifo_MEMRADDR(1), A_ADDR(1) => 
        fifo_MEMRADDR(0), A_ADDR(0) => GND_net_1, A_WEN(1) => 
        GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => GND_net_1, B_DIN(2) => GND_net_1, B_DIN(1)
         => RX_FIFO_DIN_pipe(5), B_DIN(0) => RX_FIFO_DIN_pipe(4), 
        B_ADDR(13) => fifo_MEMWADDR(12), B_ADDR(12) => 
        fifo_MEMWADDR(11), B_ADDR(11) => fifo_MEMWADDR(10), 
        B_ADDR(10) => fifo_MEMWADDR(9), B_ADDR(9) => 
        fifo_MEMWADDR(8), B_ADDR(8) => fifo_MEMWADDR(7), 
        B_ADDR(7) => fifo_MEMWADDR(6), B_ADDR(6) => 
        fifo_MEMWADDR(5), B_ADDR(5) => fifo_MEMWADDR(4), 
        B_ADDR(4) => fifo_MEMWADDR(3), B_ADDR(3) => 
        fifo_MEMWADDR(2), B_ADDR(2) => fifo_MEMWADDR(1), 
        B_ADDR(1) => fifo_MEMWADDR(0), B_ADDR(0) => GND_net_1, 
        B_WEN(1) => GND_net_1, B_WEN(0) => VCC_net_1, A_EN => 
        VCC_net_1, A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => 
        GND_net_1, A_WIDTH(1) => GND_net_1, A_WIDTH(0) => 
        VCC_net_1, A_WMODE => GND_net_1, B_EN => VCC_net_1, 
        B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => GND_net_1, 
        B_WIDTH(1) => GND_net_1, B_WIDTH(0) => VCC_net_1, B_WMODE
         => GND_net_1, SII_LOCK => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C1 : RAM1K18
      port map(A_DOUT(17) => nc158, A_DOUT(16) => nc162, 
        A_DOUT(15) => nc11, A_DOUT(14) => nc131, A_DOUT(13) => 
        nc96, A_DOUT(12) => nc79, A_DOUT(11) => nc146, A_DOUT(10)
         => nc89, A_DOUT(9) => nc119, A_DOUT(8) => nc48, 
        A_DOUT(7) => nc126, A_DOUT(6) => nc15, A_DOUT(5) => nc102, 
        A_DOUT(4) => nc3, A_DOUT(3) => nc47, A_DOUT(2) => nc90, 
        A_DOUT(1) => RDATA_int(3), A_DOUT(0) => RDATA_int(2), 
        B_DOUT(17) => nc159, B_DOUT(16) => nc136, B_DOUT(15) => 
        nc59, B_DOUT(14) => nc18, B_DOUT(13) => nc44, B_DOUT(12)
         => nc117, B_DOUT(11) => nc164, B_DOUT(10) => nc148, 
        B_DOUT(9) => nc42, B_DOUT(8) => nc17, B_DOUT(7) => nc2, 
        B_DOUT(6) => nc110, B_DOUT(5) => nc128, B_DOUT(4) => nc43, 
        B_DOUT(3) => nc157, B_DOUT(2) => nc36, B_DOUT(1) => nc61, 
        B_DOUT(0) => nc104, BUSY => OPEN, A_CLK => 
        m2s010_som_sb_0_CCC_71MHz, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => fifo_MEMRE, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => fifo_MEMRADDR(12), A_ADDR(12) => fifo_MEMRADDR(11), 
        A_ADDR(11) => fifo_MEMRADDR(10), A_ADDR(10) => 
        fifo_MEMRADDR(9), A_ADDR(9) => fifo_MEMRADDR(8), 
        A_ADDR(8) => fifo_MEMRADDR(7), A_ADDR(7) => 
        fifo_MEMRADDR(6), A_ADDR(6) => fifo_MEMRADDR(5), 
        A_ADDR(5) => fifo_MEMRADDR(4), A_ADDR(4) => 
        fifo_MEMRADDR(3), A_ADDR(3) => fifo_MEMRADDR(2), 
        A_ADDR(2) => fifo_MEMRADDR(1), A_ADDR(1) => 
        fifo_MEMRADDR(0), A_ADDR(0) => GND_net_1, A_WEN(1) => 
        GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => GND_net_1, B_DIN(2) => GND_net_1, B_DIN(1)
         => RX_FIFO_DIN_pipe(3), B_DIN(0) => RX_FIFO_DIN_pipe(2), 
        B_ADDR(13) => fifo_MEMWADDR(12), B_ADDR(12) => 
        fifo_MEMWADDR(11), B_ADDR(11) => fifo_MEMWADDR(10), 
        B_ADDR(10) => fifo_MEMWADDR(9), B_ADDR(9) => 
        fifo_MEMWADDR(8), B_ADDR(8) => fifo_MEMWADDR(7), 
        B_ADDR(7) => fifo_MEMWADDR(6), B_ADDR(6) => 
        fifo_MEMWADDR(5), B_ADDR(5) => fifo_MEMWADDR(4), 
        B_ADDR(4) => fifo_MEMWADDR(3), B_ADDR(3) => 
        fifo_MEMWADDR(2), B_ADDR(2) => fifo_MEMWADDR(1), 
        B_ADDR(1) => fifo_MEMWADDR(0), B_ADDR(0) => GND_net_1, 
        B_WEN(1) => GND_net_1, B_WEN(0) => VCC_net_1, A_EN => 
        VCC_net_1, A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => 
        GND_net_1, A_WIDTH(1) => GND_net_1, A_WIDTH(0) => 
        VCC_net_1, A_WMODE => GND_net_1, B_EN => VCC_net_1, 
        B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => GND_net_1, 
        B_WIDTH(1) => GND_net_1, B_WIDTH(0) => VCC_net_1, B_WMODE
         => GND_net_1, SII_LOCK => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C4 : RAM1K18
      port map(A_DOUT(17) => nc138, A_DOUT(16) => nc14, 
        A_DOUT(15) => nc150, A_DOUT(14) => nc149, A_DOUT(13) => 
        nc12, A_DOUT(12) => nc30, A_DOUT(11) => nc65, A_DOUT(10)
         => nc7, A_DOUT(9) => nc129, A_DOUT(8) => nc8, A_DOUT(7)
         => nc13, A_DOUT(6) => nc26, A_DOUT(5) => nc139, 
        A_DOUT(4) => nc163, A_DOUT(3) => nc112, A_DOUT(2) => nc68, 
        A_DOUT(1) => nc49, A_DOUT(0) => RDATA_int(8), B_DOUT(17)
         => nc170, B_DOUT(16) => nc91, B_DOUT(15) => nc5, 
        B_DOUT(14) => nc20, B_DOUT(13) => nc147, B_DOUT(12) => 
        nc67, B_DOUT(11) => nc152, B_DOUT(10) => nc127, B_DOUT(9)
         => nc103, B_DOUT(8) => nc76, B_DOUT(7) => nc140, 
        B_DOUT(6) => nc86, B_DOUT(5) => nc95, B_DOUT(4) => nc120, 
        B_DOUT(3) => nc165, B_DOUT(2) => nc137, B_DOUT(1) => nc64, 
        B_DOUT(0) => nc19, BUSY => OPEN, A_CLK => 
        m2s010_som_sb_0_CCC_71MHz, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => fifo_MEMRE, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => fifo_MEMRADDR(12), A_ADDR(12) => fifo_MEMRADDR(11), 
        A_ADDR(11) => fifo_MEMRADDR(10), A_ADDR(10) => 
        fifo_MEMRADDR(9), A_ADDR(9) => fifo_MEMRADDR(8), 
        A_ADDR(8) => fifo_MEMRADDR(7), A_ADDR(7) => 
        fifo_MEMRADDR(6), A_ADDR(6) => fifo_MEMRADDR(5), 
        A_ADDR(5) => fifo_MEMRADDR(4), A_ADDR(4) => 
        fifo_MEMRADDR(3), A_ADDR(3) => fifo_MEMRADDR(2), 
        A_ADDR(2) => fifo_MEMRADDR(1), A_ADDR(1) => 
        fifo_MEMRADDR(0), A_ADDR(0) => GND_net_1, A_WEN(1) => 
        GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => GND_net_1, B_DIN(2) => GND_net_1, B_DIN(1)
         => GND_net_1, B_DIN(0) => RX_FIFO_DIN_pipe(8), 
        B_ADDR(13) => fifo_MEMWADDR(12), B_ADDR(12) => 
        fifo_MEMWADDR(11), B_ADDR(11) => fifo_MEMWADDR(10), 
        B_ADDR(10) => fifo_MEMWADDR(9), B_ADDR(9) => 
        fifo_MEMWADDR(8), B_ADDR(8) => fifo_MEMWADDR(7), 
        B_ADDR(7) => fifo_MEMWADDR(6), B_ADDR(6) => 
        fifo_MEMWADDR(5), B_ADDR(5) => fifo_MEMWADDR(4), 
        B_ADDR(4) => fifo_MEMWADDR(3), B_ADDR(3) => 
        fifo_MEMWADDR(2), B_ADDR(2) => fifo_MEMWADDR(1), 
        B_ADDR(1) => fifo_MEMWADDR(0), B_ADDR(0) => GND_net_1, 
        B_WEN(1) => GND_net_1, B_WEN(0) => VCC_net_1, A_EN => 
        VCC_net_1, A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => 
        GND_net_1, A_WIDTH(1) => GND_net_1, A_WIDTH(0) => 
        VCC_net_1, A_WMODE => GND_net_1, B_EN => VCC_net_1, 
        B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => GND_net_1, 
        B_WIDTH(1) => GND_net_1, B_WIDTH(0) => VCC_net_1, B_WMODE
         => GND_net_1, SII_LOCK => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C3 : RAM1K18
      port map(A_DOUT(17) => nc70, A_DOUT(16) => nc62, A_DOUT(15)
         => nc80, A_DOUT(14) => nc130, A_DOUT(13) => nc98, 
        A_DOUT(12) => nc114, A_DOUT(11) => nc56, A_DOUT(10) => 
        nc105, A_DOUT(9) => nc63, A_DOUT(8) => nc97, A_DOUT(7)
         => nc161, A_DOUT(6) => nc31, A_DOUT(5) => nc154, 
        A_DOUT(4) => nc50, A_DOUT(3) => nc142, A_DOUT(2) => nc94, 
        A_DOUT(1) => RDATA_int(7), A_DOUT(0) => RDATA_int(6), 
        B_DOUT(17) => nc122, B_DOUT(16) => nc35, B_DOUT(15) => 
        nc4, B_DOUT(14) => nc92, B_DOUT(13) => nc101, B_DOUT(12)
         => nc166, B_DOUT(11) => nc132, B_DOUT(10) => nc21, 
        B_DOUT(9) => nc93, B_DOUT(8) => nc69, B_DOUT(7) => nc38, 
        B_DOUT(6) => nc113, B_DOUT(5) => nc106, B_DOUT(4) => nc25, 
        B_DOUT(3) => nc1, B_DOUT(2) => nc37, B_DOUT(1) => nc144, 
        B_DOUT(0) => nc153, BUSY => OPEN, A_CLK => 
        m2s010_som_sb_0_CCC_71MHz, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => fifo_MEMRE, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => fifo_MEMRADDR(12), A_ADDR(12) => fifo_MEMRADDR(11), 
        A_ADDR(11) => fifo_MEMRADDR(10), A_ADDR(10) => 
        fifo_MEMRADDR(9), A_ADDR(9) => fifo_MEMRADDR(8), 
        A_ADDR(8) => fifo_MEMRADDR(7), A_ADDR(7) => 
        fifo_MEMRADDR(6), A_ADDR(6) => fifo_MEMRADDR(5), 
        A_ADDR(5) => fifo_MEMRADDR(4), A_ADDR(4) => 
        fifo_MEMRADDR(3), A_ADDR(3) => fifo_MEMRADDR(2), 
        A_ADDR(2) => fifo_MEMRADDR(1), A_ADDR(1) => 
        fifo_MEMRADDR(0), A_ADDR(0) => GND_net_1, A_WEN(1) => 
        GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => GND_net_1, B_DIN(2) => GND_net_1, B_DIN(1)
         => RX_FIFO_DIN_pipe(7), B_DIN(0) => RX_FIFO_DIN_pipe(6), 
        B_ADDR(13) => fifo_MEMWADDR(12), B_ADDR(12) => 
        fifo_MEMWADDR(11), B_ADDR(11) => fifo_MEMWADDR(10), 
        B_ADDR(10) => fifo_MEMWADDR(9), B_ADDR(9) => 
        fifo_MEMWADDR(8), B_ADDR(8) => fifo_MEMWADDR(7), 
        B_ADDR(7) => fifo_MEMWADDR(6), B_ADDR(6) => 
        fifo_MEMWADDR(5), B_ADDR(5) => fifo_MEMWADDR(4), 
        B_ADDR(4) => fifo_MEMWADDR(3), B_ADDR(3) => 
        fifo_MEMWADDR(2), B_ADDR(2) => fifo_MEMWADDR(1), 
        B_ADDR(1) => fifo_MEMWADDR(0), B_ADDR(0) => GND_net_1, 
        B_WEN(1) => GND_net_1, B_WEN(0) => VCC_net_1, A_EN => 
        VCC_net_1, A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => 
        GND_net_1, A_WIDTH(1) => GND_net_1, A_WIDTH(0) => 
        VCC_net_1, A_WMODE => GND_net_1, B_EN => VCC_net_1, 
        B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => GND_net_1, 
        B_WIDTH(1) => GND_net_1, B_WIDTH(0) => VCC_net_1, B_WMODE
         => GND_net_1, SII_LOCK => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C0 : RAM1K18
      port map(A_DOUT(17) => nc46, A_DOUT(16) => nc71, A_DOUT(15)
         => nc124, A_DOUT(14) => nc81, A_DOUT(13) => nc168, 
        A_DOUT(12) => nc34, A_DOUT(11) => nc28, A_DOUT(10) => 
        nc115, A_DOUT(9) => nc134, A_DOUT(8) => nc32, A_DOUT(7)
         => nc40, A_DOUT(6) => nc99, A_DOUT(5) => nc75, A_DOUT(4)
         => nc85, A_DOUT(3) => nc27, A_DOUT(2) => nc108, 
        A_DOUT(1) => RDATA_int(1), A_DOUT(0) => RDATA_int(0), 
        B_DOUT(17) => nc16, B_DOUT(16) => nc155, B_DOUT(15) => 
        nc51, B_DOUT(14) => nc33, B_DOUT(13) => nc169, B_DOUT(12)
         => nc78, B_DOUT(11) => nc24, B_DOUT(10) => nc88, 
        B_DOUT(9) => nc111, B_DOUT(8) => nc55, B_DOUT(7) => nc10, 
        B_DOUT(6) => nc22, B_DOUT(5) => nc143, B_DOUT(4) => nc77, 
        B_DOUT(3) => nc6, B_DOUT(2) => nc109, B_DOUT(1) => nc87, 
        B_DOUT(0) => nc123, BUSY => OPEN, A_CLK => 
        m2s010_som_sb_0_CCC_71MHz, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => fifo_MEMRE, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => fifo_MEMRADDR(12), A_ADDR(12) => fifo_MEMRADDR(11), 
        A_ADDR(11) => fifo_MEMRADDR(10), A_ADDR(10) => 
        fifo_MEMRADDR(9), A_ADDR(9) => fifo_MEMRADDR(8), 
        A_ADDR(8) => fifo_MEMRADDR(7), A_ADDR(7) => 
        fifo_MEMRADDR(6), A_ADDR(6) => fifo_MEMRADDR(5), 
        A_ADDR(5) => fifo_MEMRADDR(4), A_ADDR(4) => 
        fifo_MEMRADDR(3), A_ADDR(3) => fifo_MEMRADDR(2), 
        A_ADDR(2) => fifo_MEMRADDR(1), A_ADDR(1) => 
        fifo_MEMRADDR(0), A_ADDR(0) => GND_net_1, A_WEN(1) => 
        GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => GND_net_1, B_DIN(2) => GND_net_1, B_DIN(1)
         => RX_FIFO_DIN_pipe(1), B_DIN(0) => RX_FIFO_DIN_pipe(0), 
        B_ADDR(13) => fifo_MEMWADDR(12), B_ADDR(12) => 
        fifo_MEMWADDR(11), B_ADDR(11) => fifo_MEMWADDR(10), 
        B_ADDR(10) => fifo_MEMWADDR(9), B_ADDR(9) => 
        fifo_MEMWADDR(8), B_ADDR(8) => fifo_MEMWADDR(7), 
        B_ADDR(7) => fifo_MEMWADDR(6), B_ADDR(6) => 
        fifo_MEMWADDR(5), B_ADDR(5) => fifo_MEMWADDR(4), 
        B_ADDR(4) => fifo_MEMWADDR(3), B_ADDR(3) => 
        fifo_MEMWADDR(2), B_ADDR(2) => fifo_MEMWADDR(1), 
        B_ADDR(1) => fifo_MEMWADDR(0), B_ADDR(0) => GND_net_1, 
        B_WEN(1) => GND_net_1, B_WEN(0) => VCC_net_1, A_EN => 
        VCC_net_1, A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => 
        GND_net_1, A_WIDTH(1) => GND_net_1, A_WIDTH(0) => 
        VCC_net_1, A_WMODE => GND_net_1, B_EN => VCC_net_1, 
        B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => GND_net_1, 
        B_WIDTH(1) => GND_net_1, B_WIDTH(0) => VCC_net_1, B_WMODE
         => GND_net_1, SII_LOCK => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_0 is

    port( fifo_MEMRADDR             : in    std_logic_vector(12 downto 0);
          fifo_MEMWADDR             : in    std_logic_vector(12 downto 0);
          RDATA_int                 : out   std_logic_vector(8 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          fifo_MEMRE                : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          fifo_MEMWE                : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_0;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_0
    port( RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          RDATA_int                 : out   std_logic_vector(8 downto 0);
          fifo_MEMWADDR             : in    std_logic_vector(12 downto 0) := (others => 'U');
          fifo_MEMRADDR             : in    std_logic_vector(12 downto 0) := (others => 'U');
          fifo_MEMWE                : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          fifo_MEMRE                : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_0
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_0(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    L1_asyncnonpipe : FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_0
      port map(RX_FIFO_DIN_pipe(8) => RX_FIFO_DIN_pipe(8), 
        RX_FIFO_DIN_pipe(7) => RX_FIFO_DIN_pipe(7), 
        RX_FIFO_DIN_pipe(6) => RX_FIFO_DIN_pipe(6), 
        RX_FIFO_DIN_pipe(5) => RX_FIFO_DIN_pipe(5), 
        RX_FIFO_DIN_pipe(4) => RX_FIFO_DIN_pipe(4), 
        RX_FIFO_DIN_pipe(3) => RX_FIFO_DIN_pipe(3), 
        RX_FIFO_DIN_pipe(2) => RX_FIFO_DIN_pipe(2), 
        RX_FIFO_DIN_pipe(1) => RX_FIFO_DIN_pipe(1), 
        RX_FIFO_DIN_pipe(0) => RX_FIFO_DIN_pipe(0), RDATA_int(8)
         => RDATA_int(8), RDATA_int(7) => RDATA_int(7), 
        RDATA_int(6) => RDATA_int(6), RDATA_int(5) => 
        RDATA_int(5), RDATA_int(4) => RDATA_int(4), RDATA_int(3)
         => RDATA_int(3), RDATA_int(2) => RDATA_int(2), 
        RDATA_int(1) => RDATA_int(1), RDATA_int(0) => 
        RDATA_int(0), fifo_MEMWADDR(12) => fifo_MEMWADDR(12), 
        fifo_MEMWADDR(11) => fifo_MEMWADDR(11), fifo_MEMWADDR(10)
         => fifo_MEMWADDR(10), fifo_MEMWADDR(9) => 
        fifo_MEMWADDR(9), fifo_MEMWADDR(8) => fifo_MEMWADDR(8), 
        fifo_MEMWADDR(7) => fifo_MEMWADDR(7), fifo_MEMWADDR(6)
         => fifo_MEMWADDR(6), fifo_MEMWADDR(5) => 
        fifo_MEMWADDR(5), fifo_MEMWADDR(4) => fifo_MEMWADDR(4), 
        fifo_MEMWADDR(3) => fifo_MEMWADDR(3), fifo_MEMWADDR(2)
         => fifo_MEMWADDR(2), fifo_MEMWADDR(1) => 
        fifo_MEMWADDR(1), fifo_MEMWADDR(0) => fifo_MEMWADDR(0), 
        fifo_MEMRADDR(12) => fifo_MEMRADDR(12), fifo_MEMRADDR(11)
         => fifo_MEMRADDR(11), fifo_MEMRADDR(10) => 
        fifo_MEMRADDR(10), fifo_MEMRADDR(9) => fifo_MEMRADDR(9), 
        fifo_MEMRADDR(8) => fifo_MEMRADDR(8), fifo_MEMRADDR(7)
         => fifo_MEMRADDR(7), fifo_MEMRADDR(6) => 
        fifo_MEMRADDR(6), fifo_MEMRADDR(5) => fifo_MEMRADDR(5), 
        fifo_MEMRADDR(4) => fifo_MEMRADDR(4), fifo_MEMRADDR(3)
         => fifo_MEMRADDR(3), fifo_MEMRADDR(2) => 
        fifo_MEMRADDR(2), fifo_MEMRADDR(1) => fifo_MEMRADDR(1), 
        fifo_MEMRADDR(0) => fifo_MEMRADDR(0), fifo_MEMWE => 
        fifo_MEMWE, CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, 
        fifo_MEMRE => fifo_MEMRE, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_2 is

    port( wptr_bin_sync  : inout std_logic_vector(13 downto 0) := (others => 'Z');
          wptr_gray_sync : in    std_logic_vector(12 downto 0)
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_2;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_2 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    \bin_out_xhdl1_0_a2[1]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(3), B => wptr_gray_sync(1), C
         => wptr_bin_sync(4), D => wptr_gray_sync(2), Y => 
        wptr_bin_sync(1));
    
    \bin_out_xhdl1_0_a2[10]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(12), B => wptr_gray_sync(11), 
        C => wptr_gray_sync(10), D => wptr_bin_sync(13), Y => 
        wptr_bin_sync(10));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \bin_out_xhdl1_0_a2[5]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(7), B => wptr_gray_sync(6), C
         => wptr_gray_sync(5), D => wptr_bin_sync(8), Y => 
        wptr_bin_sync(5));
    
    \bin_out_xhdl1_0_a2[2]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(4), B => wptr_gray_sync(3), C
         => wptr_gray_sync(2), D => wptr_bin_sync(5), Y => 
        wptr_bin_sync(2));
    
    \bin_out_xhdl1_0_a2[0]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(2), B => wptr_bin_sync(3), C
         => wptr_gray_sync(0), D => wptr_gray_sync(1), Y => 
        wptr_bin_sync(0));
    
    \bin_out_xhdl1_0_a2[9]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(11), B => wptr_gray_sync(10), 
        C => wptr_gray_sync(9), D => wptr_bin_sync(12), Y => 
        wptr_bin_sync(9));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \bin_out_xhdl1_i_o2[12]\ : CFG2
      generic map(INIT => x"6")

      port map(A => wptr_bin_sync(13), B => wptr_gray_sync(12), Y
         => wptr_bin_sync(12));
    
    \bin_out_xhdl1_0_a2[6]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(8), B => wptr_gray_sync(7), C
         => wptr_gray_sync(6), D => wptr_bin_sync(9), Y => 
        wptr_bin_sync(6));
    
    \bin_out_xhdl1_0_a2[4]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(6), B => wptr_gray_sync(5), C
         => wptr_gray_sync(4), D => wptr_bin_sync(7), Y => 
        wptr_bin_sync(4));
    
    \bin_out_xhdl1_i_o2[11]\ : CFG3
      generic map(INIT => x"96")

      port map(A => wptr_gray_sync(12), B => wptr_gray_sync(11), 
        C => wptr_bin_sync(13), Y => wptr_bin_sync(11));
    
    \bin_out_xhdl1_0_a2[8]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(10), B => wptr_gray_sync(9), C
         => wptr_gray_sync(8), D => wptr_bin_sync(11), Y => 
        wptr_bin_sync(8));
    
    \bin_out_xhdl1_0_a2[7]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(9), B => wptr_gray_sync(8), C
         => wptr_gray_sync(7), D => wptr_bin_sync(10), Y => 
        wptr_bin_sync(7));
    
    \bin_out_xhdl1_0_a2[3]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(5), B => wptr_gray_sync(4), C
         => wptr_gray_sync(3), D => wptr_bin_sync(6), Y => 
        wptr_bin_sync(3));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_1 is

    port( wptr_gray                 : in    std_logic_vector(13 downto 0);
          wptr_gray_sync            : out   std_logic_vector(12 downto 0);
          wptr_bin_sync_0           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          irx_fifo_rst_i            : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_1;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_1 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \sync_int[11]_net_1\, GND_net_1, 
        \sync_int[12]_net_1\, \sync_int[13]_net_1\, 
        \sync_int[10]_net_1\, \sync_int[0]_net_1\, 
        \sync_int[1]_net_1\, \sync_int[2]_net_1\, 
        \sync_int[3]_net_1\, \sync_int[4]_net_1\, 
        \sync_int[5]_net_1\, \sync_int[6]_net_1\, 
        \sync_int[7]_net_1\, \sync_int[8]_net_1\, 
        \sync_int[9]_net_1\ : std_logic;

begin 


    \sync_int[9]\ : SLE
      port map(D => wptr_gray(9), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[9]_net_1\);
    
    \sync_int[4]\ : SLE
      port map(D => wptr_gray(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[4]_net_1\);
    
    \sync_out_xhdl1[10]\ : SLE
      port map(D => \sync_int[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(10));
    
    \sync_int[1]\ : SLE
      port map(D => wptr_gray(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[1]_net_1\);
    
    \sync_int[11]\ : SLE
      port map(D => wptr_gray(11), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[11]_net_1\);
    
    \sync_out_xhdl1[6]\ : SLE
      port map(D => \sync_int[6]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(6));
    
    \sync_out_xhdl1[3]\ : SLE
      port map(D => \sync_int[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(3));
    
    \sync_int[6]\ : SLE
      port map(D => wptr_gray(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[6]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \sync_out_xhdl1[11]\ : SLE
      port map(D => \sync_int[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(11));
    
    \sync_int[13]\ : SLE
      port map(D => wptr_gray(13), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[13]_net_1\);
    
    \sync_int[3]\ : SLE
      port map(D => wptr_gray(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[3]_net_1\);
    
    \sync_int[12]\ : SLE
      port map(D => wptr_gray(12), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[12]_net_1\);
    
    \sync_out_xhdl1[4]\ : SLE
      port map(D => \sync_int[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(4));
    
    \sync_int[0]\ : SLE
      port map(D => wptr_gray(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[0]_net_1\);
    
    \sync_out_xhdl1[1]\ : SLE
      port map(D => \sync_int[1]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(1));
    
    \sync_int[5]\ : SLE
      port map(D => wptr_gray(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[5]_net_1\);
    
    \sync_int[2]\ : SLE
      port map(D => wptr_gray(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[2]_net_1\);
    
    \sync_out_xhdl1[12]\ : SLE
      port map(D => \sync_int[12]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(12));
    
    \sync_out_xhdl1[9]\ : SLE
      port map(D => \sync_int[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(9));
    
    \sync_out_xhdl1[2]\ : SLE
      port map(D => \sync_int[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(2));
    
    \sync_int[8]\ : SLE
      port map(D => wptr_gray(8), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[8]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sync_out_xhdl1[7]\ : SLE
      port map(D => \sync_int[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(7));
    
    \sync_out_xhdl1[5]\ : SLE
      port map(D => \sync_int[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(5));
    
    \sync_out_xhdl1[0]\ : SLE
      port map(D => \sync_int[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(0));
    
    \sync_out_xhdl1[8]\ : SLE
      port map(D => \sync_int[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(8));
    
    \sync_int[7]\ : SLE
      port map(D => wptr_gray(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[7]_net_1\);
    
    \sync_int[10]\ : SLE
      port map(D => wptr_gray(10), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[10]_net_1\);
    
    \sync_out_xhdl1[13]\ : SLE
      port map(D => \sync_int[13]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_bin_sync_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_0 is

    port( rptr_gray           : in    std_logic_vector(13 downto 0);
          rptr_gray_sync      : out   std_logic_vector(12 downto 0);
          rptr_bin_sync_0     : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          irx_fifo_rst_i      : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_0;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_0 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \sync_int[13]_net_1\, GND_net_1, 
        \sync_int[12]_net_1\, \sync_int[0]_net_1\, 
        \sync_int[1]_net_1\, \sync_int[2]_net_1\, 
        \sync_int[3]_net_1\, \sync_int[4]_net_1\, 
        \sync_int[5]_net_1\, \sync_int[6]_net_1\, 
        \sync_int[7]_net_1\, \sync_int[8]_net_1\, 
        \sync_int[9]_net_1\, \sync_int[10]_net_1\, 
        \sync_int[11]_net_1\ : std_logic;

begin 


    \sync_int[9]\ : SLE
      port map(D => rptr_gray(9), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[9]_net_1\);
    
    \sync_int[4]\ : SLE
      port map(D => rptr_gray(4), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[4]_net_1\);
    
    \sync_out_xhdl1[10]\ : SLE
      port map(D => \sync_int[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(10));
    
    \sync_int[1]\ : SLE
      port map(D => rptr_gray(1), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[1]_net_1\);
    
    \sync_int[11]\ : SLE
      port map(D => rptr_gray(11), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[11]_net_1\);
    
    \sync_out_xhdl1[6]\ : SLE
      port map(D => \sync_int[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(6));
    
    \sync_out_xhdl1[3]\ : SLE
      port map(D => \sync_int[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(3));
    
    \sync_int[6]\ : SLE
      port map(D => rptr_gray(6), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[6]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \sync_out_xhdl1[11]\ : SLE
      port map(D => \sync_int[11]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(11));
    
    \sync_int[13]\ : SLE
      port map(D => rptr_gray(13), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[13]_net_1\);
    
    \sync_int[3]\ : SLE
      port map(D => rptr_gray(3), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[3]_net_1\);
    
    \sync_int[12]\ : SLE
      port map(D => rptr_gray(12), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[12]_net_1\);
    
    \sync_out_xhdl1[4]\ : SLE
      port map(D => \sync_int[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(4));
    
    \sync_int[0]\ : SLE
      port map(D => rptr_gray(0), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[0]_net_1\);
    
    \sync_out_xhdl1[1]\ : SLE
      port map(D => \sync_int[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(1));
    
    \sync_int[5]\ : SLE
      port map(D => rptr_gray(5), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[5]_net_1\);
    
    \sync_int[2]\ : SLE
      port map(D => rptr_gray(2), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[2]_net_1\);
    
    \sync_out_xhdl1[12]\ : SLE
      port map(D => \sync_int[12]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(12));
    
    \sync_out_xhdl1[9]\ : SLE
      port map(D => \sync_int[9]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(9));
    
    \sync_out_xhdl1[2]\ : SLE
      port map(D => \sync_int[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(2));
    
    \sync_int[8]\ : SLE
      port map(D => rptr_gray(8), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[8]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sync_out_xhdl1[7]\ : SLE
      port map(D => \sync_int[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(7));
    
    \sync_out_xhdl1[5]\ : SLE
      port map(D => \sync_int[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(5));
    
    \sync_out_xhdl1[0]\ : SLE
      port map(D => \sync_int[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(0));
    
    \sync_out_xhdl1[8]\ : SLE
      port map(D => \sync_int[8]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(8));
    
    \sync_int[7]\ : SLE
      port map(D => rptr_gray(7), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[7]_net_1\);
    
    \sync_int[10]\ : SLE
      port map(D => rptr_gray(10), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[10]_net_1\);
    
    \sync_out_xhdl1[13]\ : SLE
      port map(D => \sync_int[13]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_bin_sync_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_1 is

    port( rptr_bin_sync  : inout std_logic_vector(13 downto 0) := (others => 'Z');
          rptr_gray_sync : in    std_logic_vector(12 downto 0);
          bin_N_6_i      : out   std_logic;
          bin_N_4_0_i    : out   std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_1;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_1 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \bin_m5_5\, \bin_m5_4\, \bin_m3_0_3\, \bin_N_4_0_i\, 
        GND_net_1, VCC_net_1 : std_logic;

begin 

    bin_N_4_0_i <= \bin_N_4_0_i\;

    bin_m5_4 : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(4), B => rptr_gray_sync(6), C
         => rptr_gray_sync(5), D => rptr_gray_sync(10), Y => 
        \bin_m5_4\);
    
    \bin_out_xhdl1_0_a2[10]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(12), B => rptr_gray_sync(10), 
        C => rptr_gray_sync(11), D => rptr_bin_sync(13), Y => 
        rptr_bin_sync(10));
    
    \bin_out_xhdl1_0_a2[8]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(8), B => rptr_gray_sync(9), C
         => rptr_bin_sync(10), Y => rptr_bin_sync(8));
    
    bin_m5_5 : CFG4
      generic map(INIT => x"9669")

      port map(A => rptr_gray_sync(8), B => rptr_gray_sync(9), C
         => rptr_gray_sync(7), D => rptr_gray_sync(11), Y => 
        \bin_m5_5\);
    
    bin_m3_0_3 : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(7), B => rptr_gray_sync(9), C
         => rptr_gray_sync(6), D => rptr_gray_sync(10), Y => 
        \bin_m3_0_3\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \bin_out_xhdl1_0_a2[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(3), B => rptr_gray_sync(2), Y
         => rptr_bin_sync(2));
    
    \bin_out_xhdl1_0_a2[1]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(1), B => rptr_gray_sync(2), C
         => rptr_bin_sync(3), Y => rptr_bin_sync(1));
    
    \bin_out_xhdl1_0_a2[0]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(1), B => rptr_gray_sync(0), C
         => rptr_bin_sync(3), D => rptr_gray_sync(2), Y => 
        rptr_bin_sync(0));
    
    \bin_out_xhdl1_i_o2_RNIA8NV1[12]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(8), B => rptr_gray_sync(11), C
         => rptr_bin_sync(12), D => \bin_m3_0_3\, Y => 
        \bin_N_4_0_i\);
    
    \bin_out_xhdl1_i_o2[11]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(11), B => rptr_bin_sync(13), C
         => rptr_gray_sync(12), Y => rptr_bin_sync(11));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \bin_out_xhdl1_0_a2[7]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(9), B => rptr_bin_sync(10), C
         => rptr_gray_sync(7), D => rptr_gray_sync(8), Y => 
        rptr_bin_sync(7));
    
    \bin_out_xhdl1_0_a2[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \bin_N_4_0_i\, B => rptr_gray_sync(5), Y => 
        rptr_bin_sync(5));
    
    \bin_out_xhdl1_i_o2_RNIPGFI2[12]\ : CFG3
      generic map(INIT => x"69")

      port map(A => \bin_m5_5\, B => \bin_m5_4\, C => 
        rptr_bin_sync(12), Y => bin_N_6_i);
    
    \bin_out_xhdl1_i_o2[12]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(13), B => rptr_gray_sync(12), Y
         => rptr_bin_sync(12));
    
    \bin_out_xhdl1_0_a2[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(10), B => rptr_gray_sync(9), Y
         => rptr_bin_sync(9));
    
    \bin_out_xhdl1_0_a2[3]\ : CFG4
      generic map(INIT => x"9669")

      port map(A => rptr_bin_sync(12), B => \bin_m5_5\, C => 
        rptr_gray_sync(3), D => \bin_m5_4\, Y => rptr_bin_sync(3));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_0 is

    port( fifo_MEMRADDR             : out   std_logic_vector(12 downto 0);
          fifo_MEMWADDR             : out   std_logic_vector(12 downto 0);
          iRX_FIFO_wr_en_0_0        : in    std_logic;
          iRX_FIFO_rd_en_0          : in    std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          RX_FIFO_TxColDetDis_wr_en : in    std_logic;
          fifo_MEMRE                : out   std_logic;
          fifo_MEMWE                : out   std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          irx_fifo_rst_i            : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_0;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_0 is 

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_2
    port( wptr_bin_sync  : inout   std_logic_vector(13 downto 0);
          wptr_gray_sync : in    std_logic_vector(12 downto 0) := (others => 'U')
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_1
    port( wptr_gray                 : in    std_logic_vector(13 downto 0) := (others => 'U');
          wptr_gray_sync            : out   std_logic_vector(12 downto 0);
          wptr_bin_sync_0           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          irx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_0
    port( rptr_gray           : in    std_logic_vector(13 downto 0) := (others => 'U');
          rptr_gray_sync      : out   std_logic_vector(12 downto 0);
          rptr_bin_sync_0     : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          irx_fifo_rst_i      : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_1
    port( rptr_bin_sync  : inout   std_logic_vector(13 downto 0);
          rptr_gray_sync : in    std_logic_vector(12 downto 0) := (others => 'U');
          bin_N_6_i      : out   std_logic;
          bin_N_4_0_i    : out   std_logic
        );
  end component;

    signal \rptr[0]_net_1\, \rptr_s[0]\, \wptr[0]_net_1\, 
        \wptr_s[0]\, \fifo_MEMRADDR[0]\, \fifo_MEMRADDR_i[0]\, 
        \fifo_MEMWADDR[0]\, \fifo_MEMWADDR_i[0]\, 
        \rptr_gray[1]_net_1\, VCC_net_1, \rptr_gray_1[1]_net_1\, 
        GND_net_1, \rptr_gray[2]_net_1\, \rptr_gray_1[2]_net_1\, 
        \rptr_gray[3]_net_1\, \rptr_gray_1[3]_net_1\, 
        \rptr_gray[4]_net_1\, \rptr_gray_1[4]_net_1\, 
        \rptr_gray[5]_net_1\, \rptr_gray_1[5]_net_1\, 
        \rptr_gray[6]_net_1\, \rptr_gray_1[6]_net_1\, 
        \rptr_gray[7]_net_1\, \rptr_gray_1[7]_net_1\, 
        \rptr_gray[8]_net_1\, \rptr_gray_1[8]_net_1\, 
        \rptr_gray[9]_net_1\, \rptr_gray_1[9]_net_1\, 
        \rptr_gray[10]_net_1\, \rptr_gray_1[10]_net_1\, 
        \rptr_gray[11]_net_1\, \rptr_gray_1[11]_net_1\, 
        \rptr_gray[12]_net_1\, \rptr_gray_1[12]_net_1\, 
        \rptr_gray[13]_net_1\, \rptr[13]_net_1\, 
        \wptr_gray[0]_net_1\, \wptr_gray_1[0]_net_1\, 
        \wptr_gray[1]_net_1\, \wptr_gray_1[1]_net_1\, 
        \wptr_gray[2]_net_1\, \wptr_gray_1[2]_net_1\, 
        \wptr_gray[3]_net_1\, \wptr_gray_1[3]_net_1\, 
        \wptr_gray[4]_net_1\, \wptr_gray_1[4]_net_1\, 
        \wptr_gray[5]_net_1\, \wptr_gray_1[5]_net_1\, 
        \wptr_gray[6]_net_1\, \wptr_gray_1[6]_net_1\, 
        \wptr_gray[7]_net_1\, \wptr_gray_1[7]_net_1\, 
        \wptr_gray[8]_net_1\, \wptr_gray_1[8]_net_1\, 
        \wptr_gray[9]_net_1\, \wptr_gray_1[9]_net_1\, 
        \wptr_gray[10]_net_1\, \wptr_gray_1[10]_net_1\, 
        \wptr_gray[11]_net_1\, \wptr_gray_1[11]_net_1\, 
        \wptr_gray[12]_net_1\, \wptr_gray_1[12]_net_1\, 
        \wptr_gray[13]_net_1\, \wptr[13]_net_1\, 
        \rptr_gray[0]_net_1\, \rptr_gray_1[0]_net_1\, rdiff_bus, 
        \wptr_bin_sync[0]\, \wptr_bin_sync2[1]_net_1\, 
        \wptr_bin_sync[1]\, \wptr_bin_sync2[2]_net_1\, 
        \wptr_bin_sync[2]\, \wptr_bin_sync2[3]_net_1\, 
        \wptr_bin_sync[3]\, \wptr_bin_sync2[4]_net_1\, 
        \wptr_bin_sync[4]\, \wptr_bin_sync2[5]_net_1\, 
        \wptr_bin_sync[5]\, \wptr_bin_sync2[6]_net_1\, 
        \wptr_bin_sync[6]\, \wptr_bin_sync2[7]_net_1\, 
        \wptr_bin_sync[7]\, \wptr_bin_sync2[8]_net_1\, 
        \wptr_bin_sync[8]\, \wptr_bin_sync2[9]_net_1\, 
        \wptr_bin_sync[9]\, \wptr_bin_sync2[10]_net_1\, 
        \wptr_bin_sync[10]\, \wptr_bin_sync2[11]_net_1\, 
        \wptr_bin_sync[11]\, \wptr_bin_sync2[12]_net_1\, 
        \wptr_bin_sync[12]\, \wptr_bin_sync2[13]_net_1\, 
        \wptr_bin_sync[13]\, \rptr_bin_sync2[9]_net_1\, 
        \rptr_bin_sync[9]\, \rptr_bin_sync2[10]_net_1\, 
        \rptr_bin_sync[10]\, \rptr_bin_sync2[11]_net_1\, 
        \rptr_bin_sync[11]\, \rptr_bin_sync2[12]_net_1\, 
        \rptr_bin_sync[12]\, \rptr_bin_sync2[13]_net_1\, 
        \rptr_bin_sync[13]\, \fifo_MEMWADDR[7]\, 
        \memwaddr_r_2[7]_net_1\, \fifo_MEMWE\, \fifo_MEMWADDR[8]\, 
        \memwaddr_r_2[8]_net_1\, \fifo_MEMWADDR[9]\, 
        \memwaddr_r_2[9]_net_1\, \fifo_MEMWADDR[10]\, 
        \memwaddr_r_2[10]_net_1\, \fifo_MEMWADDR[11]\, 
        \memwaddr_r_2[11]_net_1\, \fifo_MEMWADDR[12]\, 
        \memwaddr_r_2[12]_net_1\, \rptr_bin_sync2[0]_net_1\, 
        \rptr_bin_sync[0]\, \rptr_bin_sync2[1]_net_1\, 
        \rptr_bin_sync[1]\, \rptr_bin_sync2[2]_net_1\, 
        \rptr_bin_sync[2]\, \rptr_bin_sync2[3]_net_1\, 
        \rptr_bin_sync[3]\, \rptr_bin_sync2[4]_net_1\, bin_N_6_i, 
        \rptr_bin_sync2[5]_net_1\, \rptr_bin_sync[5]\, 
        \rptr_bin_sync2[6]_net_1\, bin_N_4_0_i, 
        \rptr_bin_sync2[7]_net_1\, \rptr_bin_sync[7]\, 
        \rptr_bin_sync2[8]_net_1\, \rptr_bin_sync[8]\, 
        \fifo_MEMRADDR[5]\, \memraddr_r_2[5]_net_1\, \fifo_MEMRE\, 
        \fifo_MEMRADDR[6]\, un1_memraddr_r_cry_6_S_0, 
        \fifo_MEMRADDR[7]\, \memraddr_r_2[7]_net_1\, 
        \fifo_MEMRADDR[8]\, \memraddr_r_2[8]_net_1\, 
        \fifo_MEMRADDR[9]\, \memraddr_r_2[9]_net_1\, 
        \fifo_MEMRADDR[10]\, \memraddr_r_2[10]_net_1\, 
        \fifo_MEMRADDR[11]\, \memraddr_r_2[11]_net_1\, 
        \fifo_MEMRADDR[12]\, \memraddr_r_2[12]_net_1\, 
        \fifo_MEMWADDR[1]\, un1_memwaddr_r_cry_1_S_0, 
        \fifo_MEMWADDR[2]\, un1_memwaddr_r_cry_2_S_0, 
        \fifo_MEMWADDR[3]\, un1_memwaddr_r_cry_3_S_0, 
        \fifo_MEMWADDR[4]\, un1_memwaddr_r_cry_4_S_0, 
        \fifo_MEMWADDR[5]\, \memwaddr_r_2[5]_net_1\, 
        \fifo_MEMWADDR[6]\, un1_memwaddr_r_cry_6_S_0, 
        \fifo_MEMRADDR[1]\, un1_memraddr_r_cry_1_S_0, 
        \fifo_MEMRADDR[2]\, un1_memraddr_r_cry_2_S_0, 
        \fifo_MEMRADDR[3]\, un1_memraddr_r_cry_3_S_0, 
        \fifo_MEMRADDR[4]\, un1_memraddr_r_cry_4_S_0, 
        \iRX_FIFO_Full_0\, fulli, N_6_i, N_5_i, 
        \iRX_FIFO_Empty_0\, empty_r_3, \wptr[1]_net_1\, 
        \wptr_s[1]\, \wptr[2]_net_1\, \wptr_s[2]\, 
        \wptr[3]_net_1\, \wptr_s[3]\, \wptr[4]_net_1\, 
        \wptr_s[4]\, \wptr[5]_net_1\, \wptr_s[5]\, 
        \wptr[6]_net_1\, \wptr_s[6]\, \wptr[7]_net_1\, 
        \wptr_s[7]\, \wptr[8]_net_1\, \wptr_s[8]\, 
        \wptr[9]_net_1\, \wptr_s[9]\, \wptr[10]_net_1\, 
        \wptr_s[10]\, \wptr[11]_net_1\, \wptr_s[11]\, 
        \wptr[12]_net_1\, \wptr_s[12]\, \wptr_s[13]_net_1\, 
        \rptr[1]_net_1\, \rptr_s[1]\, \rptr[2]_net_1\, 
        \rptr_s[2]\, \rptr[3]_net_1\, \rptr_s[3]\, 
        \rptr[4]_net_1\, \rptr_s[4]\, \rptr[5]_net_1\, 
        \rptr_s[5]\, \rptr[6]_net_1\, \rptr_s[6]\, 
        \rptr[7]_net_1\, \rptr_s[7]\, \rptr[8]_net_1\, 
        \rptr_s[8]\, \rptr[9]_net_1\, \rptr_s[9]\, 
        \rptr[10]_net_1\, \rptr_s[10]\, \rptr[11]_net_1\, 
        \rptr_s[11]\, \rptr[12]_net_1\, \rptr_s[12]\, 
        \rptr_s[13]_net_1\, \rdiff_bus_cry_0\, 
        rdiff_bus_cry_0_Y_1, \rdiff_bus_cry_1\, \rdiff_bus[1]\, 
        \rdiff_bus_cry_2\, \rdiff_bus[2]\, \rdiff_bus_cry_3\, 
        \rdiff_bus[3]\, \rdiff_bus_cry_4\, \rdiff_bus[4]\, 
        \rdiff_bus_cry_5\, \rdiff_bus[5]\, \rdiff_bus_cry_6\, 
        \rdiff_bus[6]\, \rdiff_bus_cry_7\, \rdiff_bus[7]\, 
        \rdiff_bus_cry_8\, \rdiff_bus[8]\, \rdiff_bus_cry_9\, 
        \rdiff_bus[9]\, \rdiff_bus_cry_10\, \rdiff_bus[10]\, 
        \rdiff_bus_cry_11\, \rdiff_bus[11]\, \rdiff_bus[13]\, 
        \rdiff_bus_cry_12\, \rdiff_bus[12]\, \wdiff_bus_cry_0\, 
        wdiff_bus_cry_0_Y_1, \wdiff_bus_cry_1\, \wdiff_bus[1]\, 
        \wdiff_bus_cry_2\, \wdiff_bus[2]\, \wdiff_bus_cry_3\, 
        \wdiff_bus[3]\, \wdiff_bus_cry_4\, \wdiff_bus[4]\, 
        \wdiff_bus_cry_5\, \wdiff_bus[5]\, \wdiff_bus_cry_6\, 
        \wdiff_bus[6]\, \wdiff_bus_cry_7\, \wdiff_bus[7]\, 
        \wdiff_bus_cry_8\, \wdiff_bus[8]\, \wdiff_bus_cry_9\, 
        \wdiff_bus[9]\, \wdiff_bus_cry_10\, \wdiff_bus[10]\, 
        \wdiff_bus_cry_11\, \wdiff_bus[11]\, \wdiff_bus[13]\, 
        \wdiff_bus_cry_12\, \wdiff_bus[12]\, rptr_s_906_FCO, 
        \rptr_cry[1]_net_1\, \rptr_cry[2]_net_1\, 
        \rptr_cry[3]_net_1\, \rptr_cry[4]_net_1\, 
        \rptr_cry[5]_net_1\, \rptr_cry[6]_net_1\, 
        \rptr_cry[7]_net_1\, \rptr_cry[8]_net_1\, 
        \rptr_cry[9]_net_1\, \rptr_cry[10]_net_1\, 
        \rptr_cry[11]_net_1\, \rptr_cry[12]_net_1\, 
        wptr_s_907_FCO, \wptr_cry[1]_net_1\, \wptr_cry[2]_net_1\, 
        \wptr_cry[3]_net_1\, \wptr_cry[4]_net_1\, 
        \wptr_cry[5]_net_1\, \wptr_cry[6]_net_1\, 
        \wptr_cry[7]_net_1\, \wptr_cry[8]_net_1\, 
        \wptr_cry[9]_net_1\, \wptr_cry[10]_net_1\, 
        \wptr_cry[11]_net_1\, \wptr_cry[12]_net_1\, 
        un1_memraddr_r_s_1_925_FCO, \un1_memraddr_r_cry_1\, 
        \un1_memraddr_r_cry_2\, \un1_memraddr_r_cry_3\, 
        \un1_memraddr_r_cry_4\, \un1_memraddr_r_cry_5\, 
        un1_memraddr_r_cry_5_S_0, \un1_memraddr_r_cry_6\, 
        \un1_memraddr_r_cry_7\, un1_memraddr_r_cry_7_S_0, 
        \un1_memraddr_r_cry_8\, un1_memraddr_r_cry_8_S_0, 
        \un1_memraddr_r_cry_9\, un1_memraddr_r_cry_9_S_0, 
        \un1_memraddr_r_cry_10\, un1_memraddr_r_cry_10_S_0, 
        un1_memraddr_r_s_12_S_0, \un1_memraddr_r_cry_11\, 
        un1_memraddr_r_cry_11_S_0, un1_memwaddr_r_s_1_926_FCO, 
        \un1_memwaddr_r_cry_1\, \un1_memwaddr_r_cry_2\, 
        \un1_memwaddr_r_cry_3\, \un1_memwaddr_r_cry_4\, 
        \un1_memwaddr_r_cry_5\, un1_memwaddr_r_cry_5_S_0, 
        \un1_memwaddr_r_cry_6\, \un1_memwaddr_r_cry_7\, 
        un1_memwaddr_r_cry_7_S_0, \un1_memwaddr_r_cry_8\, 
        un1_memwaddr_r_cry_8_S_0, \un1_memwaddr_r_cry_9\, 
        un1_memwaddr_r_cry_9_S_0, \un1_memwaddr_r_cry_10\, 
        un1_memwaddr_r_cry_10_S_0, un1_memwaddr_r_s_12_S_0, 
        \un1_memwaddr_r_cry_11\, un1_memwaddr_r_cry_11_S_0, 
        \fulli_0_a3_5_1\, \fulli_0_a3_4_3\, \fulli_0_a3_d_4\, 
        un4_re_i_0, un4_we_i_0, empty_r_3_0_a2_9, 
        empty_r_3_0_a2_8, empty_r_3_0_a2_7, un4_re_i_8, 
        un4_re_i_7, un4_we_i_8, un4_we_i_7, un4_re_i_9, 
        un4_we_i_9, \fulli_0_a3_d_3\, empty_r_3_0_a2_6, 
        \wptr_gray_sync[0]\, \wptr_gray_sync[1]\, 
        \wptr_gray_sync[2]\, \wptr_gray_sync[3]\, 
        \wptr_gray_sync[4]\, \wptr_gray_sync[5]\, 
        \wptr_gray_sync[6]\, \wptr_gray_sync[7]\, 
        \wptr_gray_sync[8]\, \wptr_gray_sync[9]\, 
        \wptr_gray_sync[10]\, \wptr_gray_sync[11]\, 
        \wptr_gray_sync[12]\, \rptr_gray_sync[0]\, 
        \rptr_gray_sync[1]\, \rptr_gray_sync[2]\, 
        \rptr_gray_sync[3]\, \rptr_gray_sync[4]\, 
        \rptr_gray_sync[5]\, \rptr_gray_sync[6]\, 
        \rptr_gray_sync[7]\, \rptr_gray_sync[8]\, 
        \rptr_gray_sync[9]\, \rptr_gray_sync[10]\, 
        \rptr_gray_sync[11]\, \rptr_gray_sync[12]\ : std_logic;
    signal nc2, nc1 : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_2
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_2(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_1
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_1(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_0
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_0(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_1
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_1(DEF_ARCH);
begin 

    fifo_MEMRADDR(12) <= \fifo_MEMRADDR[12]\;
    fifo_MEMRADDR(11) <= \fifo_MEMRADDR[11]\;
    fifo_MEMRADDR(10) <= \fifo_MEMRADDR[10]\;
    fifo_MEMRADDR(9) <= \fifo_MEMRADDR[9]\;
    fifo_MEMRADDR(8) <= \fifo_MEMRADDR[8]\;
    fifo_MEMRADDR(7) <= \fifo_MEMRADDR[7]\;
    fifo_MEMRADDR(6) <= \fifo_MEMRADDR[6]\;
    fifo_MEMRADDR(5) <= \fifo_MEMRADDR[5]\;
    fifo_MEMRADDR(4) <= \fifo_MEMRADDR[4]\;
    fifo_MEMRADDR(3) <= \fifo_MEMRADDR[3]\;
    fifo_MEMRADDR(2) <= \fifo_MEMRADDR[2]\;
    fifo_MEMRADDR(1) <= \fifo_MEMRADDR[1]\;
    fifo_MEMRADDR(0) <= \fifo_MEMRADDR[0]\;
    fifo_MEMWADDR(12) <= \fifo_MEMWADDR[12]\;
    fifo_MEMWADDR(11) <= \fifo_MEMWADDR[11]\;
    fifo_MEMWADDR(10) <= \fifo_MEMWADDR[10]\;
    fifo_MEMWADDR(9) <= \fifo_MEMWADDR[9]\;
    fifo_MEMWADDR(8) <= \fifo_MEMWADDR[8]\;
    fifo_MEMWADDR(7) <= \fifo_MEMWADDR[7]\;
    fifo_MEMWADDR(6) <= \fifo_MEMWADDR[6]\;
    fifo_MEMWADDR(5) <= \fifo_MEMWADDR[5]\;
    fifo_MEMWADDR(4) <= \fifo_MEMWADDR[4]\;
    fifo_MEMWADDR(3) <= \fifo_MEMWADDR[3]\;
    fifo_MEMWADDR(2) <= \fifo_MEMWADDR[2]\;
    fifo_MEMWADDR(1) <= \fifo_MEMWADDR[1]\;
    fifo_MEMWADDR(0) <= \fifo_MEMWADDR[0]\;
    iRX_FIFO_Empty_0 <= \iRX_FIFO_Empty_0\;
    iRX_FIFO_Full_0 <= \iRX_FIFO_Full_0\;
    fifo_MEMRE <= \fifo_MEMRE\;
    fifo_MEMWE <= \fifo_MEMWE\;

    \rptr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[4]_net_1\, S
         => \rptr_s[5]\, Y => OPEN, FCO => \rptr_cry[5]_net_1\);
    
    \memwaddr_r_2[9]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_9_S_0, D => un4_we_i_9, Y => 
        \memwaddr_r_2[9]_net_1\);
    
    wdiff_bus_cry_8 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[8]_net_1\, B => 
        \rptr_bin_sync2[8]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_7\, S => \wdiff_bus[8]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_8\);
    
    \wptr_bin_sync2[12]\ : SLE
      port map(D => \wptr_bin_sync[12]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[12]_net_1\);
    
    wdiff_bus_cry_11 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[11]_net_1\, B => 
        \rptr_bin_sync2[11]_net_1\, C => GND_net_1, D => 
        GND_net_1, FCI => \wdiff_bus_cry_10\, S => 
        \wdiff_bus[11]\, Y => OPEN, FCO => \wdiff_bus_cry_11\);
    
    \wptr_gray[4]\ : SLE
      port map(D => \wptr_gray_1[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[4]_net_1\);
    
    \rptr_gray_1[3]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[3]_net_1\, B => \rptr[4]_net_1\, Y => 
        \rptr_gray_1[3]_net_1\);
    
    wptr_s_907 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => wptr_s_907_FCO);
    
    \rptr_bin_sync2[6]\ : SLE
      port map(D => bin_N_4_0_i, CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_bin_sync2[6]_net_1\);
    
    \rptr[1]\ : SLE
      port map(D => \rptr_s[1]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[1]_net_1\);
    
    \wptr_gray_1[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[9]_net_1\, B => \wptr[10]_net_1\, Y => 
        \wptr_gray_1[9]_net_1\);
    
    \rptr_gray_1[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[5]_net_1\, B => \rptr[6]_net_1\, Y => 
        \rptr_gray_1[5]_net_1\);
    
    \rptr_gray[9]\ : SLE
      port map(D => \rptr_gray_1[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[9]_net_1\);
    
    un1_memwaddr_r_cry_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_6\, 
        S => un1_memwaddr_r_cry_7_S_0, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_7\);
    
    \rptr_gray[8]\ : SLE
      port map(D => \rptr_gray_1[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[8]_net_1\);
    
    un1_memraddr_r_cry_11 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[11]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_10\, 
        S => un1_memraddr_r_cry_11_S_0, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_11\);
    
    \rptr_gray_1[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[2]_net_1\, B => \rptr[3]_net_1\, Y => 
        \rptr_gray_1[2]_net_1\);
    
    \rptr_bin_sync2[7]\ : SLE
      port map(D => \rptr_bin_sync[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[7]_net_1\);
    
    \memwaddr_r[1]\ : SLE
      port map(D => un1_memwaddr_r_cry_1_S_0, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[1]\);
    
    \wptr_gray_1[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[7]_net_1\, B => \wptr[8]_net_1\, Y => 
        \wptr_gray_1[7]_net_1\);
    
    \rptr_gray[13]\ : SLE
      port map(D => \rptr[13]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[13]_net_1\);
    
    \memraddr_r[0]\ : SLE
      port map(D => \fifo_MEMRADDR_i[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[0]\);
    
    \memraddr_r_2[9]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => 
        un1_memraddr_r_cry_9_S_0, D => un4_re_i_9, Y => 
        \memraddr_r_2[9]_net_1\);
    
    \wptr[0]\ : SLE
      port map(D => \wptr_s[0]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[0]_net_1\);
    
    \rptr_bin_sync2[8]\ : SLE
      port map(D => \rptr_bin_sync[8]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[8]_net_1\);
    
    \rptr_gray_1[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[1]_net_1\, B => \rptr[2]_net_1\, Y => 
        \rptr_gray_1[1]_net_1\);
    
    \rptr_gray[10]\ : SLE
      port map(D => \rptr_gray_1[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[10]_net_1\);
    
    \wptr_gray_1[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[0]_net_1\, B => \wptr[1]_net_1\, Y => 
        \wptr_gray_1[0]_net_1\);
    
    wdiff_bus_cry_9 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[9]_net_1\, B => 
        \rptr_bin_sync2[9]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_8\, S => \wdiff_bus[9]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_9\);
    
    \rptr[5]\ : SLE
      port map(D => \rptr_s[5]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[5]_net_1\);
    
    \rptr_gray[3]\ : SLE
      port map(D => \rptr_gray_1[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[3]_net_1\);
    
    \rptr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[5]_net_1\, S
         => \rptr_s[6]\, Y => OPEN, FCO => \rptr_cry[6]_net_1\);
    
    \wptr_gray[3]\ : SLE
      port map(D => \wptr_gray_1[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[3]_net_1\);
    
    \rptr_gray_1[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[10]_net_1\, B => \rptr[11]_net_1\, Y
         => \rptr_gray_1[10]_net_1\);
    
    un1_memraddr_r_cry_10 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_9\, 
        S => un1_memraddr_r_cry_10_S_0, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_10\);
    
    \rptr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[7]_net_1\, S
         => \rptr_s[8]\, Y => OPEN, FCO => \rptr_cry[8]_net_1\);
    
    \rptr[7]\ : SLE
      port map(D => \rptr_s[7]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[7]_net_1\);
    
    rdiff_bus_cry_4 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[4]_net_1\, B => 
        \rptr[4]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_3\, S => \rdiff_bus[4]\, Y => OPEN, FCO
         => \rdiff_bus_cry_4\);
    
    \rptr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[9]_net_1\, S
         => \rptr_s[10]\, Y => OPEN, FCO => \rptr_cry[10]_net_1\);
    
    \rptr_bin_sync2[12]\ : SLE
      port map(D => \rptr_bin_sync[12]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[12]_net_1\);
    
    memwe_0_a3 : CFG3
      generic map(INIT => x"20")

      port map(A => RX_FIFO_TxColDetDis_wr_en, B => 
        \iRX_FIFO_Full_0\, C => iRX_FIFO_wr_en_0_0, Y => 
        \fifo_MEMWE\);
    
    \rptr_bin_sync2[0]\ : SLE
      port map(D => \rptr_bin_sync[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[0]_net_1\);
    
    \L1.empty_r_3_0_a2_7\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \rdiff_bus[1]\, B => \rdiff_bus[4]\, C => 
        \rdiff_bus[3]\, D => \rdiff_bus[2]\, Y => 
        empty_r_3_0_a2_7);
    
    \wptr[11]\ : SLE
      port map(D => \wptr_s[11]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[11]_net_1\);
    
    rdiff_bus_cry_1 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[1]_net_1\, B => 
        \rptr[1]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_0\, S => \rdiff_bus[1]\, Y => OPEN, FCO
         => \rdiff_bus_cry_1\);
    
    \memraddr_r[1]\ : SLE
      port map(D => un1_memraddr_r_cry_1_S_0, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[1]\);
    
    \L1.empty_r_3_0_a2_9\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \rdiff_bus[9]\, B => \rdiff_bus[10]\, C => 
        \rdiff_bus[11]\, D => \rdiff_bus[12]\, Y => 
        empty_r_3_0_a2_9);
    
    \rptr_bin_sync2[2]\ : SLE
      port map(D => \rptr_bin_sync[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[2]_net_1\);
    
    \memraddr_r_2[7]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => 
        un1_memraddr_r_cry_7_S_0, D => un4_re_i_9, Y => 
        \memraddr_r_2[7]_net_1\);
    
    un1_memwaddr_r_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_5\, 
        S => un1_memwaddr_r_cry_6_S_0, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_6\);
    
    rdiff_bus_cry_6 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[6]_net_1\, B => 
        \rptr[6]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_5\, S => \rdiff_bus[6]\, Y => OPEN, FCO
         => \rdiff_bus_cry_6\);
    
    \memwaddr_r_2[10]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_10_S_0, D => un4_we_i_9, Y => 
        \memwaddr_r_2[10]_net_1\);
    
    \memraddr_r_2[5]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => 
        un1_memraddr_r_cry_5_S_0, D => un4_re_i_9, Y => 
        \memraddr_r_2[5]_net_1\);
    
    un1_memraddr_r_s_1_925 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[0]\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => un1_memraddr_r_s_1_925_FCO);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    un1_memwaddr_r_cry_9 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[9]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_8\, 
        S => un1_memwaddr_r_cry_9_S_0, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_9\);
    
    \rptr_gray[1]\ : SLE
      port map(D => \rptr_gray_1[1]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[1]_net_1\);
    
    \memwaddr_r[7]\ : SLE
      port map(D => \memwaddr_r_2[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[7]\);
    
    \wptr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[3]_net_1\, S
         => \wptr_s[4]\, Y => OPEN, FCO => \wptr_cry[4]_net_1\);
    
    \wptr_gray_1[12]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[13]_net_1\, B => \wptr[12]_net_1\, Y
         => \wptr_gray_1[12]_net_1\);
    
    \wptr[12]\ : SLE
      port map(D => \wptr_s[12]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[12]_net_1\);
    
    \wptr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[9]_net_1\, S
         => \wptr_s[10]\, Y => OPEN, FCO => \wptr_cry[10]_net_1\);
    
    wdiff_bus_cry_5 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[5]_net_1\, B => 
        \rptr_bin_sync2[5]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_4\, S => \wdiff_bus[5]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_5\);
    
    \rptr_gray[12]\ : SLE
      port map(D => \rptr_gray_1[12]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[12]_net_1\);
    
    \memwaddr_r[4]\ : SLE
      port map(D => un1_memwaddr_r_cry_4_S_0, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[4]\);
    
    \wptr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[1]_net_1\, S
         => \wptr_s[2]\, Y => OPEN, FCO => \wptr_cry[2]_net_1\);
    
    \memraddr_r_2[10]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => 
        un1_memraddr_r_cry_10_S_0, D => un4_re_i_9, Y => 
        \memraddr_r_2[10]_net_1\);
    
    rdiff_bus_cry_11 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[11]_net_1\, B => 
        \rptr[11]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_10\, S => \rdiff_bus[11]\, Y => OPEN, FCO
         => \rdiff_bus_cry_11\);
    
    wdiff_bus_cry_0 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[0]_net_1\, B => 
        \rptr_bin_sync2[0]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => VCC_net_1, S => OPEN, Y => wdiff_bus_cry_0_Y_1, 
        FCO => \wdiff_bus_cry_0\);
    
    \wptr[1]\ : SLE
      port map(D => \wptr_s[1]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[1]_net_1\);
    
    \rptr_bin_sync2[4]\ : SLE
      port map(D => bin_N_6_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[4]_net_1\);
    
    \wptr_bin_sync2[6]\ : SLE
      port map(D => \wptr_bin_sync[6]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[6]_net_1\);
    
    \rptr[3]\ : SLE
      port map(D => \rptr_s[3]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[3]_net_1\);
    
    fulli_0_a3_4_3 : CFG4
      generic map(INIT => x"8000")

      port map(A => \wdiff_bus[7]\, B => \wdiff_bus[8]\, C => 
        \wdiff_bus[9]\, D => \wdiff_bus[10]\, Y => 
        \fulli_0_a3_4_3\);
    
    \wptr_gray[13]\ : SLE
      port map(D => \wptr[13]_net_1\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr_gray[13]_net_1\);
    
    \wptr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[2]_net_1\, S
         => \wptr_s[3]\, Y => OPEN, FCO => \wptr_cry[3]_net_1\);
    
    \L1.empty_r_3_0_a2_8\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \rdiff_bus[5]\, B => \rdiff_bus[6]\, C => 
        \rdiff_bus[7]\, D => \rdiff_bus[8]\, Y => 
        empty_r_3_0_a2_8);
    
    \rptr[6]\ : SLE
      port map(D => \rptr_s[6]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[6]_net_1\);
    
    rdiff_bus_cry_8 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[8]_net_1\, B => 
        \rptr[8]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_7\, S => \rdiff_bus[8]\, Y => OPEN, FCO
         => \rdiff_bus_cry_8\);
    
    \wptr_gray[10]\ : SLE
      port map(D => \wptr_gray_1[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[10]_net_1\);
    
    rdiff_bus_cry_7 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[7]_net_1\, B => 
        \rptr[7]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_6\, S => \rdiff_bus[7]\, Y => OPEN, FCO
         => \rdiff_bus_cry_7\);
    
    \wptr_bin_sync2[7]\ : SLE
      port map(D => \wptr_bin_sync[7]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[7]_net_1\);
    
    \rptr_gray_1[11]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[11]_net_1\, B => \rptr[12]_net_1\, Y
         => \rptr_gray_1[11]_net_1\);
    
    \rptr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[8]_net_1\, S
         => \rptr_s[9]\, Y => OPEN, FCO => \rptr_cry[9]_net_1\);
    
    un1_memwaddr_r_cry_1 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[1]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        un1_memwaddr_r_s_1_926_FCO, S => un1_memwaddr_r_cry_1_S_0, 
        Y => OPEN, FCO => \un1_memwaddr_r_cry_1\);
    
    \rptr_gray[5]\ : SLE
      port map(D => \rptr_gray_1[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[5]_net_1\);
    
    un1_memwaddr_r_s_12 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[12]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_11\, 
        S => un1_memwaddr_r_s_12_S_0, Y => OPEN, FCO => OPEN);
    
    \wptr_gray_1[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[2]_net_1\, B => \wptr[3]_net_1\, Y => 
        \wptr_gray_1[2]_net_1\);
    
    \wptr[5]\ : SLE
      port map(D => \wptr_s[5]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[5]_net_1\);
    
    rdiff_bus_cry_5 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[5]_net_1\, B => 
        \rptr[5]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_4\, S => \rdiff_bus[5]\, Y => OPEN, FCO
         => \rdiff_bus_cry_5\);
    
    \wptr_bin_sync2[8]\ : SLE
      port map(D => \wptr_bin_sync[8]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[8]_net_1\);
    
    \wptr[7]\ : SLE
      port map(D => \wptr_s[7]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[7]_net_1\);
    
    un1_memwaddr_r_cry_2 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[2]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_1\, 
        S => un1_memwaddr_r_cry_2_S_0, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_2\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \wptr_gray[1]\ : SLE
      port map(D => \wptr_gray_1[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[1]_net_1\);
    
    \rptr_gray_1[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[9]_net_1\, B => \rptr[10]_net_1\, Y => 
        \rptr_gray_1[9]_net_1\);
    
    \rptr_bin_sync2[5]\ : SLE
      port map(D => \rptr_bin_sync[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[5]_net_1\);
    
    \rptr_bin_sync2[1]\ : SLE
      port map(D => \rptr_bin_sync[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[1]_net_1\);
    
    \memwaddr_r[10]\ : SLE
      port map(D => \memwaddr_r_2[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[10]\);
    
    wdiff_bus_cry_7 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[7]_net_1\, B => 
        \rptr_bin_sync2[7]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_6\, S => \wdiff_bus[7]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_7\);
    
    \wptr_bin_sync2[0]\ : SLE
      port map(D => \wptr_bin_sync[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rdiff_bus);
    
    un1_memwaddr_r_cry_8 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[8]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_7\, 
        S => un1_memwaddr_r_cry_8_S_0, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_8\);
    
    \wptr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => wptr_s_907_FCO, S => 
        \wptr_s[1]\, Y => OPEN, FCO => \wptr_cry[1]_net_1\);
    
    un1_memwaddr_r_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_3\, 
        S => un1_memwaddr_r_cry_4_S_0, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_4\);
    
    un1_memwaddr_r_cry_3 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[3]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_2\, 
        S => un1_memwaddr_r_cry_3_S_0, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_3\);
    
    \memraddr_r[8]\ : SLE
      port map(D => \memraddr_r_2[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[8]\);
    
    \rptr[9]\ : SLE
      port map(D => \rptr_s[9]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[9]_net_1\);
    
    \wptr_gray_1[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[6]_net_1\, B => \wptr[7]_net_1\, Y => 
        \wptr_gray_1[6]_net_1\);
    
    \wptr_gray[12]\ : SLE
      port map(D => \wptr_gray_1[12]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[12]_net_1\);
    
    \wptr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[6]_net_1\, S
         => \wptr_s[7]\, Y => OPEN, FCO => \wptr_cry[7]_net_1\);
    
    \wptr_bin_sync2[2]\ : SLE
      port map(D => \wptr_bin_sync[2]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[2]_net_1\);
    
    \L1.un4_re_i_9\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \fifo_MEMRADDR[4]\, B => \fifo_MEMRADDR[3]\, 
        C => \fifo_MEMRADDR[0]\, D => un4_re_i_0, Y => un4_re_i_9);
    
    un1_memraddr_r_cry_3 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[3]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_2\, 
        S => un1_memraddr_r_cry_3_S_0, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_3\);
    
    \rptr_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \rptr[0]_net_1\, Y => \rptr_s[0]\);
    
    un1_memraddr_r_cry_1 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[1]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        un1_memraddr_r_s_1_925_FCO, S => un1_memraddr_r_cry_1_S_0, 
        Y => OPEN, FCO => \un1_memraddr_r_cry_1\);
    
    \rptr[4]\ : SLE
      port map(D => \rptr_s[4]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[4]_net_1\);
    
    \memwaddr_r_2[5]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_5_S_0, D => un4_we_i_9, Y => 
        \memwaddr_r_2[5]_net_1\);
    
    \wptr_gray[6]\ : SLE
      port map(D => \wptr_gray_1[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[6]_net_1\);
    
    \wptr_gray_1[3]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[3]_net_1\, B => \wptr[4]_net_1\, Y => 
        \wptr_gray_1[3]_net_1\);
    
    \wptr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[4]_net_1\, S
         => \wptr_s[5]\, Y => OPEN, FCO => \wptr_cry[5]_net_1\);
    
    un1_memraddr_r_cry_9 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[9]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_8\, 
        S => un1_memraddr_r_cry_9_S_0, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_9\);
    
    fulli_0_a3_5_1 : CFG4
      generic map(INIT => x"0F1F")

      port map(A => \wdiff_bus[5]\, B => \wdiff_bus[6]\, C => 
        \fulli_0_a3_4_3\, D => \fulli_0_a3_d_4\, Y => 
        \fulli_0_a3_5_1\);
    
    \rptr_gray[4]\ : SLE
      port map(D => \rptr_gray_1[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[4]_net_1\);
    
    un1_memraddr_r_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_4\, 
        S => un1_memraddr_r_cry_5_S_0, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_5\);
    
    \wptr_bin_sync2[4]\ : SLE
      port map(D => \wptr_bin_sync[4]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[4]_net_1\);
    
    \L1.empty_r_3_0_a2_6\ : CFG3
      generic map(INIT => x"0E")

      port map(A => iRX_FIFO_rd_en_0, B => rdiff_bus_cry_0_Y_1, C
         => \rdiff_bus[13]\, Y => empty_r_3_0_a2_6);
    
    \wptr[3]\ : SLE
      port map(D => \wptr_s[3]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[3]_net_1\);
    
    \L1.un4_we_i_9\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \fifo_MEMWADDR[4]\, B => \fifo_MEMWADDR[3]\, 
        C => \fifo_MEMWADDR[0]\, D => un4_we_i_0, Y => un4_we_i_9);
    
    \memwaddr_r[6]\ : SLE
      port map(D => un1_memwaddr_r_cry_6_S_0, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[6]\);
    
    \wptr[6]\ : SLE
      port map(D => \wptr_s[6]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[6]_net_1\);
    
    \memwaddr_r[9]\ : SLE
      port map(D => \memwaddr_r_2[9]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[9]\);
    
    \memraddr_r[10]\ : SLE
      port map(D => \memraddr_r_2[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[10]\);
    
    \L1.un4_re_i_8\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \fifo_MEMRADDR[10]\, B => \fifo_MEMRADDR[9]\, 
        C => \fifo_MEMRADDR[8]\, D => \fifo_MEMRADDR[7]\, Y => 
        un4_re_i_8);
    
    \memwaddr_r[3]\ : SLE
      port map(D => un1_memwaddr_r_cry_3_S_0, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[3]\);
    
    \rptr_gray_1[12]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[13]_net_1\, B => \rptr[12]_net_1\, Y
         => \rptr_gray_1[12]_net_1\);
    
    full_r : SLE
      port map(D => fulli, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \iRX_FIFO_Full_0\);
    
    \rptr_bin_sync2[3]\ : SLE
      port map(D => \rptr_bin_sync[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[3]_net_1\);
    
    un1_memwaddr_r_s_1_926 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[0]\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => un1_memwaddr_r_s_1_926_FCO);
    
    \wptr_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \wptr[0]_net_1\, Y => \wptr_s[0]\);
    
    \rptr[2]\ : SLE
      port map(D => \rptr_s[2]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[2]_net_1\);
    
    \memraddr_r[3]\ : SLE
      port map(D => un1_memraddr_r_cry_3_S_0, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[3]\);
    
    \wptr[13]\ : SLE
      port map(D => \wptr_s[13]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \wptr[13]_net_1\);
    
    \rptr_bin_sync2[9]\ : SLE
      port map(D => \rptr_bin_sync[9]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[9]_net_1\);
    
    \wptr_bin_sync2[13]\ : SLE
      port map(D => \wptr_bin_sync[13]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[13]_net_1\);
    
    \rptr[11]\ : SLE
      port map(D => \rptr_s[11]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rptr[11]_net_1\);
    
    \wptr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[5]_net_1\, S
         => \wptr_s[6]\, Y => OPEN, FCO => \wptr_cry[6]_net_1\);
    
    \rptr_bin_sync2[11]\ : SLE
      port map(D => \rptr_bin_sync[11]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[11]_net_1\);
    
    \wptr_bin_sync2[5]\ : SLE
      port map(D => \wptr_bin_sync[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[5]_net_1\);
    
    \L1.un4_we_i_8\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \fifo_MEMWADDR[10]\, B => \fifo_MEMWADDR[9]\, 
        C => \fifo_MEMWADDR[8]\, D => \fifo_MEMWADDR[7]\, Y => 
        un4_we_i_8);
    
    \wptr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[7]_net_1\, S
         => \wptr_s[8]\, Y => OPEN, FCO => \wptr_cry[8]_net_1\);
    
    \wptr_bin_sync2[1]\ : SLE
      port map(D => \wptr_bin_sync[1]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[1]_net_1\);
    
    Wr_corefifo_grayToBinConv : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_2
      port map(wptr_bin_sync(13) => \wptr_bin_sync[13]\, 
        wptr_bin_sync(12) => \wptr_bin_sync[12]\, 
        wptr_bin_sync(11) => \wptr_bin_sync[11]\, 
        wptr_bin_sync(10) => \wptr_bin_sync[10]\, 
        wptr_bin_sync(9) => \wptr_bin_sync[9]\, wptr_bin_sync(8)
         => \wptr_bin_sync[8]\, wptr_bin_sync(7) => 
        \wptr_bin_sync[7]\, wptr_bin_sync(6) => 
        \wptr_bin_sync[6]\, wptr_bin_sync(5) => 
        \wptr_bin_sync[5]\, wptr_bin_sync(4) => 
        \wptr_bin_sync[4]\, wptr_bin_sync(3) => 
        \wptr_bin_sync[3]\, wptr_bin_sync(2) => 
        \wptr_bin_sync[2]\, wptr_bin_sync(1) => 
        \wptr_bin_sync[1]\, wptr_bin_sync(0) => 
        \wptr_bin_sync[0]\, wptr_gray_sync(12) => 
        \wptr_gray_sync[12]\, wptr_gray_sync(11) => 
        \wptr_gray_sync[11]\, wptr_gray_sync(10) => 
        \wptr_gray_sync[10]\, wptr_gray_sync(9) => 
        \wptr_gray_sync[9]\, wptr_gray_sync(8) => 
        \wptr_gray_sync[8]\, wptr_gray_sync(7) => 
        \wptr_gray_sync[7]\, wptr_gray_sync(6) => 
        \wptr_gray_sync[6]\, wptr_gray_sync(5) => 
        \wptr_gray_sync[5]\, wptr_gray_sync(4) => 
        \wptr_gray_sync[4]\, wptr_gray_sync(3) => 
        \wptr_gray_sync[3]\, wptr_gray_sync(2) => 
        \wptr_gray_sync[2]\, wptr_gray_sync(1) => 
        \wptr_gray_sync[1]\, wptr_gray_sync(0) => 
        \wptr_gray_sync[0]\);
    
    \wptr_gray_1[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[4]_net_1\, B => \wptr[5]_net_1\, Y => 
        \wptr_gray_1[4]_net_1\);
    
    \rptr_bin_sync2[13]\ : SLE
      port map(D => \rptr_bin_sync[13]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[13]_net_1\);
    
    \L1.un4_re_i_7\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \fifo_MEMRADDR[12]\, B => \fifo_MEMRADDR[11]\, 
        C => \fifo_MEMRADDR[6]\, D => \fifo_MEMRADDR[5]\, Y => 
        un4_re_i_7);
    
    overflow_r : SLE
      port map(D => N_6_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        iRX_FIFO_OVERFLOW_0);
    
    \memraddr_r_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \fifo_MEMRADDR[0]\, Y => \fifo_MEMRADDR_i[0]\);
    
    \memraddr_r_2[8]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => 
        un1_memraddr_r_cry_8_S_0, D => un4_re_i_9, Y => 
        \memraddr_r_2[8]_net_1\);
    
    \rptr_gray[11]\ : SLE
      port map(D => \rptr_gray_1[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[11]_net_1\);
    
    \wptr_bin_sync2[10]\ : SLE
      port map(D => \wptr_bin_sync[10]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[10]_net_1\);
    
    \rptr[10]\ : SLE
      port map(D => \rptr_s[10]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rptr[10]_net_1\);
    
    \wptr[9]\ : SLE
      port map(D => \wptr_s[9]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[9]_net_1\);
    
    Wr_corefifo_doubleSync : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_1
      port map(wptr_gray(13) => \wptr_gray[13]_net_1\, 
        wptr_gray(12) => \wptr_gray[12]_net_1\, wptr_gray(11) => 
        \wptr_gray[11]_net_1\, wptr_gray(10) => 
        \wptr_gray[10]_net_1\, wptr_gray(9) => 
        \wptr_gray[9]_net_1\, wptr_gray(8) => 
        \wptr_gray[8]_net_1\, wptr_gray(7) => 
        \wptr_gray[7]_net_1\, wptr_gray(6) => 
        \wptr_gray[6]_net_1\, wptr_gray(5) => 
        \wptr_gray[5]_net_1\, wptr_gray(4) => 
        \wptr_gray[4]_net_1\, wptr_gray(3) => 
        \wptr_gray[3]_net_1\, wptr_gray(2) => 
        \wptr_gray[2]_net_1\, wptr_gray(1) => 
        \wptr_gray[1]_net_1\, wptr_gray(0) => 
        \wptr_gray[0]_net_1\, wptr_gray_sync(12) => 
        \wptr_gray_sync[12]\, wptr_gray_sync(11) => 
        \wptr_gray_sync[11]\, wptr_gray_sync(10) => 
        \wptr_gray_sync[10]\, wptr_gray_sync(9) => 
        \wptr_gray_sync[9]\, wptr_gray_sync(8) => 
        \wptr_gray_sync[8]\, wptr_gray_sync(7) => 
        \wptr_gray_sync[7]\, wptr_gray_sync(6) => 
        \wptr_gray_sync[6]\, wptr_gray_sync(5) => 
        \wptr_gray_sync[5]\, wptr_gray_sync(4) => 
        \wptr_gray_sync[4]\, wptr_gray_sync(3) => 
        \wptr_gray_sync[3]\, wptr_gray_sync(2) => 
        \wptr_gray_sync[2]\, wptr_gray_sync(1) => 
        \wptr_gray_sync[1]\, wptr_gray_sync(0) => 
        \wptr_gray_sync[0]\, wptr_bin_sync_0 => 
        \wptr_bin_sync[13]\, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, irx_fifo_rst_i => 
        irx_fifo_rst_i);
    
    un1_memwaddr_r_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_4\, 
        S => un1_memwaddr_r_cry_5_S_0, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_5\);
    
    \rptr_gray[0]\ : SLE
      port map(D => \rptr_gray_1[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[0]_net_1\);
    
    empty_r : SLE
      port map(D => empty_r_3, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \iRX_FIFO_Empty_0\);
    
    \memwaddr_r_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \fifo_MEMWADDR[0]\, Y => \fifo_MEMWADDR_i[0]\);
    
    \memwaddr_r_2[12]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_s_12_S_0, D => un4_we_i_9, Y => 
        \memwaddr_r_2[12]_net_1\);
    
    \rptr_gray_1[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[7]_net_1\, B => \rptr[8]_net_1\, Y => 
        \rptr_gray_1[7]_net_1\);
    
    fulli_0_a3_5 : CFG4
      generic map(INIT => x"BAAA")

      port map(A => \wdiff_bus[13]\, B => \fulli_0_a3_5_1\, C => 
        \wdiff_bus[11]\, D => \wdiff_bus[12]\, Y => fulli);
    
    un1_memraddr_r_cry_2 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[2]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_1\, 
        S => un1_memraddr_r_cry_2_S_0, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_2\);
    
    wdiff_bus_cry_12 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[12]_net_1\, B => 
        \rptr_bin_sync2[12]_net_1\, C => GND_net_1, D => 
        GND_net_1, FCI => \wdiff_bus_cry_11\, S => 
        \wdiff_bus[12]\, Y => OPEN, FCO => \wdiff_bus_cry_12\);
    
    \wptr[4]\ : SLE
      port map(D => \wptr_s[4]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[4]_net_1\);
    
    un1_memraddr_r_cry_8 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[8]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_7\, 
        S => un1_memraddr_r_cry_8_S_0, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_8\);
    
    \rptr_s[13]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[13]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[12]_net_1\, S
         => \rptr_s[13]_net_1\, Y => OPEN, FCO => OPEN);
    
    \memwaddr_r[8]\ : SLE
      port map(D => \memwaddr_r_2[8]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[8]\);
    
    \memwaddr_r[2]\ : SLE
      port map(D => un1_memwaddr_r_cry_2_S_0, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[2]\);
    
    \wptr_bin_sync2[11]\ : SLE
      port map(D => \wptr_bin_sync[11]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[11]_net_1\);
    
    \L1.un4_we_i_7\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \fifo_MEMWADDR[12]\, B => \fifo_MEMWADDR[11]\, 
        C => \fifo_MEMWADDR[6]\, D => \fifo_MEMWADDR[5]\, Y => 
        un4_we_i_7);
    
    \wptr_gray_1[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[1]_net_1\, B => \wptr[2]_net_1\, Y => 
        \wptr_gray_1[1]_net_1\);
    
    underflow_r : SLE
      port map(D => N_5_i, CLK => m2s010_som_sb_0_CCC_71MHz, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => iRX_FIFO_UNDERRUN_0);
    
    \memwaddr_r_2[11]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_11_S_0, D => un4_we_i_9, Y => 
        \memwaddr_r_2[11]_net_1\);
    
    \memraddr_r_2[12]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => 
        un1_memraddr_r_s_12_S_0, D => un4_re_i_9, Y => 
        \memraddr_r_2[12]_net_1\);
    
    \wptr_gray[5]\ : SLE
      port map(D => \wptr_gray_1[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[5]_net_1\);
    
    overflow_r_RNO : CFG3
      generic map(INIT => x"80")

      port map(A => RX_FIFO_TxColDetDis_wr_en, B => 
        \iRX_FIFO_Full_0\, C => iRX_FIFO_wr_en_0_0, Y => N_6_i);
    
    \memraddr_r[7]\ : SLE
      port map(D => \memraddr_r_2[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[7]\);
    
    un1_memraddr_r_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_5\, 
        S => un1_memraddr_r_cry_6_S_0, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_6\);
    
    \rptr_bin_sync2[10]\ : SLE
      port map(D => \rptr_bin_sync[10]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[10]_net_1\);
    
    wdiff_bus_s_13 : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \rptr_bin_sync2[13]_net_1\, C
         => \wptr[13]_net_1\, D => GND_net_1, FCI => 
        \wdiff_bus_cry_12\, S => \wdiff_bus[13]\, Y => OPEN, FCO
         => OPEN);
    
    wdiff_bus_cry_10 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[10]_net_1\, B => 
        \rptr_bin_sync2[10]_net_1\, C => GND_net_1, D => 
        GND_net_1, FCI => \wdiff_bus_cry_9\, S => \wdiff_bus[10]\, 
        Y => OPEN, FCO => \wdiff_bus_cry_10\);
    
    \memwaddr_r[11]\ : SLE
      port map(D => \memwaddr_r_2[11]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[11]\);
    
    \wptr_gray[8]\ : SLE
      port map(D => \wptr_gray_1[8]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[8]_net_1\);
    
    \memraddr_r_2[11]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => 
        un1_memraddr_r_cry_11_S_0, D => un4_re_i_9, Y => 
        \memraddr_r_2[11]_net_1\);
    
    un1_memraddr_r_s_12 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[12]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_11\, 
        S => un1_memraddr_r_s_12_S_0, Y => OPEN, FCO => OPEN);
    
    \wptr_gray[7]\ : SLE
      port map(D => \wptr_gray_1[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[7]_net_1\);
    
    \wptr_gray_1[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[5]_net_1\, B => \wptr[6]_net_1\, Y => 
        \wptr_gray_1[5]_net_1\);
    
    \memwaddr_r[5]\ : SLE
      port map(D => \memwaddr_r_2[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[5]\);
    
    \L1.empty_r_3_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => empty_r_3_0_a2_6, B => empty_r_3_0_a2_7, C
         => empty_r_3_0_a2_9, D => empty_r_3_0_a2_8, Y => 
        empty_r_3);
    
    un1_memraddr_r_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_3\, 
        S => un1_memraddr_r_cry_4_S_0, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_4\);
    
    \rptr[8]\ : SLE
      port map(D => \rptr_s[8]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[8]_net_1\);
    
    Rd_corefifo_doubleSync : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_0
      port map(rptr_gray(13) => \rptr_gray[13]_net_1\, 
        rptr_gray(12) => \rptr_gray[12]_net_1\, rptr_gray(11) => 
        \rptr_gray[11]_net_1\, rptr_gray(10) => 
        \rptr_gray[10]_net_1\, rptr_gray(9) => 
        \rptr_gray[9]_net_1\, rptr_gray(8) => 
        \rptr_gray[8]_net_1\, rptr_gray(7) => 
        \rptr_gray[7]_net_1\, rptr_gray(6) => 
        \rptr_gray[6]_net_1\, rptr_gray(5) => 
        \rptr_gray[5]_net_1\, rptr_gray(4) => 
        \rptr_gray[4]_net_1\, rptr_gray(3) => 
        \rptr_gray[3]_net_1\, rptr_gray(2) => 
        \rptr_gray[2]_net_1\, rptr_gray(1) => 
        \rptr_gray[1]_net_1\, rptr_gray(0) => 
        \rptr_gray[0]_net_1\, rptr_gray_sync(12) => 
        \rptr_gray_sync[12]\, rptr_gray_sync(11) => 
        \rptr_gray_sync[11]\, rptr_gray_sync(10) => 
        \rptr_gray_sync[10]\, rptr_gray_sync(9) => 
        \rptr_gray_sync[9]\, rptr_gray_sync(8) => 
        \rptr_gray_sync[8]\, rptr_gray_sync(7) => 
        \rptr_gray_sync[7]\, rptr_gray_sync(6) => 
        \rptr_gray_sync[6]\, rptr_gray_sync(5) => 
        \rptr_gray_sync[5]\, rptr_gray_sync(4) => 
        \rptr_gray_sync[4]\, rptr_gray_sync(3) => 
        \rptr_gray_sync[3]\, rptr_gray_sync(2) => 
        \rptr_gray_sync[2]\, rptr_gray_sync(1) => 
        \rptr_gray_sync[1]\, rptr_gray_sync(0) => 
        \rptr_gray_sync[0]\, rptr_bin_sync_0 => 
        \rptr_bin_sync[13]\, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, irx_fifo_rst_i => irx_fifo_rst_i);
    
    underflow_r_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => iRX_FIFO_rd_en_0, B => \iRX_FIFO_Empty_0\, Y
         => N_5_i);
    
    \rptr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[3]_net_1\, S
         => \rptr_s[4]\, Y => OPEN, FCO => \rptr_cry[4]_net_1\);
    
    wdiff_bus_cry_2 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[2]_net_1\, B => 
        \rptr_bin_sync2[2]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_1\, S => \wdiff_bus[2]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_2\);
    
    \rptr_gray[2]\ : SLE
      port map(D => \rptr_gray_1[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[2]_net_1\);
    
    \wptr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[8]_net_1\, S
         => \wptr_s[9]\, Y => OPEN, FCO => \wptr_cry[9]_net_1\);
    
    \wptr_bin_sync2[3]\ : SLE
      port map(D => \wptr_bin_sync[3]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[3]_net_1\);
    
    \rptr[12]\ : SLE
      port map(D => \rptr_s[12]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rptr[12]_net_1\);
    
    fulli_0_a3_d_4 : CFG4
      generic map(INIT => x"4000")

      port map(A => wdiff_bus_cry_0_Y_1, B => \wdiff_bus[1]\, C
         => \wdiff_bus[4]\, D => \fulli_0_a3_d_3\, Y => 
        \fulli_0_a3_d_4\);
    
    \wptr[2]\ : SLE
      port map(D => \wptr_s[2]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[2]_net_1\);
    
    \rptr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[1]_net_1\, S
         => \rptr_s[2]\, Y => OPEN, FCO => \rptr_cry[2]_net_1\);
    
    rdiff_bus_cry_9 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[9]_net_1\, B => 
        \rptr[9]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_8\, S => \rdiff_bus[9]\, Y => OPEN, FCO
         => \rdiff_bus_cry_9\);
    
    \memwaddr_r[0]\ : SLE
      port map(D => \fifo_MEMWADDR_i[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[0]\);
    
    fulli_0_a3_d_3 : CFG4
      generic map(INIT => x"8000")

      port map(A => \wdiff_bus[2]\, B => 
        RX_FIFO_TxColDetDis_wr_en, C => iRX_FIFO_wr_en_0_0, D => 
        \wdiff_bus[3]\, Y => \fulli_0_a3_d_3\);
    
    \wptr_gray[2]\ : SLE
      port map(D => \wptr_gray_1[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[2]_net_1\);
    
    \wptr_cry[12]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[12]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[11]_net_1\, S
         => \wptr_s[12]\, Y => OPEN, FCO => \wptr_cry[12]_net_1\);
    
    \memwaddr_r_2[7]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_7_S_0, D => un4_we_i_9, Y => 
        \memwaddr_r_2[7]_net_1\);
    
    wdiff_bus_cry_4 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[4]_net_1\, B => 
        \rptr_bin_sync2[4]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_3\, S => \wdiff_bus[4]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_4\);
    
    un1_memraddr_r_cry_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_6\, 
        S => un1_memraddr_r_cry_7_S_0, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_7\);
    
    \wptr_s[13]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[13]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[12]_net_1\, S
         => \wptr_s[13]_net_1\, Y => OPEN, FCO => OPEN);
    
    \wptr_gray[11]\ : SLE
      port map(D => \wptr_gray_1[11]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[11]_net_1\);
    
    \wptr_bin_sync2[9]\ : SLE
      port map(D => \wptr_bin_sync[9]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[9]_net_1\);
    
    rptr_s_906 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => rptr_s_906_FCO);
    
    \rptr_gray_1[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[6]_net_1\, B => \rptr[7]_net_1\, Y => 
        \rptr_gray_1[6]_net_1\);
    
    \wptr_gray_1[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[10]_net_1\, B => \wptr[11]_net_1\, Y
         => \wptr_gray_1[10]_net_1\);
    
    wdiff_bus_cry_6 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[6]_net_1\, B => 
        \rptr_bin_sync2[6]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_5\, S => \wdiff_bus[6]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_6\);
    
    \rptr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[2]_net_1\, S
         => \rptr_s[3]\, Y => OPEN, FCO => \rptr_cry[3]_net_1\);
    
    \memraddr_r[4]\ : SLE
      port map(D => un1_memraddr_r_cry_4_S_0, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[4]\);
    
    \rptr[13]\ : SLE
      port map(D => \rptr_s[13]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rptr[13]_net_1\);
    
    \wptr_cry[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[10]_net_1\, S
         => \wptr_s[11]\, Y => OPEN, FCO => \wptr_cry[11]_net_1\);
    
    \memwaddr_r_2[8]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_8_S_0, D => un4_we_i_9, Y => 
        \memwaddr_r_2[8]_net_1\);
    
    \memwaddr_r[12]\ : SLE
      port map(D => \memwaddr_r_2[12]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[12]\);
    
    \L1.un4_re_i_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => \fifo_MEMRADDR[1]\, B => \fifo_MEMRADDR[2]\, 
        Y => un4_re_i_0);
    
    \rptr_cry[12]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[12]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[11]_net_1\, S
         => \rptr_s[12]\, Y => OPEN, FCO => \rptr_cry[12]_net_1\);
    
    memre_0_a2 : CFG2
      generic map(INIT => x"2")

      port map(A => iRX_FIFO_rd_en_0, B => \iRX_FIFO_Empty_0\, Y
         => \fifo_MEMRE\);
    
    \memraddr_r[11]\ : SLE
      port map(D => \memraddr_r_2[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[11]\);
    
    rdiff_bus_cry_12 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[12]_net_1\, B => 
        \rptr[12]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_11\, S => \rdiff_bus[12]\, Y => OPEN, FCO
         => \rdiff_bus_cry_12\);
    
    \memraddr_r[5]\ : SLE
      port map(D => \memraddr_r_2[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[5]\);
    
    \rptr_gray[6]\ : SLE
      port map(D => \rptr_gray_1[6]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[6]_net_1\);
    
    \memraddr_r[9]\ : SLE
      port map(D => \memraddr_r_2[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[9]\);
    
    \rptr[0]\ : SLE
      port map(D => \rptr_s[0]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[0]_net_1\);
    
    \wptr[10]\ : SLE
      port map(D => \wptr_s[10]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[10]_net_1\);
    
    \L1.un4_we_i_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => \fifo_MEMWADDR[1]\, B => \fifo_MEMWADDR[2]\, 
        Y => un4_we_i_0);
    
    wdiff_bus_cry_1 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[1]_net_1\, B => 
        \rptr_bin_sync2[1]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_0\, S => \wdiff_bus[1]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_1\);
    
    rdiff_bus_cry_2 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[2]_net_1\, B => 
        \rptr[2]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_1\, S => \rdiff_bus[2]\, Y => OPEN, FCO
         => \rdiff_bus_cry_2\);
    
    \wptr_gray[9]\ : SLE
      port map(D => \wptr_gray_1[9]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[9]_net_1\);
    
    \rptr_gray_1[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[4]_net_1\, B => \rptr[5]_net_1\, Y => 
        \rptr_gray_1[4]_net_1\);
    
    \wptr_gray_1[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[8]_net_1\, B => \wptr[9]_net_1\, Y => 
        \wptr_gray_1[8]_net_1\);
    
    Rd_corefifo_grayToBinConv : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_1
      port map(rptr_bin_sync(13) => \rptr_bin_sync[13]\, 
        rptr_bin_sync(12) => \rptr_bin_sync[12]\, 
        rptr_bin_sync(11) => \rptr_bin_sync[11]\, 
        rptr_bin_sync(10) => \rptr_bin_sync[10]\, 
        rptr_bin_sync(9) => \rptr_bin_sync[9]\, rptr_bin_sync(8)
         => \rptr_bin_sync[8]\, rptr_bin_sync(7) => 
        \rptr_bin_sync[7]\, rptr_bin_sync(6) => nc2, 
        rptr_bin_sync(5) => \rptr_bin_sync[5]\, rptr_bin_sync(4)
         => nc1, rptr_bin_sync(3) => \rptr_bin_sync[3]\, 
        rptr_bin_sync(2) => \rptr_bin_sync[2]\, rptr_bin_sync(1)
         => \rptr_bin_sync[1]\, rptr_bin_sync(0) => 
        \rptr_bin_sync[0]\, rptr_gray_sync(12) => 
        \rptr_gray_sync[12]\, rptr_gray_sync(11) => 
        \rptr_gray_sync[11]\, rptr_gray_sync(10) => 
        \rptr_gray_sync[10]\, rptr_gray_sync(9) => 
        \rptr_gray_sync[9]\, rptr_gray_sync(8) => 
        \rptr_gray_sync[8]\, rptr_gray_sync(7) => 
        \rptr_gray_sync[7]\, rptr_gray_sync(6) => 
        \rptr_gray_sync[6]\, rptr_gray_sync(5) => 
        \rptr_gray_sync[5]\, rptr_gray_sync(4) => 
        \rptr_gray_sync[4]\, rptr_gray_sync(3) => 
        \rptr_gray_sync[3]\, rptr_gray_sync(2) => 
        \rptr_gray_sync[2]\, rptr_gray_sync(1) => 
        \rptr_gray_sync[1]\, rptr_gray_sync(0) => 
        \rptr_gray_sync[0]\, bin_N_6_i => bin_N_6_i, bin_N_4_0_i
         => bin_N_4_0_i);
    
    \rptr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => rptr_s_906_FCO, S => 
        \rptr_s[1]\, Y => OPEN, FCO => \rptr_cry[1]_net_1\);
    
    \rptr_cry[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[10]_net_1\, S
         => \rptr_s[11]\, Y => OPEN, FCO => \rptr_cry[11]_net_1\);
    
    rdiff_bus_cry_3 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[3]_net_1\, B => 
        \rptr[3]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_2\, S => \rdiff_bus[3]\, Y => OPEN, FCO
         => \rdiff_bus_cry_3\);
    
    rdiff_bus_cry_10 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[10]_net_1\, B => 
        \rptr[10]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_9\, S => \rdiff_bus[10]\, Y => OPEN, FCO
         => \rdiff_bus_cry_10\);
    
    un1_memwaddr_r_cry_11 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[11]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_10\, 
        S => un1_memwaddr_r_cry_11_S_0, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_11\);
    
    \memraddr_r[6]\ : SLE
      port map(D => un1_memraddr_r_cry_6_S_0, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[6]\);
    
    \rptr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[6]_net_1\, S
         => \rptr_s[7]\, Y => OPEN, FCO => \rptr_cry[7]_net_1\);
    
    rdiff_bus_cry_0 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => rdiff_bus, B => \rptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => rdiff_bus_cry_0_Y_1, FCO => \rdiff_bus_cry_0\);
    
    \memraddr_r[2]\ : SLE
      port map(D => un1_memraddr_r_cry_2_S_0, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[2]\);
    
    \wptr[8]\ : SLE
      port map(D => \wptr_s[8]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[8]_net_1\);
    
    wdiff_bus_cry_3 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[3]_net_1\, B => 
        \rptr_bin_sync2[3]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_2\, S => \wdiff_bus[3]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_3\);
    
    rdiff_bus_s_13 : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \rptr[13]_net_1\, C => 
        \wptr_bin_sync2[13]_net_1\, D => GND_net_1, FCI => 
        \rdiff_bus_cry_12\, S => \rdiff_bus[13]\, Y => OPEN, FCO
         => OPEN);
    
    \memraddr_r[12]\ : SLE
      port map(D => \memraddr_r_2[12]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[12]\);
    
    \wptr_gray_1[11]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[11]_net_1\, B => \wptr[12]_net_1\, Y
         => \wptr_gray_1[11]_net_1\);
    
    \rptr_gray[7]\ : SLE
      port map(D => \rptr_gray_1[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[7]_net_1\);
    
    \wptr_gray[0]\ : SLE
      port map(D => \wptr_gray_1[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[0]_net_1\);
    
    \rptr_gray_1[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[0]_net_1\, B => \rptr[1]_net_1\, Y => 
        \rptr_gray_1[0]_net_1\);
    
    un1_memwaddr_r_cry_10 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_9\, 
        S => un1_memwaddr_r_cry_10_S_0, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_10\);
    
    \rptr_gray_1[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[8]_net_1\, B => \rptr[9]_net_1\, Y => 
        \rptr_gray_1[8]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_0 is

    port( RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          RX_FIFO_DOUT_1            : out   std_logic_vector(8 downto 0);
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_wr_en_0_0        : in    std_logic;
          iRX_FIFO_rd_en_0          : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          RX_FIFO_TxColDetDis_wr_en : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          irx_fifo_rst_i            : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_0;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_0 is 

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_0
    port( fifo_MEMRADDR             : in    std_logic_vector(12 downto 0) := (others => 'U');
          fifo_MEMWADDR             : in    std_logic_vector(12 downto 0) := (others => 'U');
          RDATA_int                 : out   std_logic_vector(8 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          fifo_MEMRE                : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          fifo_MEMWE                : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_0
    port( fifo_MEMRADDR             : out   std_logic_vector(12 downto 0);
          fifo_MEMWADDR             : out   std_logic_vector(12 downto 0);
          iRX_FIFO_wr_en_0_0        : in    std_logic := 'U';
          iRX_FIFO_rd_en_0          : in    std_logic := 'U';
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          RX_FIFO_TxColDetDis_wr_en : in    std_logic := 'U';
          fifo_MEMRE                : out   std_logic;
          fifo_MEMWE                : out   std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          irx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \RDATA_r[0]_net_1\, VCC_net_1, \RDATA_int[0]\, 
        un6_fifo_memre_0, GND_net_1, \RDATA_r[1]_net_1\, 
        \RDATA_int[1]\, \RDATA_r[2]_net_1\, \RDATA_int[2]\, 
        \RDATA_r[3]_net_1\, \RDATA_int[3]\, \RDATA_r[4]_net_1\, 
        \RDATA_int[4]\, \RDATA_r[5]_net_1\, \RDATA_int[5]\, 
        \RDATA_r[6]_net_1\, \RDATA_int[6]\, \RDATA_r[7]_net_1\, 
        \RDATA_int[7]\, \RDATA_r[8]_net_1\, \RDATA_int[8]\, 
        \re_set\, \REN_d1\, un9_fifo_memre_0, fifo_MEMRE, \RE_d1\, 
        \re_pulse_d1\, \re_pulse\, \fifo_MEMRADDR[0]\, 
        \fifo_MEMRADDR[1]\, \fifo_MEMRADDR[2]\, 
        \fifo_MEMRADDR[3]\, \fifo_MEMRADDR[4]\, 
        \fifo_MEMRADDR[5]\, \fifo_MEMRADDR[6]\, 
        \fifo_MEMRADDR[7]\, \fifo_MEMRADDR[8]\, 
        \fifo_MEMRADDR[9]\, \fifo_MEMRADDR[10]\, 
        \fifo_MEMRADDR[11]\, \fifo_MEMRADDR[12]\, 
        \fifo_MEMWADDR[0]\, \fifo_MEMWADDR[1]\, 
        \fifo_MEMWADDR[2]\, \fifo_MEMWADDR[3]\, 
        \fifo_MEMWADDR[4]\, \fifo_MEMWADDR[5]\, 
        \fifo_MEMWADDR[6]\, \fifo_MEMWADDR[7]\, 
        \fifo_MEMWADDR[8]\, \fifo_MEMWADDR[9]\, 
        \fifo_MEMWADDR[10]\, \fifo_MEMWADDR[11]\, 
        \fifo_MEMWADDR[12]\, fifo_MEMWE : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_0
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_0(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_0
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_0(DEF_ARCH);
begin 


    re_pulse : CFG3
      generic map(INIT => x"DC")

      port map(A => fifo_MEMRE, B => \re_set\, C => \REN_d1\, Y
         => \re_pulse\);
    
    \RDATA_r[3]\ : SLE
      port map(D => \RDATA_int[3]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un6_fifo_memre_0, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[3]_net_1\);
    
    \Q[6]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[6]_net_1\, C => 
        \RDATA_int[6]\, D => \RE_d1\, Y => RX_FIFO_DOUT_1(6));
    
    re_pulse_d1 : SLE
      port map(D => \re_pulse\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \re_pulse_d1\);
    
    \RDATA_r[5]\ : SLE
      port map(D => \RDATA_int[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un6_fifo_memre_0, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[5]_net_1\);
    
    un9_fifo_memre : CFG2
      generic map(INIT => x"6")

      port map(A => fifo_MEMRE, B => \REN_d1\, Y => 
        un9_fifo_memre_0);
    
    \RDATA_r[8]\ : SLE
      port map(D => \RDATA_int[8]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un6_fifo_memre_0, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[8]_net_1\);
    
    \Q[2]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[2]_net_1\, C => 
        \RDATA_int[2]\, D => \RE_d1\, Y => RX_FIFO_DOUT_1(2));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \RW1.UI_ram_wrapper_1\ : FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_0
      port map(fifo_MEMRADDR(12) => \fifo_MEMRADDR[12]\, 
        fifo_MEMRADDR(11) => \fifo_MEMRADDR[11]\, 
        fifo_MEMRADDR(10) => \fifo_MEMRADDR[10]\, 
        fifo_MEMRADDR(9) => \fifo_MEMRADDR[9]\, fifo_MEMRADDR(8)
         => \fifo_MEMRADDR[8]\, fifo_MEMRADDR(7) => 
        \fifo_MEMRADDR[7]\, fifo_MEMRADDR(6) => 
        \fifo_MEMRADDR[6]\, fifo_MEMRADDR(5) => 
        \fifo_MEMRADDR[5]\, fifo_MEMRADDR(4) => 
        \fifo_MEMRADDR[4]\, fifo_MEMRADDR(3) => 
        \fifo_MEMRADDR[3]\, fifo_MEMRADDR(2) => 
        \fifo_MEMRADDR[2]\, fifo_MEMRADDR(1) => 
        \fifo_MEMRADDR[1]\, fifo_MEMRADDR(0) => 
        \fifo_MEMRADDR[0]\, fifo_MEMWADDR(12) => 
        \fifo_MEMWADDR[12]\, fifo_MEMWADDR(11) => 
        \fifo_MEMWADDR[11]\, fifo_MEMWADDR(10) => 
        \fifo_MEMWADDR[10]\, fifo_MEMWADDR(9) => 
        \fifo_MEMWADDR[9]\, fifo_MEMWADDR(8) => 
        \fifo_MEMWADDR[8]\, fifo_MEMWADDR(7) => 
        \fifo_MEMWADDR[7]\, fifo_MEMWADDR(6) => 
        \fifo_MEMWADDR[6]\, fifo_MEMWADDR(5) => 
        \fifo_MEMWADDR[5]\, fifo_MEMWADDR(4) => 
        \fifo_MEMWADDR[4]\, fifo_MEMWADDR(3) => 
        \fifo_MEMWADDR[3]\, fifo_MEMWADDR(2) => 
        \fifo_MEMWADDR[2]\, fifo_MEMWADDR(1) => 
        \fifo_MEMWADDR[1]\, fifo_MEMWADDR(0) => 
        \fifo_MEMWADDR[0]\, RDATA_int(8) => \RDATA_int[8]\, 
        RDATA_int(7) => \RDATA_int[7]\, RDATA_int(6) => 
        \RDATA_int[6]\, RDATA_int(5) => \RDATA_int[5]\, 
        RDATA_int(4) => \RDATA_int[4]\, RDATA_int(3) => 
        \RDATA_int[3]\, RDATA_int(2) => \RDATA_int[2]\, 
        RDATA_int(1) => \RDATA_int[1]\, RDATA_int(0) => 
        \RDATA_int[0]\, RX_FIFO_DIN_pipe(8) => 
        RX_FIFO_DIN_pipe(8), RX_FIFO_DIN_pipe(7) => 
        RX_FIFO_DIN_pipe(7), RX_FIFO_DIN_pipe(6) => 
        RX_FIFO_DIN_pipe(6), RX_FIFO_DIN_pipe(5) => 
        RX_FIFO_DIN_pipe(5), RX_FIFO_DIN_pipe(4) => 
        RX_FIFO_DIN_pipe(4), RX_FIFO_DIN_pipe(3) => 
        RX_FIFO_DIN_pipe(3), RX_FIFO_DIN_pipe(2) => 
        RX_FIFO_DIN_pipe(2), RX_FIFO_DIN_pipe(1) => 
        RX_FIFO_DIN_pipe(1), RX_FIFO_DIN_pipe(0) => 
        RX_FIFO_DIN_pipe(0), m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, fifo_MEMRE => fifo_MEMRE, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, fifo_MEMWE
         => fifo_MEMWE);
    
    \RDATA_r[0]\ : SLE
      port map(D => \RDATA_int[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un6_fifo_memre_0, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[0]_net_1\);
    
    \Q[4]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[4]_net_1\, C => 
        \RDATA_int[4]\, D => \RE_d1\, Y => RX_FIFO_DOUT_1(4));
    
    \RDATA_r[2]\ : SLE
      port map(D => \RDATA_int[2]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un6_fifo_memre_0, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[2]_net_1\);
    
    \RDATA_r[6]\ : SLE
      port map(D => \RDATA_int[6]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un6_fifo_memre_0, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[6]_net_1\);
    
    \L31.U_corefifo_async\ : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_0
      port map(fifo_MEMRADDR(12) => \fifo_MEMRADDR[12]\, 
        fifo_MEMRADDR(11) => \fifo_MEMRADDR[11]\, 
        fifo_MEMRADDR(10) => \fifo_MEMRADDR[10]\, 
        fifo_MEMRADDR(9) => \fifo_MEMRADDR[9]\, fifo_MEMRADDR(8)
         => \fifo_MEMRADDR[8]\, fifo_MEMRADDR(7) => 
        \fifo_MEMRADDR[7]\, fifo_MEMRADDR(6) => 
        \fifo_MEMRADDR[6]\, fifo_MEMRADDR(5) => 
        \fifo_MEMRADDR[5]\, fifo_MEMRADDR(4) => 
        \fifo_MEMRADDR[4]\, fifo_MEMRADDR(3) => 
        \fifo_MEMRADDR[3]\, fifo_MEMRADDR(2) => 
        \fifo_MEMRADDR[2]\, fifo_MEMRADDR(1) => 
        \fifo_MEMRADDR[1]\, fifo_MEMRADDR(0) => 
        \fifo_MEMRADDR[0]\, fifo_MEMWADDR(12) => 
        \fifo_MEMWADDR[12]\, fifo_MEMWADDR(11) => 
        \fifo_MEMWADDR[11]\, fifo_MEMWADDR(10) => 
        \fifo_MEMWADDR[10]\, fifo_MEMWADDR(9) => 
        \fifo_MEMWADDR[9]\, fifo_MEMWADDR(8) => 
        \fifo_MEMWADDR[8]\, fifo_MEMWADDR(7) => 
        \fifo_MEMWADDR[7]\, fifo_MEMWADDR(6) => 
        \fifo_MEMWADDR[6]\, fifo_MEMWADDR(5) => 
        \fifo_MEMWADDR[5]\, fifo_MEMWADDR(4) => 
        \fifo_MEMWADDR[4]\, fifo_MEMWADDR(3) => 
        \fifo_MEMWADDR[3]\, fifo_MEMWADDR(2) => 
        \fifo_MEMWADDR[2]\, fifo_MEMWADDR(1) => 
        \fifo_MEMWADDR[1]\, fifo_MEMWADDR(0) => 
        \fifo_MEMWADDR[0]\, iRX_FIFO_wr_en_0_0 => 
        iRX_FIFO_wr_en_0_0, iRX_FIFO_rd_en_0 => iRX_FIFO_rd_en_0, 
        iRX_FIFO_Empty_0 => iRX_FIFO_Empty_0, iRX_FIFO_UNDERRUN_0
         => iRX_FIFO_UNDERRUN_0, iRX_FIFO_OVERFLOW_0 => 
        iRX_FIFO_OVERFLOW_0, iRX_FIFO_Full_0 => iRX_FIFO_Full_0, 
        RX_FIFO_TxColDetDis_wr_en => RX_FIFO_TxColDetDis_wr_en, 
        fifo_MEMRE => fifo_MEMRE, fifo_MEMWE => fifo_MEMWE, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz, 
        irx_fifo_rst_i => irx_fifo_rst_i);
    
    re_set : SLE
      port map(D => \REN_d1\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => un9_fifo_memre_0, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \re_set\);
    
    \Q[3]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[3]_net_1\, C => 
        \RDATA_int[3]\, D => \RE_d1\, Y => RX_FIFO_DOUT_1(3));
    
    \Q[7]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[7]_net_1\, C => 
        \RDATA_int[7]\, D => \RE_d1\, Y => RX_FIFO_DOUT_1(7));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \Q[8]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[8]_net_1\, C => 
        \RDATA_int[8]\, D => \RE_d1\, Y => RX_FIFO_DOUT_1(8));
    
    RE_d1 : SLE
      port map(D => iRX_FIFO_rd_en_0, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RE_d1\);
    
    \RDATA_r[7]\ : SLE
      port map(D => \RDATA_int[7]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un6_fifo_memre_0, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[7]_net_1\);
    
    \RDATA_r[4]\ : SLE
      port map(D => \RDATA_int[4]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un6_fifo_memre_0, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[4]_net_1\);
    
    \Q[1]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[1]_net_1\, C => 
        \RDATA_int[1]\, D => \RE_d1\, Y => RX_FIFO_DOUT_1(1));
    
    \Q[0]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[0]_net_1\, C => 
        \RDATA_int[0]\, D => \RE_d1\, Y => RX_FIFO_DOUT_1(0));
    
    REN_d1 : SLE
      port map(D => fifo_MEMRE, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \REN_d1\);
    
    \Q[5]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[5]_net_1\, C => 
        \RDATA_int[5]\, D => \RE_d1\, Y => RX_FIFO_DOUT_1(5));
    
    un6_fifo_memre : CFG2
      generic map(INIT => x"4")

      port map(A => fifo_MEMRE, B => \REN_d1\, Y => 
        un6_fifo_memre_0);
    
    \RDATA_r[1]\ : SLE
      port map(D => \RDATA_int[1]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un6_fifo_memre_0, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[1]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_0 is

    port( RX_FIFO_DOUT_1            : out   std_logic_vector(8 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          iRX_FIFO_rd_en_0          : in    std_logic;
          iRX_FIFO_wr_en_0_0        : in    std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          irx_fifo_rst_i            : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          RX_FIFO_TxColDetDis_wr_en : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic
        );

end FIFO_8Kx9_0;

architecture DEF_ARCH of FIFO_8Kx9_0 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_0
    port( RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          RX_FIFO_DOUT_1            : out   std_logic_vector(8 downto 0);
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_wr_en_0_0        : in    std_logic := 'U';
          iRX_FIFO_rd_en_0          : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          RX_FIFO_TxColDetDis_wr_en : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          irx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_0
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_0(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    FIFO_8Kx9_0 : FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_0
      port map(RX_FIFO_DIN_pipe(8) => RX_FIFO_DIN_pipe(8), 
        RX_FIFO_DIN_pipe(7) => RX_FIFO_DIN_pipe(7), 
        RX_FIFO_DIN_pipe(6) => RX_FIFO_DIN_pipe(6), 
        RX_FIFO_DIN_pipe(5) => RX_FIFO_DIN_pipe(5), 
        RX_FIFO_DIN_pipe(4) => RX_FIFO_DIN_pipe(4), 
        RX_FIFO_DIN_pipe(3) => RX_FIFO_DIN_pipe(3), 
        RX_FIFO_DIN_pipe(2) => RX_FIFO_DIN_pipe(2), 
        RX_FIFO_DIN_pipe(1) => RX_FIFO_DIN_pipe(1), 
        RX_FIFO_DIN_pipe(0) => RX_FIFO_DIN_pipe(0), 
        RX_FIFO_DOUT_1(8) => RX_FIFO_DOUT_1(8), RX_FIFO_DOUT_1(7)
         => RX_FIFO_DOUT_1(7), RX_FIFO_DOUT_1(6) => 
        RX_FIFO_DOUT_1(6), RX_FIFO_DOUT_1(5) => RX_FIFO_DOUT_1(5), 
        RX_FIFO_DOUT_1(4) => RX_FIFO_DOUT_1(4), RX_FIFO_DOUT_1(3)
         => RX_FIFO_DOUT_1(3), RX_FIFO_DOUT_1(2) => 
        RX_FIFO_DOUT_1(2), RX_FIFO_DOUT_1(1) => RX_FIFO_DOUT_1(1), 
        RX_FIFO_DOUT_1(0) => RX_FIFO_DOUT_1(0), iRX_FIFO_Full_0
         => iRX_FIFO_Full_0, iRX_FIFO_OVERFLOW_0 => 
        iRX_FIFO_OVERFLOW_0, iRX_FIFO_UNDERRUN_0 => 
        iRX_FIFO_UNDERRUN_0, iRX_FIFO_Empty_0 => iRX_FIFO_Empty_0, 
        iRX_FIFO_wr_en_0_0 => iRX_FIFO_wr_en_0_0, 
        iRX_FIFO_rd_en_0 => iRX_FIFO_rd_en_0, CommsFPGA_CCC_0_GL0
         => CommsFPGA_CCC_0_GL0, RX_FIFO_TxColDetDis_wr_en => 
        RX_FIFO_TxColDetDis_wr_en, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, irx_fifo_rst_i => 
        irx_fifo_rst_i);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_1 is

    port( RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          RDATA_int                 : out   std_logic_vector(8 downto 0);
          fifo_MEMWADDR             : in    std_logic_vector(12 downto 0);
          fifo_MEMRADDR             : in    std_logic_vector(12 downto 0);
          fifo_MEMWE                : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          fifo_MEMRE                : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_1;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_1 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component RAM1K18
    generic (MEMORYFILE:string := "");

    port( A_DOUT        : out   std_logic_vector(17 downto 0);
          B_DOUT        : out   std_logic_vector(17 downto 0);
          BUSY          : out   std_logic;
          A_CLK         : in    std_logic := 'U';
          A_DOUT_CLK    : in    std_logic := 'U';
          A_ARST_N      : in    std_logic := 'U';
          A_DOUT_EN     : in    std_logic := 'U';
          A_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_DOUT_ARST_N : in    std_logic := 'U';
          A_DOUT_SRST_N : in    std_logic := 'U';
          A_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          A_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          A_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          B_CLK         : in    std_logic := 'U';
          B_DOUT_CLK    : in    std_logic := 'U';
          B_ARST_N      : in    std_logic := 'U';
          B_DOUT_EN     : in    std_logic := 'U';
          B_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_DOUT_ARST_N : in    std_logic := 'U';
          B_DOUT_SRST_N : in    std_logic := 'U';
          B_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          B_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          B_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          A_EN          : in    std_logic := 'U';
          A_DOUT_LAT    : in    std_logic := 'U';
          A_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_WMODE       : in    std_logic := 'U';
          B_EN          : in    std_logic := 'U';
          B_DOUT_LAT    : in    std_logic := 'U';
          B_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_WMODE       : in    std_logic := 'U';
          SII_LOCK      : in    std_logic := 'U'
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;
    signal nc151, nc23, nc58, nc116, nc74, nc133, nc167, nc84, 
        nc39, nc72, nc82, nc145, nc160, nc57, nc156, nc125, nc73, 
        nc107, nc66, nc83, nc9, nc171, nc54, nc135, nc41, nc100, 
        nc52, nc29, nc118, nc60, nc141, nc45, nc53, nc121, nc158, 
        nc162, nc11, nc131, nc96, nc79, nc146, nc89, nc119, nc48, 
        nc126, nc15, nc102, nc3, nc47, nc90, nc159, nc136, nc59, 
        nc18, nc44, nc117, nc164, nc148, nc42, nc17, nc2, nc110, 
        nc128, nc43, nc157, nc36, nc61, nc104, nc138, nc14, nc150, 
        nc149, nc12, nc30, nc65, nc7, nc129, nc8, nc13, nc26, 
        nc139, nc163, nc112, nc68, nc49, nc170, nc91, nc5, nc20, 
        nc147, nc67, nc152, nc127, nc103, nc76, nc140, nc86, nc95, 
        nc120, nc165, nc137, nc64, nc19, nc70, nc62, nc80, nc130, 
        nc98, nc114, nc56, nc105, nc63, nc97, nc161, nc31, nc154, 
        nc50, nc142, nc94, nc122, nc35, nc4, nc92, nc101, nc166, 
        nc132, nc21, nc93, nc69, nc38, nc113, nc106, nc25, nc1, 
        nc37, nc144, nc153, nc46, nc71, nc124, nc81, nc168, nc34, 
        nc28, nc115, nc134, nc32, nc40, nc99, nc75, nc85, nc27, 
        nc108, nc16, nc155, nc51, nc33, nc169, nc78, nc24, nc88, 
        nc111, nc55, nc10, nc22, nc143, nc77, nc6, nc109, nc87, 
        nc123 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C2 : RAM1K18
      port map(A_DOUT(17) => nc151, A_DOUT(16) => nc23, 
        A_DOUT(15) => nc58, A_DOUT(14) => nc116, A_DOUT(13) => 
        nc74, A_DOUT(12) => nc133, A_DOUT(11) => nc167, 
        A_DOUT(10) => nc84, A_DOUT(9) => nc39, A_DOUT(8) => nc72, 
        A_DOUT(7) => nc82, A_DOUT(6) => nc145, A_DOUT(5) => nc160, 
        A_DOUT(4) => nc57, A_DOUT(3) => nc156, A_DOUT(2) => nc125, 
        A_DOUT(1) => RDATA_int(5), A_DOUT(0) => RDATA_int(4), 
        B_DOUT(17) => nc73, B_DOUT(16) => nc107, B_DOUT(15) => 
        nc66, B_DOUT(14) => nc83, B_DOUT(13) => nc9, B_DOUT(12)
         => nc171, B_DOUT(11) => nc54, B_DOUT(10) => nc135, 
        B_DOUT(9) => nc41, B_DOUT(8) => nc100, B_DOUT(7) => nc52, 
        B_DOUT(6) => nc29, B_DOUT(5) => nc118, B_DOUT(4) => nc60, 
        B_DOUT(3) => nc141, B_DOUT(2) => nc45, B_DOUT(1) => nc53, 
        B_DOUT(0) => nc121, BUSY => OPEN, A_CLK => 
        m2s010_som_sb_0_CCC_71MHz, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => fifo_MEMRE, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => fifo_MEMRADDR(12), A_ADDR(12) => fifo_MEMRADDR(11), 
        A_ADDR(11) => fifo_MEMRADDR(10), A_ADDR(10) => 
        fifo_MEMRADDR(9), A_ADDR(9) => fifo_MEMRADDR(8), 
        A_ADDR(8) => fifo_MEMRADDR(7), A_ADDR(7) => 
        fifo_MEMRADDR(6), A_ADDR(6) => fifo_MEMRADDR(5), 
        A_ADDR(5) => fifo_MEMRADDR(4), A_ADDR(4) => 
        fifo_MEMRADDR(3), A_ADDR(3) => fifo_MEMRADDR(2), 
        A_ADDR(2) => fifo_MEMRADDR(1), A_ADDR(1) => 
        fifo_MEMRADDR(0), A_ADDR(0) => GND_net_1, A_WEN(1) => 
        GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => GND_net_1, B_DIN(2) => GND_net_1, B_DIN(1)
         => RX_FIFO_DIN_pipe(5), B_DIN(0) => RX_FIFO_DIN_pipe(4), 
        B_ADDR(13) => fifo_MEMWADDR(12), B_ADDR(12) => 
        fifo_MEMWADDR(11), B_ADDR(11) => fifo_MEMWADDR(10), 
        B_ADDR(10) => fifo_MEMWADDR(9), B_ADDR(9) => 
        fifo_MEMWADDR(8), B_ADDR(8) => fifo_MEMWADDR(7), 
        B_ADDR(7) => fifo_MEMWADDR(6), B_ADDR(6) => 
        fifo_MEMWADDR(5), B_ADDR(5) => fifo_MEMWADDR(4), 
        B_ADDR(4) => fifo_MEMWADDR(3), B_ADDR(3) => 
        fifo_MEMWADDR(2), B_ADDR(2) => fifo_MEMWADDR(1), 
        B_ADDR(1) => fifo_MEMWADDR(0), B_ADDR(0) => GND_net_1, 
        B_WEN(1) => GND_net_1, B_WEN(0) => VCC_net_1, A_EN => 
        VCC_net_1, A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => 
        GND_net_1, A_WIDTH(1) => GND_net_1, A_WIDTH(0) => 
        VCC_net_1, A_WMODE => GND_net_1, B_EN => VCC_net_1, 
        B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => GND_net_1, 
        B_WIDTH(1) => GND_net_1, B_WIDTH(0) => VCC_net_1, B_WMODE
         => GND_net_1, SII_LOCK => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C1 : RAM1K18
      port map(A_DOUT(17) => nc158, A_DOUT(16) => nc162, 
        A_DOUT(15) => nc11, A_DOUT(14) => nc131, A_DOUT(13) => 
        nc96, A_DOUT(12) => nc79, A_DOUT(11) => nc146, A_DOUT(10)
         => nc89, A_DOUT(9) => nc119, A_DOUT(8) => nc48, 
        A_DOUT(7) => nc126, A_DOUT(6) => nc15, A_DOUT(5) => nc102, 
        A_DOUT(4) => nc3, A_DOUT(3) => nc47, A_DOUT(2) => nc90, 
        A_DOUT(1) => RDATA_int(3), A_DOUT(0) => RDATA_int(2), 
        B_DOUT(17) => nc159, B_DOUT(16) => nc136, B_DOUT(15) => 
        nc59, B_DOUT(14) => nc18, B_DOUT(13) => nc44, B_DOUT(12)
         => nc117, B_DOUT(11) => nc164, B_DOUT(10) => nc148, 
        B_DOUT(9) => nc42, B_DOUT(8) => nc17, B_DOUT(7) => nc2, 
        B_DOUT(6) => nc110, B_DOUT(5) => nc128, B_DOUT(4) => nc43, 
        B_DOUT(3) => nc157, B_DOUT(2) => nc36, B_DOUT(1) => nc61, 
        B_DOUT(0) => nc104, BUSY => OPEN, A_CLK => 
        m2s010_som_sb_0_CCC_71MHz, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => fifo_MEMRE, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => fifo_MEMRADDR(12), A_ADDR(12) => fifo_MEMRADDR(11), 
        A_ADDR(11) => fifo_MEMRADDR(10), A_ADDR(10) => 
        fifo_MEMRADDR(9), A_ADDR(9) => fifo_MEMRADDR(8), 
        A_ADDR(8) => fifo_MEMRADDR(7), A_ADDR(7) => 
        fifo_MEMRADDR(6), A_ADDR(6) => fifo_MEMRADDR(5), 
        A_ADDR(5) => fifo_MEMRADDR(4), A_ADDR(4) => 
        fifo_MEMRADDR(3), A_ADDR(3) => fifo_MEMRADDR(2), 
        A_ADDR(2) => fifo_MEMRADDR(1), A_ADDR(1) => 
        fifo_MEMRADDR(0), A_ADDR(0) => GND_net_1, A_WEN(1) => 
        GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => GND_net_1, B_DIN(2) => GND_net_1, B_DIN(1)
         => RX_FIFO_DIN_pipe(3), B_DIN(0) => RX_FIFO_DIN_pipe(2), 
        B_ADDR(13) => fifo_MEMWADDR(12), B_ADDR(12) => 
        fifo_MEMWADDR(11), B_ADDR(11) => fifo_MEMWADDR(10), 
        B_ADDR(10) => fifo_MEMWADDR(9), B_ADDR(9) => 
        fifo_MEMWADDR(8), B_ADDR(8) => fifo_MEMWADDR(7), 
        B_ADDR(7) => fifo_MEMWADDR(6), B_ADDR(6) => 
        fifo_MEMWADDR(5), B_ADDR(5) => fifo_MEMWADDR(4), 
        B_ADDR(4) => fifo_MEMWADDR(3), B_ADDR(3) => 
        fifo_MEMWADDR(2), B_ADDR(2) => fifo_MEMWADDR(1), 
        B_ADDR(1) => fifo_MEMWADDR(0), B_ADDR(0) => GND_net_1, 
        B_WEN(1) => GND_net_1, B_WEN(0) => VCC_net_1, A_EN => 
        VCC_net_1, A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => 
        GND_net_1, A_WIDTH(1) => GND_net_1, A_WIDTH(0) => 
        VCC_net_1, A_WMODE => GND_net_1, B_EN => VCC_net_1, 
        B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => GND_net_1, 
        B_WIDTH(1) => GND_net_1, B_WIDTH(0) => VCC_net_1, B_WMODE
         => GND_net_1, SII_LOCK => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C4 : RAM1K18
      port map(A_DOUT(17) => nc138, A_DOUT(16) => nc14, 
        A_DOUT(15) => nc150, A_DOUT(14) => nc149, A_DOUT(13) => 
        nc12, A_DOUT(12) => nc30, A_DOUT(11) => nc65, A_DOUT(10)
         => nc7, A_DOUT(9) => nc129, A_DOUT(8) => nc8, A_DOUT(7)
         => nc13, A_DOUT(6) => nc26, A_DOUT(5) => nc139, 
        A_DOUT(4) => nc163, A_DOUT(3) => nc112, A_DOUT(2) => nc68, 
        A_DOUT(1) => nc49, A_DOUT(0) => RDATA_int(8), B_DOUT(17)
         => nc170, B_DOUT(16) => nc91, B_DOUT(15) => nc5, 
        B_DOUT(14) => nc20, B_DOUT(13) => nc147, B_DOUT(12) => 
        nc67, B_DOUT(11) => nc152, B_DOUT(10) => nc127, B_DOUT(9)
         => nc103, B_DOUT(8) => nc76, B_DOUT(7) => nc140, 
        B_DOUT(6) => nc86, B_DOUT(5) => nc95, B_DOUT(4) => nc120, 
        B_DOUT(3) => nc165, B_DOUT(2) => nc137, B_DOUT(1) => nc64, 
        B_DOUT(0) => nc19, BUSY => OPEN, A_CLK => 
        m2s010_som_sb_0_CCC_71MHz, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => fifo_MEMRE, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => fifo_MEMRADDR(12), A_ADDR(12) => fifo_MEMRADDR(11), 
        A_ADDR(11) => fifo_MEMRADDR(10), A_ADDR(10) => 
        fifo_MEMRADDR(9), A_ADDR(9) => fifo_MEMRADDR(8), 
        A_ADDR(8) => fifo_MEMRADDR(7), A_ADDR(7) => 
        fifo_MEMRADDR(6), A_ADDR(6) => fifo_MEMRADDR(5), 
        A_ADDR(5) => fifo_MEMRADDR(4), A_ADDR(4) => 
        fifo_MEMRADDR(3), A_ADDR(3) => fifo_MEMRADDR(2), 
        A_ADDR(2) => fifo_MEMRADDR(1), A_ADDR(1) => 
        fifo_MEMRADDR(0), A_ADDR(0) => GND_net_1, A_WEN(1) => 
        GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => GND_net_1, B_DIN(2) => GND_net_1, B_DIN(1)
         => GND_net_1, B_DIN(0) => RX_FIFO_DIN_pipe(8), 
        B_ADDR(13) => fifo_MEMWADDR(12), B_ADDR(12) => 
        fifo_MEMWADDR(11), B_ADDR(11) => fifo_MEMWADDR(10), 
        B_ADDR(10) => fifo_MEMWADDR(9), B_ADDR(9) => 
        fifo_MEMWADDR(8), B_ADDR(8) => fifo_MEMWADDR(7), 
        B_ADDR(7) => fifo_MEMWADDR(6), B_ADDR(6) => 
        fifo_MEMWADDR(5), B_ADDR(5) => fifo_MEMWADDR(4), 
        B_ADDR(4) => fifo_MEMWADDR(3), B_ADDR(3) => 
        fifo_MEMWADDR(2), B_ADDR(2) => fifo_MEMWADDR(1), 
        B_ADDR(1) => fifo_MEMWADDR(0), B_ADDR(0) => GND_net_1, 
        B_WEN(1) => GND_net_1, B_WEN(0) => VCC_net_1, A_EN => 
        VCC_net_1, A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => 
        GND_net_1, A_WIDTH(1) => GND_net_1, A_WIDTH(0) => 
        VCC_net_1, A_WMODE => GND_net_1, B_EN => VCC_net_1, 
        B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => GND_net_1, 
        B_WIDTH(1) => GND_net_1, B_WIDTH(0) => VCC_net_1, B_WMODE
         => GND_net_1, SII_LOCK => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C3 : RAM1K18
      port map(A_DOUT(17) => nc70, A_DOUT(16) => nc62, A_DOUT(15)
         => nc80, A_DOUT(14) => nc130, A_DOUT(13) => nc98, 
        A_DOUT(12) => nc114, A_DOUT(11) => nc56, A_DOUT(10) => 
        nc105, A_DOUT(9) => nc63, A_DOUT(8) => nc97, A_DOUT(7)
         => nc161, A_DOUT(6) => nc31, A_DOUT(5) => nc154, 
        A_DOUT(4) => nc50, A_DOUT(3) => nc142, A_DOUT(2) => nc94, 
        A_DOUT(1) => RDATA_int(7), A_DOUT(0) => RDATA_int(6), 
        B_DOUT(17) => nc122, B_DOUT(16) => nc35, B_DOUT(15) => 
        nc4, B_DOUT(14) => nc92, B_DOUT(13) => nc101, B_DOUT(12)
         => nc166, B_DOUT(11) => nc132, B_DOUT(10) => nc21, 
        B_DOUT(9) => nc93, B_DOUT(8) => nc69, B_DOUT(7) => nc38, 
        B_DOUT(6) => nc113, B_DOUT(5) => nc106, B_DOUT(4) => nc25, 
        B_DOUT(3) => nc1, B_DOUT(2) => nc37, B_DOUT(1) => nc144, 
        B_DOUT(0) => nc153, BUSY => OPEN, A_CLK => 
        m2s010_som_sb_0_CCC_71MHz, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => fifo_MEMRE, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => fifo_MEMRADDR(12), A_ADDR(12) => fifo_MEMRADDR(11), 
        A_ADDR(11) => fifo_MEMRADDR(10), A_ADDR(10) => 
        fifo_MEMRADDR(9), A_ADDR(9) => fifo_MEMRADDR(8), 
        A_ADDR(8) => fifo_MEMRADDR(7), A_ADDR(7) => 
        fifo_MEMRADDR(6), A_ADDR(6) => fifo_MEMRADDR(5), 
        A_ADDR(5) => fifo_MEMRADDR(4), A_ADDR(4) => 
        fifo_MEMRADDR(3), A_ADDR(3) => fifo_MEMRADDR(2), 
        A_ADDR(2) => fifo_MEMRADDR(1), A_ADDR(1) => 
        fifo_MEMRADDR(0), A_ADDR(0) => GND_net_1, A_WEN(1) => 
        GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => GND_net_1, B_DIN(2) => GND_net_1, B_DIN(1)
         => RX_FIFO_DIN_pipe(7), B_DIN(0) => RX_FIFO_DIN_pipe(6), 
        B_ADDR(13) => fifo_MEMWADDR(12), B_ADDR(12) => 
        fifo_MEMWADDR(11), B_ADDR(11) => fifo_MEMWADDR(10), 
        B_ADDR(10) => fifo_MEMWADDR(9), B_ADDR(9) => 
        fifo_MEMWADDR(8), B_ADDR(8) => fifo_MEMWADDR(7), 
        B_ADDR(7) => fifo_MEMWADDR(6), B_ADDR(6) => 
        fifo_MEMWADDR(5), B_ADDR(5) => fifo_MEMWADDR(4), 
        B_ADDR(4) => fifo_MEMWADDR(3), B_ADDR(3) => 
        fifo_MEMWADDR(2), B_ADDR(2) => fifo_MEMWADDR(1), 
        B_ADDR(1) => fifo_MEMWADDR(0), B_ADDR(0) => GND_net_1, 
        B_WEN(1) => GND_net_1, B_WEN(0) => VCC_net_1, A_EN => 
        VCC_net_1, A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => 
        GND_net_1, A_WIDTH(1) => GND_net_1, A_WIDTH(0) => 
        VCC_net_1, A_WMODE => GND_net_1, B_EN => VCC_net_1, 
        B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => GND_net_1, 
        B_WIDTH(1) => GND_net_1, B_WIDTH(0) => VCC_net_1, B_WMODE
         => GND_net_1, SII_LOCK => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C0 : RAM1K18
      port map(A_DOUT(17) => nc46, A_DOUT(16) => nc71, A_DOUT(15)
         => nc124, A_DOUT(14) => nc81, A_DOUT(13) => nc168, 
        A_DOUT(12) => nc34, A_DOUT(11) => nc28, A_DOUT(10) => 
        nc115, A_DOUT(9) => nc134, A_DOUT(8) => nc32, A_DOUT(7)
         => nc40, A_DOUT(6) => nc99, A_DOUT(5) => nc75, A_DOUT(4)
         => nc85, A_DOUT(3) => nc27, A_DOUT(2) => nc108, 
        A_DOUT(1) => RDATA_int(1), A_DOUT(0) => RDATA_int(0), 
        B_DOUT(17) => nc16, B_DOUT(16) => nc155, B_DOUT(15) => 
        nc51, B_DOUT(14) => nc33, B_DOUT(13) => nc169, B_DOUT(12)
         => nc78, B_DOUT(11) => nc24, B_DOUT(10) => nc88, 
        B_DOUT(9) => nc111, B_DOUT(8) => nc55, B_DOUT(7) => nc10, 
        B_DOUT(6) => nc22, B_DOUT(5) => nc143, B_DOUT(4) => nc77, 
        B_DOUT(3) => nc6, B_DOUT(2) => nc109, B_DOUT(1) => nc87, 
        B_DOUT(0) => nc123, BUSY => OPEN, A_CLK => 
        m2s010_som_sb_0_CCC_71MHz, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => fifo_MEMRE, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => fifo_MEMRADDR(12), A_ADDR(12) => fifo_MEMRADDR(11), 
        A_ADDR(11) => fifo_MEMRADDR(10), A_ADDR(10) => 
        fifo_MEMRADDR(9), A_ADDR(9) => fifo_MEMRADDR(8), 
        A_ADDR(8) => fifo_MEMRADDR(7), A_ADDR(7) => 
        fifo_MEMRADDR(6), A_ADDR(6) => fifo_MEMRADDR(5), 
        A_ADDR(5) => fifo_MEMRADDR(4), A_ADDR(4) => 
        fifo_MEMRADDR(3), A_ADDR(3) => fifo_MEMRADDR(2), 
        A_ADDR(2) => fifo_MEMRADDR(1), A_ADDR(1) => 
        fifo_MEMRADDR(0), A_ADDR(0) => GND_net_1, A_WEN(1) => 
        GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => GND_net_1, B_DIN(2) => GND_net_1, B_DIN(1)
         => RX_FIFO_DIN_pipe(1), B_DIN(0) => RX_FIFO_DIN_pipe(0), 
        B_ADDR(13) => fifo_MEMWADDR(12), B_ADDR(12) => 
        fifo_MEMWADDR(11), B_ADDR(11) => fifo_MEMWADDR(10), 
        B_ADDR(10) => fifo_MEMWADDR(9), B_ADDR(9) => 
        fifo_MEMWADDR(8), B_ADDR(8) => fifo_MEMWADDR(7), 
        B_ADDR(7) => fifo_MEMWADDR(6), B_ADDR(6) => 
        fifo_MEMWADDR(5), B_ADDR(5) => fifo_MEMWADDR(4), 
        B_ADDR(4) => fifo_MEMWADDR(3), B_ADDR(3) => 
        fifo_MEMWADDR(2), B_ADDR(2) => fifo_MEMWADDR(1), 
        B_ADDR(1) => fifo_MEMWADDR(0), B_ADDR(0) => GND_net_1, 
        B_WEN(1) => GND_net_1, B_WEN(0) => VCC_net_1, A_EN => 
        VCC_net_1, A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => 
        GND_net_1, A_WIDTH(1) => GND_net_1, A_WIDTH(0) => 
        VCC_net_1, A_WMODE => GND_net_1, B_EN => VCC_net_1, 
        B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => GND_net_1, 
        B_WIDTH(1) => GND_net_1, B_WIDTH(0) => VCC_net_1, B_WMODE
         => GND_net_1, SII_LOCK => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_1 is

    port( fifo_MEMRADDR             : in    std_logic_vector(12 downto 0);
          fifo_MEMWADDR             : in    std_logic_vector(12 downto 0);
          RDATA_int                 : out   std_logic_vector(8 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          fifo_MEMRE                : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          fifo_MEMWE                : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_1;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_1 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_1
    port( RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          RDATA_int                 : out   std_logic_vector(8 downto 0);
          fifo_MEMWADDR             : in    std_logic_vector(12 downto 0) := (others => 'U');
          fifo_MEMRADDR             : in    std_logic_vector(12 downto 0) := (others => 'U');
          fifo_MEMWE                : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          fifo_MEMRE                : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_1
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_1(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    L1_asyncnonpipe : FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_1
      port map(RX_FIFO_DIN_pipe(8) => RX_FIFO_DIN_pipe(8), 
        RX_FIFO_DIN_pipe(7) => RX_FIFO_DIN_pipe(7), 
        RX_FIFO_DIN_pipe(6) => RX_FIFO_DIN_pipe(6), 
        RX_FIFO_DIN_pipe(5) => RX_FIFO_DIN_pipe(5), 
        RX_FIFO_DIN_pipe(4) => RX_FIFO_DIN_pipe(4), 
        RX_FIFO_DIN_pipe(3) => RX_FIFO_DIN_pipe(3), 
        RX_FIFO_DIN_pipe(2) => RX_FIFO_DIN_pipe(2), 
        RX_FIFO_DIN_pipe(1) => RX_FIFO_DIN_pipe(1), 
        RX_FIFO_DIN_pipe(0) => RX_FIFO_DIN_pipe(0), RDATA_int(8)
         => RDATA_int(8), RDATA_int(7) => RDATA_int(7), 
        RDATA_int(6) => RDATA_int(6), RDATA_int(5) => 
        RDATA_int(5), RDATA_int(4) => RDATA_int(4), RDATA_int(3)
         => RDATA_int(3), RDATA_int(2) => RDATA_int(2), 
        RDATA_int(1) => RDATA_int(1), RDATA_int(0) => 
        RDATA_int(0), fifo_MEMWADDR(12) => fifo_MEMWADDR(12), 
        fifo_MEMWADDR(11) => fifo_MEMWADDR(11), fifo_MEMWADDR(10)
         => fifo_MEMWADDR(10), fifo_MEMWADDR(9) => 
        fifo_MEMWADDR(9), fifo_MEMWADDR(8) => fifo_MEMWADDR(8), 
        fifo_MEMWADDR(7) => fifo_MEMWADDR(7), fifo_MEMWADDR(6)
         => fifo_MEMWADDR(6), fifo_MEMWADDR(5) => 
        fifo_MEMWADDR(5), fifo_MEMWADDR(4) => fifo_MEMWADDR(4), 
        fifo_MEMWADDR(3) => fifo_MEMWADDR(3), fifo_MEMWADDR(2)
         => fifo_MEMWADDR(2), fifo_MEMWADDR(1) => 
        fifo_MEMWADDR(1), fifo_MEMWADDR(0) => fifo_MEMWADDR(0), 
        fifo_MEMRADDR(12) => fifo_MEMRADDR(12), fifo_MEMRADDR(11)
         => fifo_MEMRADDR(11), fifo_MEMRADDR(10) => 
        fifo_MEMRADDR(10), fifo_MEMRADDR(9) => fifo_MEMRADDR(9), 
        fifo_MEMRADDR(8) => fifo_MEMRADDR(8), fifo_MEMRADDR(7)
         => fifo_MEMRADDR(7), fifo_MEMRADDR(6) => 
        fifo_MEMRADDR(6), fifo_MEMRADDR(5) => fifo_MEMRADDR(5), 
        fifo_MEMRADDR(4) => fifo_MEMRADDR(4), fifo_MEMRADDR(3)
         => fifo_MEMRADDR(3), fifo_MEMRADDR(2) => 
        fifo_MEMRADDR(2), fifo_MEMRADDR(1) => fifo_MEMRADDR(1), 
        fifo_MEMRADDR(0) => fifo_MEMRADDR(0), fifo_MEMWE => 
        fifo_MEMWE, CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, 
        fifo_MEMRE => fifo_MEMRE, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_4 is

    port( wptr_bin_sync  : inout std_logic_vector(13 downto 0) := (others => 'Z');
          wptr_gray_sync : in    std_logic_vector(12 downto 0)
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_4;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_4 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    \bin_out_xhdl1_0_a2[1]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(3), B => wptr_gray_sync(1), C
         => wptr_bin_sync(4), D => wptr_gray_sync(2), Y => 
        wptr_bin_sync(1));
    
    \bin_out_xhdl1_0_a2[10]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(12), B => wptr_gray_sync(11), 
        C => wptr_gray_sync(10), D => wptr_bin_sync(13), Y => 
        wptr_bin_sync(10));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \bin_out_xhdl1_0_a2[5]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(7), B => wptr_gray_sync(6), C
         => wptr_gray_sync(5), D => wptr_bin_sync(8), Y => 
        wptr_bin_sync(5));
    
    \bin_out_xhdl1_0_a2[2]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(4), B => wptr_gray_sync(3), C
         => wptr_gray_sync(2), D => wptr_bin_sync(5), Y => 
        wptr_bin_sync(2));
    
    \bin_out_xhdl1_0_a2[0]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(2), B => wptr_bin_sync(3), C
         => wptr_gray_sync(0), D => wptr_gray_sync(1), Y => 
        wptr_bin_sync(0));
    
    \bin_out_xhdl1_0_a2[9]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(11), B => wptr_gray_sync(10), 
        C => wptr_gray_sync(9), D => wptr_bin_sync(12), Y => 
        wptr_bin_sync(9));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \bin_out_xhdl1_i_o2[12]\ : CFG2
      generic map(INIT => x"6")

      port map(A => wptr_bin_sync(13), B => wptr_gray_sync(12), Y
         => wptr_bin_sync(12));
    
    \bin_out_xhdl1_0_a2[6]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(8), B => wptr_gray_sync(7), C
         => wptr_gray_sync(6), D => wptr_bin_sync(9), Y => 
        wptr_bin_sync(6));
    
    \bin_out_xhdl1_0_a2[4]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(6), B => wptr_gray_sync(5), C
         => wptr_gray_sync(4), D => wptr_bin_sync(7), Y => 
        wptr_bin_sync(4));
    
    \bin_out_xhdl1_i_o2[11]\ : CFG3
      generic map(INIT => x"96")

      port map(A => wptr_gray_sync(12), B => wptr_gray_sync(11), 
        C => wptr_bin_sync(13), Y => wptr_bin_sync(11));
    
    \bin_out_xhdl1_0_a2[8]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(10), B => wptr_gray_sync(9), C
         => wptr_gray_sync(8), D => wptr_bin_sync(11), Y => 
        wptr_bin_sync(8));
    
    \bin_out_xhdl1_0_a2[7]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(9), B => wptr_gray_sync(8), C
         => wptr_gray_sync(7), D => wptr_bin_sync(10), Y => 
        wptr_bin_sync(7));
    
    \bin_out_xhdl1_0_a2[3]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(5), B => wptr_gray_sync(4), C
         => wptr_gray_sync(3), D => wptr_bin_sync(6), Y => 
        wptr_bin_sync(3));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_2 is

    port( wptr_gray                 : in    std_logic_vector(13 downto 0);
          wptr_gray_sync            : out   std_logic_vector(12 downto 0);
          wptr_bin_sync_0           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          irx_fifo_rst_i            : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_2;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_2 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \sync_int[11]_net_1\, GND_net_1, 
        \sync_int[12]_net_1\, \sync_int[13]_net_1\, 
        \sync_int[10]_net_1\, \sync_int[0]_net_1\, 
        \sync_int[1]_net_1\, \sync_int[2]_net_1\, 
        \sync_int[3]_net_1\, \sync_int[4]_net_1\, 
        \sync_int[5]_net_1\, \sync_int[6]_net_1\, 
        \sync_int[7]_net_1\, \sync_int[8]_net_1\, 
        \sync_int[9]_net_1\ : std_logic;

begin 


    \sync_int[9]\ : SLE
      port map(D => wptr_gray(9), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[9]_net_1\);
    
    \sync_int[4]\ : SLE
      port map(D => wptr_gray(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[4]_net_1\);
    
    \sync_out_xhdl1[10]\ : SLE
      port map(D => \sync_int[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(10));
    
    \sync_int[1]\ : SLE
      port map(D => wptr_gray(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[1]_net_1\);
    
    \sync_int[11]\ : SLE
      port map(D => wptr_gray(11), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[11]_net_1\);
    
    \sync_out_xhdl1[6]\ : SLE
      port map(D => \sync_int[6]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(6));
    
    \sync_out_xhdl1[3]\ : SLE
      port map(D => \sync_int[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(3));
    
    \sync_int[6]\ : SLE
      port map(D => wptr_gray(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[6]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \sync_out_xhdl1[11]\ : SLE
      port map(D => \sync_int[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(11));
    
    \sync_int[13]\ : SLE
      port map(D => wptr_gray(13), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[13]_net_1\);
    
    \sync_int[3]\ : SLE
      port map(D => wptr_gray(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[3]_net_1\);
    
    \sync_int[12]\ : SLE
      port map(D => wptr_gray(12), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[12]_net_1\);
    
    \sync_out_xhdl1[4]\ : SLE
      port map(D => \sync_int[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(4));
    
    \sync_int[0]\ : SLE
      port map(D => wptr_gray(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[0]_net_1\);
    
    \sync_out_xhdl1[1]\ : SLE
      port map(D => \sync_int[1]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(1));
    
    \sync_int[5]\ : SLE
      port map(D => wptr_gray(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[5]_net_1\);
    
    \sync_int[2]\ : SLE
      port map(D => wptr_gray(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[2]_net_1\);
    
    \sync_out_xhdl1[12]\ : SLE
      port map(D => \sync_int[12]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(12));
    
    \sync_out_xhdl1[9]\ : SLE
      port map(D => \sync_int[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(9));
    
    \sync_out_xhdl1[2]\ : SLE
      port map(D => \sync_int[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(2));
    
    \sync_int[8]\ : SLE
      port map(D => wptr_gray(8), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[8]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sync_out_xhdl1[7]\ : SLE
      port map(D => \sync_int[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(7));
    
    \sync_out_xhdl1[5]\ : SLE
      port map(D => \sync_int[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(5));
    
    \sync_out_xhdl1[0]\ : SLE
      port map(D => \sync_int[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(0));
    
    \sync_out_xhdl1[8]\ : SLE
      port map(D => \sync_int[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(8));
    
    \sync_int[7]\ : SLE
      port map(D => wptr_gray(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[7]_net_1\);
    
    \sync_int[10]\ : SLE
      port map(D => wptr_gray(10), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[10]_net_1\);
    
    \sync_out_xhdl1[13]\ : SLE
      port map(D => \sync_int[13]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_bin_sync_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_1 is

    port( rptr_gray           : in    std_logic_vector(13 downto 0);
          rptr_gray_sync      : out   std_logic_vector(12 downto 0);
          rptr_bin_sync_0     : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          irx_fifo_rst_i      : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_1;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_1 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \sync_int[13]_net_1\, GND_net_1, 
        \sync_int[12]_net_1\, \sync_int[0]_net_1\, 
        \sync_int[1]_net_1\, \sync_int[2]_net_1\, 
        \sync_int[3]_net_1\, \sync_int[4]_net_1\, 
        \sync_int[5]_net_1\, \sync_int[6]_net_1\, 
        \sync_int[7]_net_1\, \sync_int[8]_net_1\, 
        \sync_int[9]_net_1\, \sync_int[10]_net_1\, 
        \sync_int[11]_net_1\ : std_logic;

begin 


    \sync_int[9]\ : SLE
      port map(D => rptr_gray(9), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[9]_net_1\);
    
    \sync_int[4]\ : SLE
      port map(D => rptr_gray(4), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[4]_net_1\);
    
    \sync_out_xhdl1[10]\ : SLE
      port map(D => \sync_int[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(10));
    
    \sync_int[1]\ : SLE
      port map(D => rptr_gray(1), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[1]_net_1\);
    
    \sync_int[11]\ : SLE
      port map(D => rptr_gray(11), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[11]_net_1\);
    
    \sync_out_xhdl1[6]\ : SLE
      port map(D => \sync_int[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(6));
    
    \sync_out_xhdl1[3]\ : SLE
      port map(D => \sync_int[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(3));
    
    \sync_int[6]\ : SLE
      port map(D => rptr_gray(6), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[6]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \sync_out_xhdl1[11]\ : SLE
      port map(D => \sync_int[11]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(11));
    
    \sync_int[13]\ : SLE
      port map(D => rptr_gray(13), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[13]_net_1\);
    
    \sync_int[3]\ : SLE
      port map(D => rptr_gray(3), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[3]_net_1\);
    
    \sync_int[12]\ : SLE
      port map(D => rptr_gray(12), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[12]_net_1\);
    
    \sync_out_xhdl1[4]\ : SLE
      port map(D => \sync_int[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(4));
    
    \sync_int[0]\ : SLE
      port map(D => rptr_gray(0), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[0]_net_1\);
    
    \sync_out_xhdl1[1]\ : SLE
      port map(D => \sync_int[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(1));
    
    \sync_int[5]\ : SLE
      port map(D => rptr_gray(5), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[5]_net_1\);
    
    \sync_int[2]\ : SLE
      port map(D => rptr_gray(2), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[2]_net_1\);
    
    \sync_out_xhdl1[12]\ : SLE
      port map(D => \sync_int[12]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(12));
    
    \sync_out_xhdl1[9]\ : SLE
      port map(D => \sync_int[9]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(9));
    
    \sync_out_xhdl1[2]\ : SLE
      port map(D => \sync_int[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(2));
    
    \sync_int[8]\ : SLE
      port map(D => rptr_gray(8), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[8]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sync_out_xhdl1[7]\ : SLE
      port map(D => \sync_int[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(7));
    
    \sync_out_xhdl1[5]\ : SLE
      port map(D => \sync_int[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(5));
    
    \sync_out_xhdl1[0]\ : SLE
      port map(D => \sync_int[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(0));
    
    \sync_out_xhdl1[8]\ : SLE
      port map(D => \sync_int[8]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(8));
    
    \sync_int[7]\ : SLE
      port map(D => rptr_gray(7), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[7]_net_1\);
    
    \sync_int[10]\ : SLE
      port map(D => rptr_gray(10), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[10]_net_1\);
    
    \sync_out_xhdl1[13]\ : SLE
      port map(D => \sync_int[13]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_bin_sync_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_3 is

    port( rptr_bin_sync  : inout std_logic_vector(13 downto 0) := (others => 'Z');
          rptr_gray_sync : in    std_logic_vector(12 downto 0);
          bin_N_6_i      : out   std_logic;
          bin_N_4_0_i    : out   std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_3;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_3 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \bin_m5_5\, \bin_m5_4\, \bin_m3_0_3\, \bin_N_4_0_i\, 
        GND_net_1, VCC_net_1 : std_logic;

begin 

    bin_N_4_0_i <= \bin_N_4_0_i\;

    bin_m5_4 : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(4), B => rptr_gray_sync(6), C
         => rptr_gray_sync(5), D => rptr_gray_sync(10), Y => 
        \bin_m5_4\);
    
    \bin_out_xhdl1_0_a2[10]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(12), B => rptr_gray_sync(10), 
        C => rptr_gray_sync(11), D => rptr_bin_sync(13), Y => 
        rptr_bin_sync(10));
    
    \bin_out_xhdl1_0_a2[8]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(8), B => rptr_gray_sync(9), C
         => rptr_bin_sync(10), Y => rptr_bin_sync(8));
    
    bin_m5_5 : CFG4
      generic map(INIT => x"9669")

      port map(A => rptr_gray_sync(8), B => rptr_gray_sync(9), C
         => rptr_gray_sync(7), D => rptr_gray_sync(11), Y => 
        \bin_m5_5\);
    
    bin_m3_0_3 : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(7), B => rptr_gray_sync(9), C
         => rptr_gray_sync(6), D => rptr_gray_sync(10), Y => 
        \bin_m3_0_3\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \bin_out_xhdl1_0_a2[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(3), B => rptr_gray_sync(2), Y
         => rptr_bin_sync(2));
    
    \bin_out_xhdl1_i_o2_RNI2LPC1[12]\ : CFG3
      generic map(INIT => x"69")

      port map(A => \bin_m5_5\, B => \bin_m5_4\, C => 
        rptr_bin_sync(12), Y => bin_N_6_i);
    
    \bin_out_xhdl1_0_a2[1]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(1), B => rptr_gray_sync(2), C
         => rptr_bin_sync(3), Y => rptr_bin_sync(1));
    
    \bin_out_xhdl1_0_a2[0]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(1), B => rptr_gray_sync(0), C
         => rptr_bin_sync(3), D => rptr_gray_sync(2), Y => 
        rptr_bin_sync(0));
    
    \bin_out_xhdl1_i_o2_RNIHO211[12]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(8), B => rptr_gray_sync(11), C
         => rptr_bin_sync(12), D => \bin_m3_0_3\, Y => 
        \bin_N_4_0_i\);
    
    \bin_out_xhdl1_i_o2[11]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(11), B => rptr_bin_sync(13), C
         => rptr_gray_sync(12), Y => rptr_bin_sync(11));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \bin_out_xhdl1_0_a2[7]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(9), B => rptr_bin_sync(10), C
         => rptr_gray_sync(7), D => rptr_gray_sync(8), Y => 
        rptr_bin_sync(7));
    
    \bin_out_xhdl1_0_a2[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \bin_N_4_0_i\, B => rptr_gray_sync(5), Y => 
        rptr_bin_sync(5));
    
    \bin_out_xhdl1_i_o2[12]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(13), B => rptr_gray_sync(12), Y
         => rptr_bin_sync(12));
    
    \bin_out_xhdl1_0_a2[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(10), B => rptr_gray_sync(9), Y
         => rptr_bin_sync(9));
    
    \bin_out_xhdl1_0_a2[3]\ : CFG4
      generic map(INIT => x"9669")

      port map(A => rptr_bin_sync(12), B => \bin_m5_5\, C => 
        rptr_gray_sync(3), D => \bin_m5_4\, Y => rptr_bin_sync(3));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_1 is

    port( fifo_MEMRADDR             : out   std_logic_vector(12 downto 0);
          fifo_MEMWADDR             : out   std_logic_vector(12 downto 0);
          iRX_FIFO_wr_en_0_0        : in    std_logic;
          iRX_FIFO_rd_en_0          : in    std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          RX_FIFO_TxColDetDis_wr_en : in    std_logic;
          fifo_MEMRE                : out   std_logic;
          fifo_MEMWE                : out   std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          irx_fifo_rst_i            : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_1;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_1 is 

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_4
    port( wptr_bin_sync  : inout   std_logic_vector(13 downto 0);
          wptr_gray_sync : in    std_logic_vector(12 downto 0) := (others => 'U')
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_2
    port( wptr_gray                 : in    std_logic_vector(13 downto 0) := (others => 'U');
          wptr_gray_sync            : out   std_logic_vector(12 downto 0);
          wptr_bin_sync_0           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          irx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_1
    port( rptr_gray           : in    std_logic_vector(13 downto 0) := (others => 'U');
          rptr_gray_sync      : out   std_logic_vector(12 downto 0);
          rptr_bin_sync_0     : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          irx_fifo_rst_i      : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_3
    port( rptr_bin_sync  : inout   std_logic_vector(13 downto 0);
          rptr_gray_sync : in    std_logic_vector(12 downto 0) := (others => 'U');
          bin_N_6_i      : out   std_logic;
          bin_N_4_0_i    : out   std_logic
        );
  end component;

    signal \rptr[0]_net_1\, \rptr_s[0]\, \wptr[0]_net_1\, 
        \wptr_s[0]\, \fifo_MEMRADDR[0]\, \fifo_MEMRADDR_i[0]\, 
        \fifo_MEMWADDR[0]\, \fifo_MEMWADDR_i[0]\, 
        \rptr_gray[1]_net_1\, VCC_net_1, \rptr_gray_1[1]_net_1\, 
        GND_net_1, \rptr_gray[2]_net_1\, \rptr_gray_1[2]_net_1\, 
        \rptr_gray[3]_net_1\, \rptr_gray_1[3]_net_1\, 
        \rptr_gray[4]_net_1\, \rptr_gray_1[4]_net_1\, 
        \rptr_gray[5]_net_1\, \rptr_gray_1[5]_net_1\, 
        \rptr_gray[6]_net_1\, \rptr_gray_1[6]_net_1\, 
        \rptr_gray[7]_net_1\, \rptr_gray_1[7]_net_1\, 
        \rptr_gray[8]_net_1\, \rptr_gray_1[8]_net_1\, 
        \rptr_gray[9]_net_1\, \rptr_gray_1[9]_net_1\, 
        \rptr_gray[10]_net_1\, \rptr_gray_1[10]_net_1\, 
        \rptr_gray[11]_net_1\, \rptr_gray_1[11]_net_1\, 
        \rptr_gray[12]_net_1\, \rptr_gray_1[12]_net_1\, 
        \rptr_gray[13]_net_1\, \rptr[13]_net_1\, 
        \wptr_gray[0]_net_1\, \wptr_gray_1[0]_net_1\, 
        \wptr_gray[1]_net_1\, \wptr_gray_1[1]_net_1\, 
        \wptr_gray[2]_net_1\, \wptr_gray_1[2]_net_1\, 
        \wptr_gray[3]_net_1\, \wptr_gray_1[3]_net_1\, 
        \wptr_gray[4]_net_1\, \wptr_gray_1[4]_net_1\, 
        \wptr_gray[5]_net_1\, \wptr_gray_1[5]_net_1\, 
        \wptr_gray[6]_net_1\, \wptr_gray_1[6]_net_1\, 
        \wptr_gray[7]_net_1\, \wptr_gray_1[7]_net_1\, 
        \wptr_gray[8]_net_1\, \wptr_gray_1[8]_net_1\, 
        \wptr_gray[9]_net_1\, \wptr_gray_1[9]_net_1\, 
        \wptr_gray[10]_net_1\, \wptr_gray_1[10]_net_1\, 
        \wptr_gray[11]_net_1\, \wptr_gray_1[11]_net_1\, 
        \wptr_gray[12]_net_1\, \wptr_gray_1[12]_net_1\, 
        \wptr_gray[13]_net_1\, \wptr[13]_net_1\, 
        \rptr_gray[0]_net_1\, \rptr_gray_1[0]_net_1\, rdiff_bus, 
        \wptr_bin_sync[0]\, \wptr_bin_sync2[1]_net_1\, 
        \wptr_bin_sync[1]\, \wptr_bin_sync2[2]_net_1\, 
        \wptr_bin_sync[2]\, \wptr_bin_sync2[3]_net_1\, 
        \wptr_bin_sync[3]\, \wptr_bin_sync2[4]_net_1\, 
        \wptr_bin_sync[4]\, \wptr_bin_sync2[5]_net_1\, 
        \wptr_bin_sync[5]\, \wptr_bin_sync2[6]_net_1\, 
        \wptr_bin_sync[6]\, \wptr_bin_sync2[7]_net_1\, 
        \wptr_bin_sync[7]\, \wptr_bin_sync2[8]_net_1\, 
        \wptr_bin_sync[8]\, \wptr_bin_sync2[9]_net_1\, 
        \wptr_bin_sync[9]\, \wptr_bin_sync2[10]_net_1\, 
        \wptr_bin_sync[10]\, \wptr_bin_sync2[11]_net_1\, 
        \wptr_bin_sync[11]\, \wptr_bin_sync2[12]_net_1\, 
        \wptr_bin_sync[12]\, \wptr_bin_sync2[13]_net_1\, 
        \wptr_bin_sync[13]\, \rptr_bin_sync2[9]_net_1\, 
        \rptr_bin_sync[9]\, \rptr_bin_sync2[10]_net_1\, 
        \rptr_bin_sync[10]\, \rptr_bin_sync2[11]_net_1\, 
        \rptr_bin_sync[11]\, \rptr_bin_sync2[12]_net_1\, 
        \rptr_bin_sync[12]\, \rptr_bin_sync2[13]_net_1\, 
        \rptr_bin_sync[13]\, \fifo_MEMWADDR[7]\, 
        \memwaddr_r_2[7]_net_1\, \fifo_MEMWE\, \fifo_MEMWADDR[8]\, 
        \memwaddr_r_2[8]_net_1\, \fifo_MEMWADDR[9]\, 
        \memwaddr_r_2[9]_net_1\, \fifo_MEMWADDR[10]\, 
        \memwaddr_r_2[10]_net_1\, \fifo_MEMWADDR[11]\, 
        \memwaddr_r_2[11]_net_1\, \fifo_MEMWADDR[12]\, 
        \memwaddr_r_2[12]_net_1\, \rptr_bin_sync2[0]_net_1\, 
        \rptr_bin_sync[0]\, \rptr_bin_sync2[1]_net_1\, 
        \rptr_bin_sync[1]\, \rptr_bin_sync2[2]_net_1\, 
        \rptr_bin_sync[2]\, \rptr_bin_sync2[3]_net_1\, 
        \rptr_bin_sync[3]\, \rptr_bin_sync2[4]_net_1\, bin_N_6_i, 
        \rptr_bin_sync2[5]_net_1\, \rptr_bin_sync[5]\, 
        \rptr_bin_sync2[6]_net_1\, bin_N_4_0_i, 
        \rptr_bin_sync2[7]_net_1\, \rptr_bin_sync[7]\, 
        \rptr_bin_sync2[8]_net_1\, \rptr_bin_sync[8]\, 
        \fifo_MEMRADDR[5]\, \memraddr_r_2[5]_net_1\, \fifo_MEMRE\, 
        \fifo_MEMRADDR[6]\, un1_memraddr_r_cry_6_S_1, 
        \fifo_MEMRADDR[7]\, \memraddr_r_2[7]_net_1\, 
        \fifo_MEMRADDR[8]\, \memraddr_r_2[8]_net_1\, 
        \fifo_MEMRADDR[9]\, \memraddr_r_2[9]_net_1\, 
        \fifo_MEMRADDR[10]\, \memraddr_r_2[10]_net_1\, 
        \fifo_MEMRADDR[11]\, \memraddr_r_2[11]_net_1\, 
        \fifo_MEMRADDR[12]\, \memraddr_r_2[12]_net_1\, 
        \fifo_MEMWADDR[1]\, un1_memwaddr_r_cry_1_S_1, 
        \fifo_MEMWADDR[2]\, un1_memwaddr_r_cry_2_S_1, 
        \fifo_MEMWADDR[3]\, un1_memwaddr_r_cry_3_S_1, 
        \fifo_MEMWADDR[4]\, un1_memwaddr_r_cry_4_S_1, 
        \fifo_MEMWADDR[5]\, \memwaddr_r_2[5]_net_1\, 
        \fifo_MEMWADDR[6]\, un1_memwaddr_r_cry_6_S_1, 
        \fifo_MEMRADDR[1]\, un1_memraddr_r_cry_1_S_1, 
        \fifo_MEMRADDR[2]\, un1_memraddr_r_cry_2_S_1, 
        \fifo_MEMRADDR[3]\, un1_memraddr_r_cry_3_S_1, 
        \fifo_MEMRADDR[4]\, un1_memraddr_r_cry_4_S_1, 
        \iRX_FIFO_Full_0\, fulli, N_6_i, N_5_i, 
        \iRX_FIFO_Empty_0\, empty_r_3, \wptr[1]_net_1\, 
        \wptr_s[1]\, \wptr[2]_net_1\, \wptr_s[2]\, 
        \wptr[3]_net_1\, \wptr_s[3]\, \wptr[4]_net_1\, 
        \wptr_s[4]\, \wptr[5]_net_1\, \wptr_s[5]\, 
        \wptr[6]_net_1\, \wptr_s[6]\, \wptr[7]_net_1\, 
        \wptr_s[7]\, \wptr[8]_net_1\, \wptr_s[8]\, 
        \wptr[9]_net_1\, \wptr_s[9]\, \wptr[10]_net_1\, 
        \wptr_s[10]\, \wptr[11]_net_1\, \wptr_s[11]\, 
        \wptr[12]_net_1\, \wptr_s[12]\, \wptr_s[13]_net_1\, 
        \rptr[1]_net_1\, \rptr_s[1]\, \rptr[2]_net_1\, 
        \rptr_s[2]\, \rptr[3]_net_1\, \rptr_s[3]\, 
        \rptr[4]_net_1\, \rptr_s[4]\, \rptr[5]_net_1\, 
        \rptr_s[5]\, \rptr[6]_net_1\, \rptr_s[6]\, 
        \rptr[7]_net_1\, \rptr_s[7]\, \rptr[8]_net_1\, 
        \rptr_s[8]\, \rptr[9]_net_1\, \rptr_s[9]\, 
        \rptr[10]_net_1\, \rptr_s[10]\, \rptr[11]_net_1\, 
        \rptr_s[11]\, \rptr[12]_net_1\, \rptr_s[12]\, 
        \rptr_s[13]_net_1\, \rdiff_bus_cry_0\, 
        rdiff_bus_cry_0_Y_2, \rdiff_bus_cry_1\, \rdiff_bus[1]\, 
        \rdiff_bus_cry_2\, \rdiff_bus[2]\, \rdiff_bus_cry_3\, 
        \rdiff_bus[3]\, \rdiff_bus_cry_4\, \rdiff_bus[4]\, 
        \rdiff_bus_cry_5\, \rdiff_bus[5]\, \rdiff_bus_cry_6\, 
        \rdiff_bus[6]\, \rdiff_bus_cry_7\, \rdiff_bus[7]\, 
        \rdiff_bus_cry_8\, \rdiff_bus[8]\, \rdiff_bus_cry_9\, 
        \rdiff_bus[9]\, \rdiff_bus_cry_10\, \rdiff_bus[10]\, 
        \rdiff_bus_cry_11\, \rdiff_bus[11]\, \rdiff_bus[13]\, 
        \rdiff_bus_cry_12\, \rdiff_bus[12]\, \wdiff_bus_cry_0\, 
        wdiff_bus_cry_0_Y_2, \wdiff_bus_cry_1\, \wdiff_bus[1]\, 
        \wdiff_bus_cry_2\, \wdiff_bus[2]\, \wdiff_bus_cry_3\, 
        \wdiff_bus[3]\, \wdiff_bus_cry_4\, \wdiff_bus[4]\, 
        \wdiff_bus_cry_5\, \wdiff_bus[5]\, \wdiff_bus_cry_6\, 
        \wdiff_bus[6]\, \wdiff_bus_cry_7\, \wdiff_bus[7]\, 
        \wdiff_bus_cry_8\, \wdiff_bus[8]\, \wdiff_bus_cry_9\, 
        \wdiff_bus[9]\, \wdiff_bus_cry_10\, \wdiff_bus[10]\, 
        \wdiff_bus_cry_11\, \wdiff_bus[11]\, \wdiff_bus[13]\, 
        \wdiff_bus_cry_12\, \wdiff_bus[12]\, rptr_s_904_FCO, 
        \rptr_cry[1]_net_1\, \rptr_cry[2]_net_1\, 
        \rptr_cry[3]_net_1\, \rptr_cry[4]_net_1\, 
        \rptr_cry[5]_net_1\, \rptr_cry[6]_net_1\, 
        \rptr_cry[7]_net_1\, \rptr_cry[8]_net_1\, 
        \rptr_cry[9]_net_1\, \rptr_cry[10]_net_1\, 
        \rptr_cry[11]_net_1\, \rptr_cry[12]_net_1\, 
        wptr_s_905_FCO, \wptr_cry[1]_net_1\, \wptr_cry[2]_net_1\, 
        \wptr_cry[3]_net_1\, \wptr_cry[4]_net_1\, 
        \wptr_cry[5]_net_1\, \wptr_cry[6]_net_1\, 
        \wptr_cry[7]_net_1\, \wptr_cry[8]_net_1\, 
        \wptr_cry[9]_net_1\, \wptr_cry[10]_net_1\, 
        \wptr_cry[11]_net_1\, \wptr_cry[12]_net_1\, 
        un1_memraddr_r_s_1_927_FCO, \un1_memraddr_r_cry_1\, 
        \un1_memraddr_r_cry_2\, \un1_memraddr_r_cry_3\, 
        \un1_memraddr_r_cry_4\, \un1_memraddr_r_cry_5\, 
        un1_memraddr_r_cry_5_S_1, \un1_memraddr_r_cry_6\, 
        \un1_memraddr_r_cry_7\, un1_memraddr_r_cry_7_S_1, 
        \un1_memraddr_r_cry_8\, un1_memraddr_r_cry_8_S_1, 
        \un1_memraddr_r_cry_9\, un1_memraddr_r_cry_9_S_1, 
        \un1_memraddr_r_cry_10\, un1_memraddr_r_cry_10_S_1, 
        un1_memraddr_r_s_12_S_1, \un1_memraddr_r_cry_11\, 
        un1_memraddr_r_cry_11_S_1, un1_memwaddr_r_s_1_928_FCO, 
        \un1_memwaddr_r_cry_1\, \un1_memwaddr_r_cry_2\, 
        \un1_memwaddr_r_cry_3\, \un1_memwaddr_r_cry_4\, 
        \un1_memwaddr_r_cry_5\, un1_memwaddr_r_cry_5_S_1, 
        \un1_memwaddr_r_cry_6\, \un1_memwaddr_r_cry_7\, 
        un1_memwaddr_r_cry_7_S_1, \un1_memwaddr_r_cry_8\, 
        un1_memwaddr_r_cry_8_S_1, \un1_memwaddr_r_cry_9\, 
        un1_memwaddr_r_cry_9_S_1, \un1_memwaddr_r_cry_10\, 
        un1_memwaddr_r_cry_10_S_1, un1_memwaddr_r_s_12_S_1, 
        \un1_memwaddr_r_cry_11\, un1_memwaddr_r_cry_11_S_1, 
        \fulli_0_1\, N_12, \fulli_0_a3_3\, empty_r_3_0_a2_3, 
        un4_we_i_0, un4_re_i_0, empty_r_3_0_a2_9, un4_we_i_8, 
        un4_we_i_7, un4_re_i_8, un4_re_i_7, empty_r_3_0_a2_11, 
        un4_we_i_9, un4_re_i_9, N_7, \fulli_0_a3_0_3\, 
        empty_r_3_0_a2_7, \wptr_gray_sync[0]\, 
        \wptr_gray_sync[1]\, \wptr_gray_sync[2]\, 
        \wptr_gray_sync[3]\, \wptr_gray_sync[4]\, 
        \wptr_gray_sync[5]\, \wptr_gray_sync[6]\, 
        \wptr_gray_sync[7]\, \wptr_gray_sync[8]\, 
        \wptr_gray_sync[9]\, \wptr_gray_sync[10]\, 
        \wptr_gray_sync[11]\, \wptr_gray_sync[12]\, 
        \rptr_gray_sync[0]\, \rptr_gray_sync[1]\, 
        \rptr_gray_sync[2]\, \rptr_gray_sync[3]\, 
        \rptr_gray_sync[4]\, \rptr_gray_sync[5]\, 
        \rptr_gray_sync[6]\, \rptr_gray_sync[7]\, 
        \rptr_gray_sync[8]\, \rptr_gray_sync[9]\, 
        \rptr_gray_sync[10]\, \rptr_gray_sync[11]\, 
        \rptr_gray_sync[12]\ : std_logic;
    signal nc2, nc1 : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_4
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_4(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_2
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_2(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_1
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_1(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_3
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_3(DEF_ARCH);
begin 

    fifo_MEMRADDR(12) <= \fifo_MEMRADDR[12]\;
    fifo_MEMRADDR(11) <= \fifo_MEMRADDR[11]\;
    fifo_MEMRADDR(10) <= \fifo_MEMRADDR[10]\;
    fifo_MEMRADDR(9) <= \fifo_MEMRADDR[9]\;
    fifo_MEMRADDR(8) <= \fifo_MEMRADDR[8]\;
    fifo_MEMRADDR(7) <= \fifo_MEMRADDR[7]\;
    fifo_MEMRADDR(6) <= \fifo_MEMRADDR[6]\;
    fifo_MEMRADDR(5) <= \fifo_MEMRADDR[5]\;
    fifo_MEMRADDR(4) <= \fifo_MEMRADDR[4]\;
    fifo_MEMRADDR(3) <= \fifo_MEMRADDR[3]\;
    fifo_MEMRADDR(2) <= \fifo_MEMRADDR[2]\;
    fifo_MEMRADDR(1) <= \fifo_MEMRADDR[1]\;
    fifo_MEMRADDR(0) <= \fifo_MEMRADDR[0]\;
    fifo_MEMWADDR(12) <= \fifo_MEMWADDR[12]\;
    fifo_MEMWADDR(11) <= \fifo_MEMWADDR[11]\;
    fifo_MEMWADDR(10) <= \fifo_MEMWADDR[10]\;
    fifo_MEMWADDR(9) <= \fifo_MEMWADDR[9]\;
    fifo_MEMWADDR(8) <= \fifo_MEMWADDR[8]\;
    fifo_MEMWADDR(7) <= \fifo_MEMWADDR[7]\;
    fifo_MEMWADDR(6) <= \fifo_MEMWADDR[6]\;
    fifo_MEMWADDR(5) <= \fifo_MEMWADDR[5]\;
    fifo_MEMWADDR(4) <= \fifo_MEMWADDR[4]\;
    fifo_MEMWADDR(3) <= \fifo_MEMWADDR[3]\;
    fifo_MEMWADDR(2) <= \fifo_MEMWADDR[2]\;
    fifo_MEMWADDR(1) <= \fifo_MEMWADDR[1]\;
    fifo_MEMWADDR(0) <= \fifo_MEMWADDR[0]\;
    iRX_FIFO_Empty_0 <= \iRX_FIFO_Empty_0\;
    iRX_FIFO_Full_0 <= \iRX_FIFO_Full_0\;
    fifo_MEMRE <= \fifo_MEMRE\;
    fifo_MEMWE <= \fifo_MEMWE\;

    \rptr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[4]_net_1\, S
         => \rptr_s[5]\, Y => OPEN, FCO => \rptr_cry[5]_net_1\);
    
    \memwaddr_r_2[9]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_9_S_1, D => un4_we_i_9, Y => 
        \memwaddr_r_2[9]_net_1\);
    
    wdiff_bus_cry_8 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[8]_net_1\, B => 
        \rptr_bin_sync2[8]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_7\, S => \wdiff_bus[8]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_8\);
    
    \wptr_bin_sync2[12]\ : SLE
      port map(D => \wptr_bin_sync[12]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[12]_net_1\);
    
    \L1.empty_r_3_0_a2_11\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \rdiff_bus[4]\, B => \rdiff_bus[5]\, C => 
        empty_r_3_0_a2_3, D => empty_r_3_0_a2_9, Y => 
        empty_r_3_0_a2_11);
    
    wdiff_bus_cry_11 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[11]_net_1\, B => 
        \rptr_bin_sync2[11]_net_1\, C => GND_net_1, D => 
        GND_net_1, FCI => \wdiff_bus_cry_10\, S => 
        \wdiff_bus[11]\, Y => OPEN, FCO => \wdiff_bus_cry_11\);
    
    \wptr_gray[4]\ : SLE
      port map(D => \wptr_gray_1[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[4]_net_1\);
    
    \rptr_gray_1[3]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[3]_net_1\, B => \rptr[4]_net_1\, Y => 
        \rptr_gray_1[3]_net_1\);
    
    \rptr_bin_sync2[6]\ : SLE
      port map(D => bin_N_4_0_i, CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_bin_sync2[6]_net_1\);
    
    \rptr[1]\ : SLE
      port map(D => \rptr_s[1]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[1]_net_1\);
    
    fulli_0_a3_0_3 : CFG4
      generic map(INIT => x"8000")

      port map(A => \wdiff_bus[2]\, B => 
        RX_FIFO_TxColDetDis_wr_en, C => iRX_FIFO_wr_en_0_0, D => 
        \wdiff_bus[3]\, Y => \fulli_0_a3_0_3\);
    
    un1_memraddr_r_s_1_927 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[0]\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => un1_memraddr_r_s_1_927_FCO);
    
    \wptr_gray_1[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[9]_net_1\, B => \wptr[10]_net_1\, Y => 
        \wptr_gray_1[9]_net_1\);
    
    \rptr_gray_1[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[5]_net_1\, B => \rptr[6]_net_1\, Y => 
        \rptr_gray_1[5]_net_1\);
    
    \rptr_gray[9]\ : SLE
      port map(D => \rptr_gray_1[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[9]_net_1\);
    
    un1_memwaddr_r_cry_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_6\, 
        S => un1_memwaddr_r_cry_7_S_1, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_7\);
    
    \rptr_gray[8]\ : SLE
      port map(D => \rptr_gray_1[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[8]_net_1\);
    
    un1_memraddr_r_cry_11 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[11]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_10\, 
        S => un1_memraddr_r_cry_11_S_1, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_11\);
    
    \rptr_gray_1[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[2]_net_1\, B => \rptr[3]_net_1\, Y => 
        \rptr_gray_1[2]_net_1\);
    
    \rptr_bin_sync2[7]\ : SLE
      port map(D => \rptr_bin_sync[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[7]_net_1\);
    
    \memwaddr_r[1]\ : SLE
      port map(D => un1_memwaddr_r_cry_1_S_1, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[1]\);
    
    \wptr_gray_1[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[7]_net_1\, B => \wptr[8]_net_1\, Y => 
        \wptr_gray_1[7]_net_1\);
    
    \rptr_gray[13]\ : SLE
      port map(D => \rptr[13]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[13]_net_1\);
    
    \memraddr_r[0]\ : SLE
      port map(D => \fifo_MEMRADDR_i[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[0]\);
    
    \memraddr_r_2[9]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => 
        un1_memraddr_r_cry_9_S_1, D => un4_re_i_9, Y => 
        \memraddr_r_2[9]_net_1\);
    
    \wptr[0]\ : SLE
      port map(D => \wptr_s[0]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[0]_net_1\);
    
    \rptr_bin_sync2[8]\ : SLE
      port map(D => \rptr_bin_sync[8]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[8]_net_1\);
    
    \rptr_gray_1[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[1]_net_1\, B => \rptr[2]_net_1\, Y => 
        \rptr_gray_1[1]_net_1\);
    
    \rptr_gray[10]\ : SLE
      port map(D => \rptr_gray_1[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[10]_net_1\);
    
    \wptr_gray_1[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[0]_net_1\, B => \wptr[1]_net_1\, Y => 
        \wptr_gray_1[0]_net_1\);
    
    wdiff_bus_cry_9 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[9]_net_1\, B => 
        \rptr_bin_sync2[9]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_8\, S => \wdiff_bus[9]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_9\);
    
    \rptr[5]\ : SLE
      port map(D => \rptr_s[5]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[5]_net_1\);
    
    \rptr_gray[3]\ : SLE
      port map(D => \rptr_gray_1[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[3]_net_1\);
    
    \rptr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[5]_net_1\, S
         => \rptr_s[6]\, Y => OPEN, FCO => \rptr_cry[6]_net_1\);
    
    \wptr_gray[3]\ : SLE
      port map(D => \wptr_gray_1[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[3]_net_1\);
    
    \rptr_gray_1[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[10]_net_1\, B => \rptr[11]_net_1\, Y
         => \rptr_gray_1[10]_net_1\);
    
    un1_memraddr_r_cry_10 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_9\, 
        S => un1_memraddr_r_cry_10_S_1, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_10\);
    
    \rptr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[7]_net_1\, S
         => \rptr_s[8]\, Y => OPEN, FCO => \rptr_cry[8]_net_1\);
    
    \rptr[7]\ : SLE
      port map(D => \rptr_s[7]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[7]_net_1\);
    
    rdiff_bus_cry_4 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[4]_net_1\, B => 
        \rptr[4]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_3\, S => \rdiff_bus[4]\, Y => OPEN, FCO
         => \rdiff_bus_cry_4\);
    
    \rptr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[9]_net_1\, S
         => \rptr_s[10]\, Y => OPEN, FCO => \rptr_cry[10]_net_1\);
    
    \rptr_bin_sync2[12]\ : SLE
      port map(D => \rptr_bin_sync[12]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[12]_net_1\);
    
    memwe_0_a3 : CFG3
      generic map(INIT => x"20")

      port map(A => RX_FIFO_TxColDetDis_wr_en, B => 
        \iRX_FIFO_Full_0\, C => iRX_FIFO_wr_en_0_0, Y => 
        \fifo_MEMWE\);
    
    \rptr_bin_sync2[0]\ : SLE
      port map(D => \rptr_bin_sync[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[0]_net_1\);
    
    \L1.empty_r_3_0_a2_7\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \rdiff_bus[3]\, B => \rdiff_bus[2]\, C => 
        \rdiff_bus[1]\, D => N_7, Y => empty_r_3_0_a2_7);
    
    \wptr[11]\ : SLE
      port map(D => \wptr_s[11]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[11]_net_1\);
    
    rdiff_bus_cry_1 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[1]_net_1\, B => 
        \rptr[1]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_0\, S => \rdiff_bus[1]\, Y => OPEN, FCO
         => \rdiff_bus_cry_1\);
    
    \memraddr_r[1]\ : SLE
      port map(D => un1_memraddr_r_cry_1_S_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[1]\);
    
    \L1.empty_r_3_0_a2_9\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \rdiff_bus[8]\, B => \rdiff_bus[9]\, C => 
        \rdiff_bus[10]\, D => \rdiff_bus[11]\, Y => 
        empty_r_3_0_a2_9);
    
    \rptr_bin_sync2[2]\ : SLE
      port map(D => \rptr_bin_sync[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[2]_net_1\);
    
    \memraddr_r_2[7]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => 
        un1_memraddr_r_cry_7_S_1, D => un4_re_i_9, Y => 
        \memraddr_r_2[7]_net_1\);
    
    un1_memwaddr_r_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_5\, 
        S => un1_memwaddr_r_cry_6_S_1, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_6\);
    
    rdiff_bus_cry_6 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[6]_net_1\, B => 
        \rptr[6]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_5\, S => \rdiff_bus[6]\, Y => OPEN, FCO
         => \rdiff_bus_cry_6\);
    
    \memwaddr_r_2[10]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_10_S_1, D => un4_we_i_9, Y => 
        \memwaddr_r_2[10]_net_1\);
    
    \memraddr_r_2[5]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => 
        un1_memraddr_r_cry_5_S_1, D => un4_re_i_9, Y => 
        \memraddr_r_2[5]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    un1_memwaddr_r_cry_9 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[9]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_8\, 
        S => un1_memwaddr_r_cry_9_S_1, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_9\);
    
    \rptr_gray[1]\ : SLE
      port map(D => \rptr_gray_1[1]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[1]_net_1\);
    
    \memwaddr_r[7]\ : SLE
      port map(D => \memwaddr_r_2[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[7]\);
    
    \wptr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[3]_net_1\, S
         => \wptr_s[4]\, Y => OPEN, FCO => \wptr_cry[4]_net_1\);
    
    \wptr_gray_1[12]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[13]_net_1\, B => \wptr[12]_net_1\, Y
         => \wptr_gray_1[12]_net_1\);
    
    \wptr[12]\ : SLE
      port map(D => \wptr_s[12]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[12]_net_1\);
    
    \L1.empty_r_3_0_o2\ : CFG2
      generic map(INIT => x"E")

      port map(A => rdiff_bus_cry_0_Y_2, B => iRX_FIFO_rd_en_0, Y
         => N_7);
    
    \wptr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[9]_net_1\, S
         => \wptr_s[10]\, Y => OPEN, FCO => \wptr_cry[10]_net_1\);
    
    wdiff_bus_cry_5 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[5]_net_1\, B => 
        \rptr_bin_sync2[5]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_4\, S => \wdiff_bus[5]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_5\);
    
    \rptr_gray[12]\ : SLE
      port map(D => \rptr_gray_1[12]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[12]_net_1\);
    
    \memwaddr_r[4]\ : SLE
      port map(D => un1_memwaddr_r_cry_4_S_1, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[4]\);
    
    \wptr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[1]_net_1\, S
         => \wptr_s[2]\, Y => OPEN, FCO => \wptr_cry[2]_net_1\);
    
    \memraddr_r_2[10]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => 
        un1_memraddr_r_cry_10_S_1, D => un4_re_i_9, Y => 
        \memraddr_r_2[10]_net_1\);
    
    rdiff_bus_cry_11 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[11]_net_1\, B => 
        \rptr[11]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_10\, S => \rdiff_bus[11]\, Y => OPEN, FCO
         => \rdiff_bus_cry_11\);
    
    wdiff_bus_cry_0 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[0]_net_1\, B => 
        \rptr_bin_sync2[0]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => VCC_net_1, S => OPEN, Y => wdiff_bus_cry_0_Y_2, 
        FCO => \wdiff_bus_cry_0\);
    
    \wptr[1]\ : SLE
      port map(D => \wptr_s[1]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[1]_net_1\);
    
    \rptr_bin_sync2[4]\ : SLE
      port map(D => bin_N_6_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[4]_net_1\);
    
    \wptr_bin_sync2[6]\ : SLE
      port map(D => \wptr_bin_sync[6]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[6]_net_1\);
    
    \rptr[3]\ : SLE
      port map(D => \rptr_s[3]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[3]_net_1\);
    
    \wptr_gray[13]\ : SLE
      port map(D => \wptr[13]_net_1\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr_gray[13]_net_1\);
    
    \wptr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[2]_net_1\, S
         => \wptr_s[3]\, Y => OPEN, FCO => \wptr_cry[3]_net_1\);
    
    \rptr[6]\ : SLE
      port map(D => \rptr_s[6]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[6]_net_1\);
    
    rdiff_bus_cry_8 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[8]_net_1\, B => 
        \rptr[8]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_7\, S => \rdiff_bus[8]\, Y => OPEN, FCO
         => \rdiff_bus_cry_8\);
    
    \wptr_gray[10]\ : SLE
      port map(D => \wptr_gray_1[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[10]_net_1\);
    
    rdiff_bus_cry_7 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[7]_net_1\, B => 
        \rptr[7]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_6\, S => \rdiff_bus[7]\, Y => OPEN, FCO
         => \rdiff_bus_cry_7\);
    
    \wptr_bin_sync2[7]\ : SLE
      port map(D => \wptr_bin_sync[7]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[7]_net_1\);
    
    \rptr_gray_1[11]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[11]_net_1\, B => \rptr[12]_net_1\, Y
         => \rptr_gray_1[11]_net_1\);
    
    \rptr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[8]_net_1\, S
         => \rptr_s[9]\, Y => OPEN, FCO => \rptr_cry[9]_net_1\);
    
    un1_memwaddr_r_cry_1 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[1]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        un1_memwaddr_r_s_1_928_FCO, S => un1_memwaddr_r_cry_1_S_1, 
        Y => OPEN, FCO => \un1_memwaddr_r_cry_1\);
    
    \rptr_gray[5]\ : SLE
      port map(D => \rptr_gray_1[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[5]_net_1\);
    
    un1_memwaddr_r_s_12 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[12]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_11\, 
        S => un1_memwaddr_r_s_12_S_1, Y => OPEN, FCO => OPEN);
    
    \wptr_gray_1[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[2]_net_1\, B => \wptr[3]_net_1\, Y => 
        \wptr_gray_1[2]_net_1\);
    
    \wptr[5]\ : SLE
      port map(D => \wptr_s[5]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[5]_net_1\);
    
    rdiff_bus_cry_5 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[5]_net_1\, B => 
        \rptr[5]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_4\, S => \rdiff_bus[5]\, Y => OPEN, FCO
         => \rdiff_bus_cry_5\);
    
    \wptr_bin_sync2[8]\ : SLE
      port map(D => \wptr_bin_sync[8]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[8]_net_1\);
    
    fulli_0_a3_3 : CFG4
      generic map(INIT => x"8000")

      port map(A => \wdiff_bus[7]\, B => \wdiff_bus[8]\, C => 
        \wdiff_bus[9]\, D => \wdiff_bus[10]\, Y => \fulli_0_a3_3\);
    
    \wptr[7]\ : SLE
      port map(D => \wptr_s[7]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[7]_net_1\);
    
    un1_memwaddr_r_cry_2 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[2]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_1\, 
        S => un1_memwaddr_r_cry_2_S_1, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_2\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \wptr_gray[1]\ : SLE
      port map(D => \wptr_gray_1[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[1]_net_1\);
    
    \rptr_gray_1[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[9]_net_1\, B => \rptr[10]_net_1\, Y => 
        \rptr_gray_1[9]_net_1\);
    
    \rptr_bin_sync2[5]\ : SLE
      port map(D => \rptr_bin_sync[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[5]_net_1\);
    
    \rptr_bin_sync2[1]\ : SLE
      port map(D => \rptr_bin_sync[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[1]_net_1\);
    
    \memwaddr_r[10]\ : SLE
      port map(D => \memwaddr_r_2[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[10]\);
    
    wdiff_bus_cry_7 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[7]_net_1\, B => 
        \rptr_bin_sync2[7]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_6\, S => \wdiff_bus[7]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_7\);
    
    \wptr_bin_sync2[0]\ : SLE
      port map(D => \wptr_bin_sync[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rdiff_bus);
    
    un1_memwaddr_r_cry_8 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[8]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_7\, 
        S => un1_memwaddr_r_cry_8_S_1, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_8\);
    
    \wptr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => wptr_s_905_FCO, S => 
        \wptr_s[1]\, Y => OPEN, FCO => \wptr_cry[1]_net_1\);
    
    un1_memwaddr_r_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_3\, 
        S => un1_memwaddr_r_cry_4_S_1, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_4\);
    
    un1_memwaddr_r_cry_3 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[3]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_2\, 
        S => un1_memwaddr_r_cry_3_S_1, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_3\);
    
    \memraddr_r[8]\ : SLE
      port map(D => \memraddr_r_2[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[8]\);
    
    \rptr[9]\ : SLE
      port map(D => \rptr_s[9]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[9]_net_1\);
    
    \wptr_gray_1[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[6]_net_1\, B => \wptr[7]_net_1\, Y => 
        \wptr_gray_1[6]_net_1\);
    
    \wptr_gray[12]\ : SLE
      port map(D => \wptr_gray_1[12]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[12]_net_1\);
    
    \wptr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[6]_net_1\, S
         => \wptr_s[7]\, Y => OPEN, FCO => \wptr_cry[7]_net_1\);
    
    \wptr_bin_sync2[2]\ : SLE
      port map(D => \wptr_bin_sync[2]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[2]_net_1\);
    
    fulli_0_1 : CFG4
      generic map(INIT => x"01FF")

      port map(A => \wdiff_bus[6]\, B => \wdiff_bus[5]\, C => 
        N_12, D => \fulli_0_a3_3\, Y => \fulli_0_1\);
    
    \L1.un4_re_i_9\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \fifo_MEMRADDR[4]\, B => \fifo_MEMRADDR[3]\, 
        C => \fifo_MEMRADDR[0]\, D => un4_re_i_0, Y => un4_re_i_9);
    
    un1_memraddr_r_cry_3 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[3]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_2\, 
        S => un1_memraddr_r_cry_3_S_1, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_3\);
    
    \rptr_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \rptr[0]_net_1\, Y => \rptr_s[0]\);
    
    un1_memraddr_r_cry_1 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[1]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        un1_memraddr_r_s_1_927_FCO, S => un1_memraddr_r_cry_1_S_1, 
        Y => OPEN, FCO => \un1_memraddr_r_cry_1\);
    
    \rptr[4]\ : SLE
      port map(D => \rptr_s[4]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[4]_net_1\);
    
    \memwaddr_r_2[5]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_5_S_1, D => un4_we_i_9, Y => 
        \memwaddr_r_2[5]_net_1\);
    
    \wptr_gray[6]\ : SLE
      port map(D => \wptr_gray_1[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[6]_net_1\);
    
    \wptr_gray_1[3]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[3]_net_1\, B => \wptr[4]_net_1\, Y => 
        \wptr_gray_1[3]_net_1\);
    
    \wptr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[4]_net_1\, S
         => \wptr_s[5]\, Y => OPEN, FCO => \wptr_cry[5]_net_1\);
    
    un1_memraddr_r_cry_9 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[9]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_8\, 
        S => un1_memraddr_r_cry_9_S_1, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_9\);
    
    fulli_0_a3_0 : CFG4
      generic map(INIT => x"4000")

      port map(A => wdiff_bus_cry_0_Y_2, B => \wdiff_bus[1]\, C
         => \wdiff_bus[4]\, D => \fulli_0_a3_0_3\, Y => N_12);
    
    \rptr_gray[4]\ : SLE
      port map(D => \rptr_gray_1[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[4]_net_1\);
    
    un1_memraddr_r_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_4\, 
        S => un1_memraddr_r_cry_5_S_1, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_5\);
    
    \wptr_bin_sync2[4]\ : SLE
      port map(D => \wptr_bin_sync[4]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[4]_net_1\);
    
    \wptr[3]\ : SLE
      port map(D => \wptr_s[3]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[3]_net_1\);
    
    \L1.un4_we_i_9\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \fifo_MEMWADDR[4]\, B => \fifo_MEMWADDR[3]\, 
        C => \fifo_MEMWADDR[0]\, D => un4_we_i_0, Y => un4_we_i_9);
    
    \memwaddr_r[6]\ : SLE
      port map(D => un1_memwaddr_r_cry_6_S_1, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[6]\);
    
    \wptr[6]\ : SLE
      port map(D => \wptr_s[6]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[6]_net_1\);
    
    \memwaddr_r[9]\ : SLE
      port map(D => \memwaddr_r_2[9]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[9]\);
    
    \memraddr_r[10]\ : SLE
      port map(D => \memraddr_r_2[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[10]\);
    
    \L1.un4_re_i_8\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \fifo_MEMRADDR[10]\, B => \fifo_MEMRADDR[9]\, 
        C => \fifo_MEMRADDR[8]\, D => \fifo_MEMRADDR[7]\, Y => 
        un4_re_i_8);
    
    \memwaddr_r[3]\ : SLE
      port map(D => un1_memwaddr_r_cry_3_S_1, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[3]\);
    
    \rptr_gray_1[12]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[13]_net_1\, B => \rptr[12]_net_1\, Y
         => \rptr_gray_1[12]_net_1\);
    
    full_r : SLE
      port map(D => fulli, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \iRX_FIFO_Full_0\);
    
    \rptr_bin_sync2[3]\ : SLE
      port map(D => \rptr_bin_sync[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[3]_net_1\);
    
    \wptr_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \wptr[0]_net_1\, Y => \wptr_s[0]\);
    
    \rptr[2]\ : SLE
      port map(D => \rptr_s[2]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[2]_net_1\);
    
    \memraddr_r[3]\ : SLE
      port map(D => un1_memraddr_r_cry_3_S_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[3]\);
    
    \wptr[13]\ : SLE
      port map(D => \wptr_s[13]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \wptr[13]_net_1\);
    
    \rptr_bin_sync2[9]\ : SLE
      port map(D => \rptr_bin_sync[9]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[9]_net_1\);
    
    \wptr_bin_sync2[13]\ : SLE
      port map(D => \wptr_bin_sync[13]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[13]_net_1\);
    
    \rptr[11]\ : SLE
      port map(D => \rptr_s[11]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rptr[11]_net_1\);
    
    \wptr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[5]_net_1\, S
         => \wptr_s[6]\, Y => OPEN, FCO => \wptr_cry[6]_net_1\);
    
    \rptr_bin_sync2[11]\ : SLE
      port map(D => \rptr_bin_sync[11]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[11]_net_1\);
    
    \wptr_bin_sync2[5]\ : SLE
      port map(D => \wptr_bin_sync[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[5]_net_1\);
    
    \L1.un4_we_i_8\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \fifo_MEMWADDR[10]\, B => \fifo_MEMWADDR[9]\, 
        C => \fifo_MEMWADDR[8]\, D => \fifo_MEMWADDR[7]\, Y => 
        un4_we_i_8);
    
    \wptr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[7]_net_1\, S
         => \wptr_s[8]\, Y => OPEN, FCO => \wptr_cry[8]_net_1\);
    
    \wptr_bin_sync2[1]\ : SLE
      port map(D => \wptr_bin_sync[1]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[1]_net_1\);
    
    Wr_corefifo_grayToBinConv : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_4
      port map(wptr_bin_sync(13) => \wptr_bin_sync[13]\, 
        wptr_bin_sync(12) => \wptr_bin_sync[12]\, 
        wptr_bin_sync(11) => \wptr_bin_sync[11]\, 
        wptr_bin_sync(10) => \wptr_bin_sync[10]\, 
        wptr_bin_sync(9) => \wptr_bin_sync[9]\, wptr_bin_sync(8)
         => \wptr_bin_sync[8]\, wptr_bin_sync(7) => 
        \wptr_bin_sync[7]\, wptr_bin_sync(6) => 
        \wptr_bin_sync[6]\, wptr_bin_sync(5) => 
        \wptr_bin_sync[5]\, wptr_bin_sync(4) => 
        \wptr_bin_sync[4]\, wptr_bin_sync(3) => 
        \wptr_bin_sync[3]\, wptr_bin_sync(2) => 
        \wptr_bin_sync[2]\, wptr_bin_sync(1) => 
        \wptr_bin_sync[1]\, wptr_bin_sync(0) => 
        \wptr_bin_sync[0]\, wptr_gray_sync(12) => 
        \wptr_gray_sync[12]\, wptr_gray_sync(11) => 
        \wptr_gray_sync[11]\, wptr_gray_sync(10) => 
        \wptr_gray_sync[10]\, wptr_gray_sync(9) => 
        \wptr_gray_sync[9]\, wptr_gray_sync(8) => 
        \wptr_gray_sync[8]\, wptr_gray_sync(7) => 
        \wptr_gray_sync[7]\, wptr_gray_sync(6) => 
        \wptr_gray_sync[6]\, wptr_gray_sync(5) => 
        \wptr_gray_sync[5]\, wptr_gray_sync(4) => 
        \wptr_gray_sync[4]\, wptr_gray_sync(3) => 
        \wptr_gray_sync[3]\, wptr_gray_sync(2) => 
        \wptr_gray_sync[2]\, wptr_gray_sync(1) => 
        \wptr_gray_sync[1]\, wptr_gray_sync(0) => 
        \wptr_gray_sync[0]\);
    
    \wptr_gray_1[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[4]_net_1\, B => \wptr[5]_net_1\, Y => 
        \wptr_gray_1[4]_net_1\);
    
    \rptr_bin_sync2[13]\ : SLE
      port map(D => \rptr_bin_sync[13]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[13]_net_1\);
    
    wptr_s_905 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => wptr_s_905_FCO);
    
    \L1.un4_re_i_7\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \fifo_MEMRADDR[12]\, B => \fifo_MEMRADDR[11]\, 
        C => \fifo_MEMRADDR[6]\, D => \fifo_MEMRADDR[5]\, Y => 
        un4_re_i_7);
    
    overflow_r : SLE
      port map(D => N_6_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        iRX_FIFO_OVERFLOW_0);
    
    fulli_0 : CFG4
      generic map(INIT => x"BAAA")

      port map(A => \wdiff_bus[13]\, B => \fulli_0_1\, C => 
        \wdiff_bus[11]\, D => \wdiff_bus[12]\, Y => fulli);
    
    \memraddr_r_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \fifo_MEMRADDR[0]\, Y => \fifo_MEMRADDR_i[0]\);
    
    \memraddr_r_2[8]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => 
        un1_memraddr_r_cry_8_S_1, D => un4_re_i_9, Y => 
        \memraddr_r_2[8]_net_1\);
    
    \rptr_gray[11]\ : SLE
      port map(D => \rptr_gray_1[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[11]_net_1\);
    
    \wptr_bin_sync2[10]\ : SLE
      port map(D => \wptr_bin_sync[10]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[10]_net_1\);
    
    \rptr[10]\ : SLE
      port map(D => \rptr_s[10]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rptr[10]_net_1\);
    
    \wptr[9]\ : SLE
      port map(D => \wptr_s[9]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[9]_net_1\);
    
    Wr_corefifo_doubleSync : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_2
      port map(wptr_gray(13) => \wptr_gray[13]_net_1\, 
        wptr_gray(12) => \wptr_gray[12]_net_1\, wptr_gray(11) => 
        \wptr_gray[11]_net_1\, wptr_gray(10) => 
        \wptr_gray[10]_net_1\, wptr_gray(9) => 
        \wptr_gray[9]_net_1\, wptr_gray(8) => 
        \wptr_gray[8]_net_1\, wptr_gray(7) => 
        \wptr_gray[7]_net_1\, wptr_gray(6) => 
        \wptr_gray[6]_net_1\, wptr_gray(5) => 
        \wptr_gray[5]_net_1\, wptr_gray(4) => 
        \wptr_gray[4]_net_1\, wptr_gray(3) => 
        \wptr_gray[3]_net_1\, wptr_gray(2) => 
        \wptr_gray[2]_net_1\, wptr_gray(1) => 
        \wptr_gray[1]_net_1\, wptr_gray(0) => 
        \wptr_gray[0]_net_1\, wptr_gray_sync(12) => 
        \wptr_gray_sync[12]\, wptr_gray_sync(11) => 
        \wptr_gray_sync[11]\, wptr_gray_sync(10) => 
        \wptr_gray_sync[10]\, wptr_gray_sync(9) => 
        \wptr_gray_sync[9]\, wptr_gray_sync(8) => 
        \wptr_gray_sync[8]\, wptr_gray_sync(7) => 
        \wptr_gray_sync[7]\, wptr_gray_sync(6) => 
        \wptr_gray_sync[6]\, wptr_gray_sync(5) => 
        \wptr_gray_sync[5]\, wptr_gray_sync(4) => 
        \wptr_gray_sync[4]\, wptr_gray_sync(3) => 
        \wptr_gray_sync[3]\, wptr_gray_sync(2) => 
        \wptr_gray_sync[2]\, wptr_gray_sync(1) => 
        \wptr_gray_sync[1]\, wptr_gray_sync(0) => 
        \wptr_gray_sync[0]\, wptr_bin_sync_0 => 
        \wptr_bin_sync[13]\, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, irx_fifo_rst_i => 
        irx_fifo_rst_i);
    
    un1_memwaddr_r_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_4\, 
        S => un1_memwaddr_r_cry_5_S_1, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_5\);
    
    \rptr_gray[0]\ : SLE
      port map(D => \rptr_gray_1[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[0]_net_1\);
    
    empty_r : SLE
      port map(D => empty_r_3, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \iRX_FIFO_Empty_0\);
    
    \memwaddr_r_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \fifo_MEMWADDR[0]\, Y => \fifo_MEMWADDR_i[0]\);
    
    \L1.empty_r_3_0_a2_3\ : CFG2
      generic map(INIT => x"1")

      port map(A => \rdiff_bus[7]\, B => \rdiff_bus[6]\, Y => 
        empty_r_3_0_a2_3);
    
    \memwaddr_r_2[12]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_s_12_S_1, D => un4_we_i_9, Y => 
        \memwaddr_r_2[12]_net_1\);
    
    un1_memwaddr_r_s_1_928 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[0]\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => un1_memwaddr_r_s_1_928_FCO);
    
    \rptr_gray_1[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[7]_net_1\, B => \rptr[8]_net_1\, Y => 
        \rptr_gray_1[7]_net_1\);
    
    un1_memraddr_r_cry_2 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[2]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_1\, 
        S => un1_memraddr_r_cry_2_S_1, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_2\);
    
    wdiff_bus_cry_12 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[12]_net_1\, B => 
        \rptr_bin_sync2[12]_net_1\, C => GND_net_1, D => 
        GND_net_1, FCI => \wdiff_bus_cry_11\, S => 
        \wdiff_bus[12]\, Y => OPEN, FCO => \wdiff_bus_cry_12\);
    
    \wptr[4]\ : SLE
      port map(D => \wptr_s[4]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[4]_net_1\);
    
    un1_memraddr_r_cry_8 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[8]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_7\, 
        S => un1_memraddr_r_cry_8_S_1, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_8\);
    
    \rptr_s[13]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[13]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[12]_net_1\, S
         => \rptr_s[13]_net_1\, Y => OPEN, FCO => OPEN);
    
    \memwaddr_r[8]\ : SLE
      port map(D => \memwaddr_r_2[8]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[8]\);
    
    \memwaddr_r[2]\ : SLE
      port map(D => un1_memwaddr_r_cry_2_S_1, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[2]\);
    
    \wptr_bin_sync2[11]\ : SLE
      port map(D => \wptr_bin_sync[11]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[11]_net_1\);
    
    \L1.un4_we_i_7\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \fifo_MEMWADDR[12]\, B => \fifo_MEMWADDR[11]\, 
        C => \fifo_MEMWADDR[6]\, D => \fifo_MEMWADDR[5]\, Y => 
        un4_we_i_7);
    
    \wptr_gray_1[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[1]_net_1\, B => \wptr[2]_net_1\, Y => 
        \wptr_gray_1[1]_net_1\);
    
    underflow_r : SLE
      port map(D => N_5_i, CLK => m2s010_som_sb_0_CCC_71MHz, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => iRX_FIFO_UNDERRUN_0);
    
    \memwaddr_r_2[11]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_11_S_1, D => un4_we_i_9, Y => 
        \memwaddr_r_2[11]_net_1\);
    
    \memraddr_r_2[12]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => 
        un1_memraddr_r_s_12_S_1, D => un4_re_i_9, Y => 
        \memraddr_r_2[12]_net_1\);
    
    \wptr_gray[5]\ : SLE
      port map(D => \wptr_gray_1[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[5]_net_1\);
    
    overflow_r_RNO : CFG3
      generic map(INIT => x"80")

      port map(A => RX_FIFO_TxColDetDis_wr_en, B => 
        \iRX_FIFO_Full_0\, C => iRX_FIFO_wr_en_0_0, Y => N_6_i);
    
    \memraddr_r[7]\ : SLE
      port map(D => \memraddr_r_2[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[7]\);
    
    un1_memraddr_r_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_5\, 
        S => un1_memraddr_r_cry_6_S_1, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_6\);
    
    rptr_s_904 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => rptr_s_904_FCO);
    
    \rptr_bin_sync2[10]\ : SLE
      port map(D => \rptr_bin_sync[10]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[10]_net_1\);
    
    wdiff_bus_s_13 : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \rptr_bin_sync2[13]_net_1\, C
         => \wptr[13]_net_1\, D => GND_net_1, FCI => 
        \wdiff_bus_cry_12\, S => \wdiff_bus[13]\, Y => OPEN, FCO
         => OPEN);
    
    wdiff_bus_cry_10 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[10]_net_1\, B => 
        \rptr_bin_sync2[10]_net_1\, C => GND_net_1, D => 
        GND_net_1, FCI => \wdiff_bus_cry_9\, S => \wdiff_bus[10]\, 
        Y => OPEN, FCO => \wdiff_bus_cry_10\);
    
    \memwaddr_r[11]\ : SLE
      port map(D => \memwaddr_r_2[11]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[11]\);
    
    \wptr_gray[8]\ : SLE
      port map(D => \wptr_gray_1[8]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[8]_net_1\);
    
    \memraddr_r_2[11]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => 
        un1_memraddr_r_cry_11_S_1, D => un4_re_i_9, Y => 
        \memraddr_r_2[11]_net_1\);
    
    un1_memraddr_r_s_12 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[12]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_11\, 
        S => un1_memraddr_r_s_12_S_1, Y => OPEN, FCO => OPEN);
    
    \wptr_gray[7]\ : SLE
      port map(D => \wptr_gray_1[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[7]_net_1\);
    
    \wptr_gray_1[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[5]_net_1\, B => \wptr[6]_net_1\, Y => 
        \wptr_gray_1[5]_net_1\);
    
    \memwaddr_r[5]\ : SLE
      port map(D => \memwaddr_r_2[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[5]\);
    
    \L1.empty_r_3_0_a2\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \rdiff_bus[12]\, B => \rdiff_bus[13]\, C => 
        empty_r_3_0_a2_7, D => empty_r_3_0_a2_11, Y => empty_r_3);
    
    un1_memraddr_r_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_3\, 
        S => un1_memraddr_r_cry_4_S_1, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_4\);
    
    \rptr[8]\ : SLE
      port map(D => \rptr_s[8]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[8]_net_1\);
    
    Rd_corefifo_doubleSync : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_1
      port map(rptr_gray(13) => \rptr_gray[13]_net_1\, 
        rptr_gray(12) => \rptr_gray[12]_net_1\, rptr_gray(11) => 
        \rptr_gray[11]_net_1\, rptr_gray(10) => 
        \rptr_gray[10]_net_1\, rptr_gray(9) => 
        \rptr_gray[9]_net_1\, rptr_gray(8) => 
        \rptr_gray[8]_net_1\, rptr_gray(7) => 
        \rptr_gray[7]_net_1\, rptr_gray(6) => 
        \rptr_gray[6]_net_1\, rptr_gray(5) => 
        \rptr_gray[5]_net_1\, rptr_gray(4) => 
        \rptr_gray[4]_net_1\, rptr_gray(3) => 
        \rptr_gray[3]_net_1\, rptr_gray(2) => 
        \rptr_gray[2]_net_1\, rptr_gray(1) => 
        \rptr_gray[1]_net_1\, rptr_gray(0) => 
        \rptr_gray[0]_net_1\, rptr_gray_sync(12) => 
        \rptr_gray_sync[12]\, rptr_gray_sync(11) => 
        \rptr_gray_sync[11]\, rptr_gray_sync(10) => 
        \rptr_gray_sync[10]\, rptr_gray_sync(9) => 
        \rptr_gray_sync[9]\, rptr_gray_sync(8) => 
        \rptr_gray_sync[8]\, rptr_gray_sync(7) => 
        \rptr_gray_sync[7]\, rptr_gray_sync(6) => 
        \rptr_gray_sync[6]\, rptr_gray_sync(5) => 
        \rptr_gray_sync[5]\, rptr_gray_sync(4) => 
        \rptr_gray_sync[4]\, rptr_gray_sync(3) => 
        \rptr_gray_sync[3]\, rptr_gray_sync(2) => 
        \rptr_gray_sync[2]\, rptr_gray_sync(1) => 
        \rptr_gray_sync[1]\, rptr_gray_sync(0) => 
        \rptr_gray_sync[0]\, rptr_bin_sync_0 => 
        \rptr_bin_sync[13]\, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, irx_fifo_rst_i => irx_fifo_rst_i);
    
    underflow_r_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => iRX_FIFO_rd_en_0, B => \iRX_FIFO_Empty_0\, Y
         => N_5_i);
    
    \rptr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[3]_net_1\, S
         => \rptr_s[4]\, Y => OPEN, FCO => \rptr_cry[4]_net_1\);
    
    wdiff_bus_cry_2 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[2]_net_1\, B => 
        \rptr_bin_sync2[2]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_1\, S => \wdiff_bus[2]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_2\);
    
    \rptr_gray[2]\ : SLE
      port map(D => \rptr_gray_1[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[2]_net_1\);
    
    \wptr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[8]_net_1\, S
         => \wptr_s[9]\, Y => OPEN, FCO => \wptr_cry[9]_net_1\);
    
    \wptr_bin_sync2[3]\ : SLE
      port map(D => \wptr_bin_sync[3]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[3]_net_1\);
    
    \rptr[12]\ : SLE
      port map(D => \rptr_s[12]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rptr[12]_net_1\);
    
    \wptr[2]\ : SLE
      port map(D => \wptr_s[2]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[2]_net_1\);
    
    \rptr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[1]_net_1\, S
         => \rptr_s[2]\, Y => OPEN, FCO => \rptr_cry[2]_net_1\);
    
    rdiff_bus_cry_9 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[9]_net_1\, B => 
        \rptr[9]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_8\, S => \rdiff_bus[9]\, Y => OPEN, FCO
         => \rdiff_bus_cry_9\);
    
    \memwaddr_r[0]\ : SLE
      port map(D => \fifo_MEMWADDR_i[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[0]\);
    
    \wptr_gray[2]\ : SLE
      port map(D => \wptr_gray_1[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[2]_net_1\);
    
    \wptr_cry[12]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[12]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[11]_net_1\, S
         => \wptr_s[12]\, Y => OPEN, FCO => \wptr_cry[12]_net_1\);
    
    \memwaddr_r_2[7]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_7_S_1, D => un4_we_i_9, Y => 
        \memwaddr_r_2[7]_net_1\);
    
    wdiff_bus_cry_4 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[4]_net_1\, B => 
        \rptr_bin_sync2[4]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_3\, S => \wdiff_bus[4]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_4\);
    
    un1_memraddr_r_cry_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_6\, 
        S => un1_memraddr_r_cry_7_S_1, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_7\);
    
    \wptr_s[13]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[13]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[12]_net_1\, S
         => \wptr_s[13]_net_1\, Y => OPEN, FCO => OPEN);
    
    \wptr_gray[11]\ : SLE
      port map(D => \wptr_gray_1[11]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[11]_net_1\);
    
    \wptr_bin_sync2[9]\ : SLE
      port map(D => \wptr_bin_sync[9]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[9]_net_1\);
    
    \rptr_gray_1[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[6]_net_1\, B => \rptr[7]_net_1\, Y => 
        \rptr_gray_1[6]_net_1\);
    
    \wptr_gray_1[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[10]_net_1\, B => \wptr[11]_net_1\, Y
         => \wptr_gray_1[10]_net_1\);
    
    wdiff_bus_cry_6 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[6]_net_1\, B => 
        \rptr_bin_sync2[6]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_5\, S => \wdiff_bus[6]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_6\);
    
    \rptr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[2]_net_1\, S
         => \rptr_s[3]\, Y => OPEN, FCO => \rptr_cry[3]_net_1\);
    
    \memraddr_r[4]\ : SLE
      port map(D => un1_memraddr_r_cry_4_S_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[4]\);
    
    \rptr[13]\ : SLE
      port map(D => \rptr_s[13]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rptr[13]_net_1\);
    
    \wptr_cry[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[10]_net_1\, S
         => \wptr_s[11]\, Y => OPEN, FCO => \wptr_cry[11]_net_1\);
    
    \memwaddr_r_2[8]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_8_S_1, D => un4_we_i_9, Y => 
        \memwaddr_r_2[8]_net_1\);
    
    \memwaddr_r[12]\ : SLE
      port map(D => \memwaddr_r_2[12]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[12]\);
    
    \L1.un4_re_i_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => \fifo_MEMRADDR[1]\, B => \fifo_MEMRADDR[2]\, 
        Y => un4_re_i_0);
    
    \rptr_cry[12]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[12]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[11]_net_1\, S
         => \rptr_s[12]\, Y => OPEN, FCO => \rptr_cry[12]_net_1\);
    
    memre_0_a2 : CFG2
      generic map(INIT => x"2")

      port map(A => iRX_FIFO_rd_en_0, B => \iRX_FIFO_Empty_0\, Y
         => \fifo_MEMRE\);
    
    \memraddr_r[11]\ : SLE
      port map(D => \memraddr_r_2[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[11]\);
    
    rdiff_bus_cry_12 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[12]_net_1\, B => 
        \rptr[12]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_11\, S => \rdiff_bus[12]\, Y => OPEN, FCO
         => \rdiff_bus_cry_12\);
    
    \memraddr_r[5]\ : SLE
      port map(D => \memraddr_r_2[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[5]\);
    
    \rptr_gray[6]\ : SLE
      port map(D => \rptr_gray_1[6]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[6]_net_1\);
    
    \memraddr_r[9]\ : SLE
      port map(D => \memraddr_r_2[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[9]\);
    
    \rptr[0]\ : SLE
      port map(D => \rptr_s[0]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[0]_net_1\);
    
    \wptr[10]\ : SLE
      port map(D => \wptr_s[10]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[10]_net_1\);
    
    \L1.un4_we_i_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => \fifo_MEMWADDR[1]\, B => \fifo_MEMWADDR[2]\, 
        Y => un4_we_i_0);
    
    wdiff_bus_cry_1 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[1]_net_1\, B => 
        \rptr_bin_sync2[1]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_0\, S => \wdiff_bus[1]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_1\);
    
    rdiff_bus_cry_2 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[2]_net_1\, B => 
        \rptr[2]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_1\, S => \rdiff_bus[2]\, Y => OPEN, FCO
         => \rdiff_bus_cry_2\);
    
    \wptr_gray[9]\ : SLE
      port map(D => \wptr_gray_1[9]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[9]_net_1\);
    
    \rptr_gray_1[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[4]_net_1\, B => \rptr[5]_net_1\, Y => 
        \rptr_gray_1[4]_net_1\);
    
    \wptr_gray_1[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[8]_net_1\, B => \wptr[9]_net_1\, Y => 
        \wptr_gray_1[8]_net_1\);
    
    Rd_corefifo_grayToBinConv : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_3
      port map(rptr_bin_sync(13) => \rptr_bin_sync[13]\, 
        rptr_bin_sync(12) => \rptr_bin_sync[12]\, 
        rptr_bin_sync(11) => \rptr_bin_sync[11]\, 
        rptr_bin_sync(10) => \rptr_bin_sync[10]\, 
        rptr_bin_sync(9) => \rptr_bin_sync[9]\, rptr_bin_sync(8)
         => \rptr_bin_sync[8]\, rptr_bin_sync(7) => 
        \rptr_bin_sync[7]\, rptr_bin_sync(6) => nc2, 
        rptr_bin_sync(5) => \rptr_bin_sync[5]\, rptr_bin_sync(4)
         => nc1, rptr_bin_sync(3) => \rptr_bin_sync[3]\, 
        rptr_bin_sync(2) => \rptr_bin_sync[2]\, rptr_bin_sync(1)
         => \rptr_bin_sync[1]\, rptr_bin_sync(0) => 
        \rptr_bin_sync[0]\, rptr_gray_sync(12) => 
        \rptr_gray_sync[12]\, rptr_gray_sync(11) => 
        \rptr_gray_sync[11]\, rptr_gray_sync(10) => 
        \rptr_gray_sync[10]\, rptr_gray_sync(9) => 
        \rptr_gray_sync[9]\, rptr_gray_sync(8) => 
        \rptr_gray_sync[8]\, rptr_gray_sync(7) => 
        \rptr_gray_sync[7]\, rptr_gray_sync(6) => 
        \rptr_gray_sync[6]\, rptr_gray_sync(5) => 
        \rptr_gray_sync[5]\, rptr_gray_sync(4) => 
        \rptr_gray_sync[4]\, rptr_gray_sync(3) => 
        \rptr_gray_sync[3]\, rptr_gray_sync(2) => 
        \rptr_gray_sync[2]\, rptr_gray_sync(1) => 
        \rptr_gray_sync[1]\, rptr_gray_sync(0) => 
        \rptr_gray_sync[0]\, bin_N_6_i => bin_N_6_i, bin_N_4_0_i
         => bin_N_4_0_i);
    
    \rptr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => rptr_s_904_FCO, S => 
        \rptr_s[1]\, Y => OPEN, FCO => \rptr_cry[1]_net_1\);
    
    \rptr_cry[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[10]_net_1\, S
         => \rptr_s[11]\, Y => OPEN, FCO => \rptr_cry[11]_net_1\);
    
    rdiff_bus_cry_3 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[3]_net_1\, B => 
        \rptr[3]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_2\, S => \rdiff_bus[3]\, Y => OPEN, FCO
         => \rdiff_bus_cry_3\);
    
    rdiff_bus_cry_10 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[10]_net_1\, B => 
        \rptr[10]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_9\, S => \rdiff_bus[10]\, Y => OPEN, FCO
         => \rdiff_bus_cry_10\);
    
    un1_memwaddr_r_cry_11 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[11]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_10\, 
        S => un1_memwaddr_r_cry_11_S_1, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_11\);
    
    \memraddr_r[6]\ : SLE
      port map(D => un1_memraddr_r_cry_6_S_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[6]\);
    
    \rptr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[6]_net_1\, S
         => \rptr_s[7]\, Y => OPEN, FCO => \rptr_cry[7]_net_1\);
    
    rdiff_bus_cry_0 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => rdiff_bus, B => \rptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => rdiff_bus_cry_0_Y_2, FCO => \rdiff_bus_cry_0\);
    
    \memraddr_r[2]\ : SLE
      port map(D => un1_memraddr_r_cry_2_S_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[2]\);
    
    \wptr[8]\ : SLE
      port map(D => \wptr_s[8]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[8]_net_1\);
    
    wdiff_bus_cry_3 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[3]_net_1\, B => 
        \rptr_bin_sync2[3]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_2\, S => \wdiff_bus[3]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_3\);
    
    rdiff_bus_s_13 : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \rptr[13]_net_1\, C => 
        \wptr_bin_sync2[13]_net_1\, D => GND_net_1, FCI => 
        \rdiff_bus_cry_12\, S => \rdiff_bus[13]\, Y => OPEN, FCO
         => OPEN);
    
    \memraddr_r[12]\ : SLE
      port map(D => \memraddr_r_2[12]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[12]\);
    
    \wptr_gray_1[11]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[11]_net_1\, B => \wptr[12]_net_1\, Y
         => \wptr_gray_1[11]_net_1\);
    
    \rptr_gray[7]\ : SLE
      port map(D => \rptr_gray_1[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[7]_net_1\);
    
    \wptr_gray[0]\ : SLE
      port map(D => \wptr_gray_1[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[0]_net_1\);
    
    \rptr_gray_1[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[0]_net_1\, B => \rptr[1]_net_1\, Y => 
        \rptr_gray_1[0]_net_1\);
    
    un1_memwaddr_r_cry_10 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_9\, 
        S => un1_memwaddr_r_cry_10_S_1, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_10\);
    
    \rptr_gray_1[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[8]_net_1\, B => \rptr[9]_net_1\, Y => 
        \rptr_gray_1[8]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_1 is

    port( RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          RX_FIFO_DOUT_2            : out   std_logic_vector(8 downto 0);
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_wr_en_0_0        : in    std_logic;
          iRX_FIFO_rd_en_0          : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          RX_FIFO_TxColDetDis_wr_en : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          irx_fifo_rst_i            : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_1;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_1 is 

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_1
    port( fifo_MEMRADDR             : in    std_logic_vector(12 downto 0) := (others => 'U');
          fifo_MEMWADDR             : in    std_logic_vector(12 downto 0) := (others => 'U');
          RDATA_int                 : out   std_logic_vector(8 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          fifo_MEMRE                : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          fifo_MEMWE                : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_1
    port( fifo_MEMRADDR             : out   std_logic_vector(12 downto 0);
          fifo_MEMWADDR             : out   std_logic_vector(12 downto 0);
          iRX_FIFO_wr_en_0_0        : in    std_logic := 'U';
          iRX_FIFO_rd_en_0          : in    std_logic := 'U';
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          RX_FIFO_TxColDetDis_wr_en : in    std_logic := 'U';
          fifo_MEMRE                : out   std_logic;
          fifo_MEMWE                : out   std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          irx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \RDATA_r[0]_net_1\, VCC_net_1, \RDATA_int[0]\, 
        un6_fifo_memre_1, GND_net_1, \RDATA_r[1]_net_1\, 
        \RDATA_int[1]\, \RDATA_r[2]_net_1\, \RDATA_int[2]\, 
        \RDATA_r[3]_net_1\, \RDATA_int[3]\, \RDATA_r[4]_net_1\, 
        \RDATA_int[4]\, \RDATA_r[5]_net_1\, \RDATA_int[5]\, 
        \RDATA_r[6]_net_1\, \RDATA_int[6]\, \RDATA_r[7]_net_1\, 
        \RDATA_int[7]\, \RDATA_r[8]_net_1\, \RDATA_int[8]\, 
        \re_set\, \REN_d1\, un9_fifo_memre_1, fifo_MEMRE, \RE_d1\, 
        \re_pulse_d1\, \re_pulse\, \fifo_MEMRADDR[0]\, 
        \fifo_MEMRADDR[1]\, \fifo_MEMRADDR[2]\, 
        \fifo_MEMRADDR[3]\, \fifo_MEMRADDR[4]\, 
        \fifo_MEMRADDR[5]\, \fifo_MEMRADDR[6]\, 
        \fifo_MEMRADDR[7]\, \fifo_MEMRADDR[8]\, 
        \fifo_MEMRADDR[9]\, \fifo_MEMRADDR[10]\, 
        \fifo_MEMRADDR[11]\, \fifo_MEMRADDR[12]\, 
        \fifo_MEMWADDR[0]\, \fifo_MEMWADDR[1]\, 
        \fifo_MEMWADDR[2]\, \fifo_MEMWADDR[3]\, 
        \fifo_MEMWADDR[4]\, \fifo_MEMWADDR[5]\, 
        \fifo_MEMWADDR[6]\, \fifo_MEMWADDR[7]\, 
        \fifo_MEMWADDR[8]\, \fifo_MEMWADDR[9]\, 
        \fifo_MEMWADDR[10]\, \fifo_MEMWADDR[11]\, 
        \fifo_MEMWADDR[12]\, fifo_MEMWE : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_1
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_1(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_1
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_1(DEF_ARCH);
begin 


    re_pulse : CFG3
      generic map(INIT => x"DC")

      port map(A => fifo_MEMRE, B => \re_set\, C => \REN_d1\, Y
         => \re_pulse\);
    
    \RDATA_r[3]\ : SLE
      port map(D => \RDATA_int[3]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un6_fifo_memre_1, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[3]_net_1\);
    
    \Q[6]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[6]_net_1\, C => 
        \RDATA_int[6]\, D => \RE_d1\, Y => RX_FIFO_DOUT_2(6));
    
    re_pulse_d1 : SLE
      port map(D => \re_pulse\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \re_pulse_d1\);
    
    \RDATA_r[5]\ : SLE
      port map(D => \RDATA_int[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un6_fifo_memre_1, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[5]_net_1\);
    
    un9_fifo_memre : CFG2
      generic map(INIT => x"6")

      port map(A => fifo_MEMRE, B => \REN_d1\, Y => 
        un9_fifo_memre_1);
    
    \RDATA_r[8]\ : SLE
      port map(D => \RDATA_int[8]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un6_fifo_memre_1, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[8]_net_1\);
    
    \Q[2]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[2]_net_1\, C => 
        \RDATA_int[2]\, D => \RE_d1\, Y => RX_FIFO_DOUT_2(2));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \RW1.UI_ram_wrapper_1\ : FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_1
      port map(fifo_MEMRADDR(12) => \fifo_MEMRADDR[12]\, 
        fifo_MEMRADDR(11) => \fifo_MEMRADDR[11]\, 
        fifo_MEMRADDR(10) => \fifo_MEMRADDR[10]\, 
        fifo_MEMRADDR(9) => \fifo_MEMRADDR[9]\, fifo_MEMRADDR(8)
         => \fifo_MEMRADDR[8]\, fifo_MEMRADDR(7) => 
        \fifo_MEMRADDR[7]\, fifo_MEMRADDR(6) => 
        \fifo_MEMRADDR[6]\, fifo_MEMRADDR(5) => 
        \fifo_MEMRADDR[5]\, fifo_MEMRADDR(4) => 
        \fifo_MEMRADDR[4]\, fifo_MEMRADDR(3) => 
        \fifo_MEMRADDR[3]\, fifo_MEMRADDR(2) => 
        \fifo_MEMRADDR[2]\, fifo_MEMRADDR(1) => 
        \fifo_MEMRADDR[1]\, fifo_MEMRADDR(0) => 
        \fifo_MEMRADDR[0]\, fifo_MEMWADDR(12) => 
        \fifo_MEMWADDR[12]\, fifo_MEMWADDR(11) => 
        \fifo_MEMWADDR[11]\, fifo_MEMWADDR(10) => 
        \fifo_MEMWADDR[10]\, fifo_MEMWADDR(9) => 
        \fifo_MEMWADDR[9]\, fifo_MEMWADDR(8) => 
        \fifo_MEMWADDR[8]\, fifo_MEMWADDR(7) => 
        \fifo_MEMWADDR[7]\, fifo_MEMWADDR(6) => 
        \fifo_MEMWADDR[6]\, fifo_MEMWADDR(5) => 
        \fifo_MEMWADDR[5]\, fifo_MEMWADDR(4) => 
        \fifo_MEMWADDR[4]\, fifo_MEMWADDR(3) => 
        \fifo_MEMWADDR[3]\, fifo_MEMWADDR(2) => 
        \fifo_MEMWADDR[2]\, fifo_MEMWADDR(1) => 
        \fifo_MEMWADDR[1]\, fifo_MEMWADDR(0) => 
        \fifo_MEMWADDR[0]\, RDATA_int(8) => \RDATA_int[8]\, 
        RDATA_int(7) => \RDATA_int[7]\, RDATA_int(6) => 
        \RDATA_int[6]\, RDATA_int(5) => \RDATA_int[5]\, 
        RDATA_int(4) => \RDATA_int[4]\, RDATA_int(3) => 
        \RDATA_int[3]\, RDATA_int(2) => \RDATA_int[2]\, 
        RDATA_int(1) => \RDATA_int[1]\, RDATA_int(0) => 
        \RDATA_int[0]\, RX_FIFO_DIN_pipe(8) => 
        RX_FIFO_DIN_pipe(8), RX_FIFO_DIN_pipe(7) => 
        RX_FIFO_DIN_pipe(7), RX_FIFO_DIN_pipe(6) => 
        RX_FIFO_DIN_pipe(6), RX_FIFO_DIN_pipe(5) => 
        RX_FIFO_DIN_pipe(5), RX_FIFO_DIN_pipe(4) => 
        RX_FIFO_DIN_pipe(4), RX_FIFO_DIN_pipe(3) => 
        RX_FIFO_DIN_pipe(3), RX_FIFO_DIN_pipe(2) => 
        RX_FIFO_DIN_pipe(2), RX_FIFO_DIN_pipe(1) => 
        RX_FIFO_DIN_pipe(1), RX_FIFO_DIN_pipe(0) => 
        RX_FIFO_DIN_pipe(0), m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, fifo_MEMRE => fifo_MEMRE, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, fifo_MEMWE
         => fifo_MEMWE);
    
    \RDATA_r[0]\ : SLE
      port map(D => \RDATA_int[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un6_fifo_memre_1, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[0]_net_1\);
    
    \Q[4]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[4]_net_1\, C => 
        \RDATA_int[4]\, D => \RE_d1\, Y => RX_FIFO_DOUT_2(4));
    
    \RDATA_r[2]\ : SLE
      port map(D => \RDATA_int[2]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un6_fifo_memre_1, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[2]_net_1\);
    
    \RDATA_r[6]\ : SLE
      port map(D => \RDATA_int[6]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un6_fifo_memre_1, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[6]_net_1\);
    
    \L31.U_corefifo_async\ : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_1
      port map(fifo_MEMRADDR(12) => \fifo_MEMRADDR[12]\, 
        fifo_MEMRADDR(11) => \fifo_MEMRADDR[11]\, 
        fifo_MEMRADDR(10) => \fifo_MEMRADDR[10]\, 
        fifo_MEMRADDR(9) => \fifo_MEMRADDR[9]\, fifo_MEMRADDR(8)
         => \fifo_MEMRADDR[8]\, fifo_MEMRADDR(7) => 
        \fifo_MEMRADDR[7]\, fifo_MEMRADDR(6) => 
        \fifo_MEMRADDR[6]\, fifo_MEMRADDR(5) => 
        \fifo_MEMRADDR[5]\, fifo_MEMRADDR(4) => 
        \fifo_MEMRADDR[4]\, fifo_MEMRADDR(3) => 
        \fifo_MEMRADDR[3]\, fifo_MEMRADDR(2) => 
        \fifo_MEMRADDR[2]\, fifo_MEMRADDR(1) => 
        \fifo_MEMRADDR[1]\, fifo_MEMRADDR(0) => 
        \fifo_MEMRADDR[0]\, fifo_MEMWADDR(12) => 
        \fifo_MEMWADDR[12]\, fifo_MEMWADDR(11) => 
        \fifo_MEMWADDR[11]\, fifo_MEMWADDR(10) => 
        \fifo_MEMWADDR[10]\, fifo_MEMWADDR(9) => 
        \fifo_MEMWADDR[9]\, fifo_MEMWADDR(8) => 
        \fifo_MEMWADDR[8]\, fifo_MEMWADDR(7) => 
        \fifo_MEMWADDR[7]\, fifo_MEMWADDR(6) => 
        \fifo_MEMWADDR[6]\, fifo_MEMWADDR(5) => 
        \fifo_MEMWADDR[5]\, fifo_MEMWADDR(4) => 
        \fifo_MEMWADDR[4]\, fifo_MEMWADDR(3) => 
        \fifo_MEMWADDR[3]\, fifo_MEMWADDR(2) => 
        \fifo_MEMWADDR[2]\, fifo_MEMWADDR(1) => 
        \fifo_MEMWADDR[1]\, fifo_MEMWADDR(0) => 
        \fifo_MEMWADDR[0]\, iRX_FIFO_wr_en_0_0 => 
        iRX_FIFO_wr_en_0_0, iRX_FIFO_rd_en_0 => iRX_FIFO_rd_en_0, 
        iRX_FIFO_Empty_0 => iRX_FIFO_Empty_0, iRX_FIFO_UNDERRUN_0
         => iRX_FIFO_UNDERRUN_0, iRX_FIFO_OVERFLOW_0 => 
        iRX_FIFO_OVERFLOW_0, iRX_FIFO_Full_0 => iRX_FIFO_Full_0, 
        RX_FIFO_TxColDetDis_wr_en => RX_FIFO_TxColDetDis_wr_en, 
        fifo_MEMRE => fifo_MEMRE, fifo_MEMWE => fifo_MEMWE, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz, 
        irx_fifo_rst_i => irx_fifo_rst_i);
    
    re_set : SLE
      port map(D => \REN_d1\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => un9_fifo_memre_1, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \re_set\);
    
    \Q[3]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[3]_net_1\, C => 
        \RDATA_int[3]\, D => \RE_d1\, Y => RX_FIFO_DOUT_2(3));
    
    \Q[7]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[7]_net_1\, C => 
        \RDATA_int[7]\, D => \RE_d1\, Y => RX_FIFO_DOUT_2(7));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \Q[8]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[8]_net_1\, C => 
        \RDATA_int[8]\, D => \RE_d1\, Y => RX_FIFO_DOUT_2(8));
    
    RE_d1 : SLE
      port map(D => iRX_FIFO_rd_en_0, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RE_d1\);
    
    \RDATA_r[7]\ : SLE
      port map(D => \RDATA_int[7]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un6_fifo_memre_1, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[7]_net_1\);
    
    \RDATA_r[4]\ : SLE
      port map(D => \RDATA_int[4]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un6_fifo_memre_1, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[4]_net_1\);
    
    \Q[1]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[1]_net_1\, C => 
        \RDATA_int[1]\, D => \RE_d1\, Y => RX_FIFO_DOUT_2(1));
    
    \Q[0]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[0]_net_1\, C => 
        \RDATA_int[0]\, D => \RE_d1\, Y => RX_FIFO_DOUT_2(0));
    
    REN_d1 : SLE
      port map(D => fifo_MEMRE, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \REN_d1\);
    
    \Q[5]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[5]_net_1\, C => 
        \RDATA_int[5]\, D => \RE_d1\, Y => RX_FIFO_DOUT_2(5));
    
    un6_fifo_memre : CFG2
      generic map(INIT => x"4")

      port map(A => fifo_MEMRE, B => \REN_d1\, Y => 
        un6_fifo_memre_1);
    
    \RDATA_r[1]\ : SLE
      port map(D => \RDATA_int[1]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un6_fifo_memre_1, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[1]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_1 is

    port( RX_FIFO_DOUT_2            : out   std_logic_vector(8 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          iRX_FIFO_rd_en_0          : in    std_logic;
          iRX_FIFO_wr_en_0_0        : in    std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          irx_fifo_rst_i            : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          RX_FIFO_TxColDetDis_wr_en : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic
        );

end FIFO_8Kx9_1;

architecture DEF_ARCH of FIFO_8Kx9_1 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_1
    port( RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          RX_FIFO_DOUT_2            : out   std_logic_vector(8 downto 0);
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_wr_en_0_0        : in    std_logic := 'U';
          iRX_FIFO_rd_en_0          : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          RX_FIFO_TxColDetDis_wr_en : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          irx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_1
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_1(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    FIFO_8Kx9_0 : FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_1
      port map(RX_FIFO_DIN_pipe(8) => RX_FIFO_DIN_pipe(8), 
        RX_FIFO_DIN_pipe(7) => RX_FIFO_DIN_pipe(7), 
        RX_FIFO_DIN_pipe(6) => RX_FIFO_DIN_pipe(6), 
        RX_FIFO_DIN_pipe(5) => RX_FIFO_DIN_pipe(5), 
        RX_FIFO_DIN_pipe(4) => RX_FIFO_DIN_pipe(4), 
        RX_FIFO_DIN_pipe(3) => RX_FIFO_DIN_pipe(3), 
        RX_FIFO_DIN_pipe(2) => RX_FIFO_DIN_pipe(2), 
        RX_FIFO_DIN_pipe(1) => RX_FIFO_DIN_pipe(1), 
        RX_FIFO_DIN_pipe(0) => RX_FIFO_DIN_pipe(0), 
        RX_FIFO_DOUT_2(8) => RX_FIFO_DOUT_2(8), RX_FIFO_DOUT_2(7)
         => RX_FIFO_DOUT_2(7), RX_FIFO_DOUT_2(6) => 
        RX_FIFO_DOUT_2(6), RX_FIFO_DOUT_2(5) => RX_FIFO_DOUT_2(5), 
        RX_FIFO_DOUT_2(4) => RX_FIFO_DOUT_2(4), RX_FIFO_DOUT_2(3)
         => RX_FIFO_DOUT_2(3), RX_FIFO_DOUT_2(2) => 
        RX_FIFO_DOUT_2(2), RX_FIFO_DOUT_2(1) => RX_FIFO_DOUT_2(1), 
        RX_FIFO_DOUT_2(0) => RX_FIFO_DOUT_2(0), iRX_FIFO_Full_0
         => iRX_FIFO_Full_0, iRX_FIFO_OVERFLOW_0 => 
        iRX_FIFO_OVERFLOW_0, iRX_FIFO_UNDERRUN_0 => 
        iRX_FIFO_UNDERRUN_0, iRX_FIFO_Empty_0 => iRX_FIFO_Empty_0, 
        iRX_FIFO_wr_en_0_0 => iRX_FIFO_wr_en_0_0, 
        iRX_FIFO_rd_en_0 => iRX_FIFO_rd_en_0, CommsFPGA_CCC_0_GL0
         => CommsFPGA_CCC_0_GL0, RX_FIFO_TxColDetDis_wr_en => 
        RX_FIFO_TxColDetDis_wr_en, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, irx_fifo_rst_i => 
        irx_fifo_rst_i);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_2 is

    port( RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          RDATA_int                 : out   std_logic_vector(8 downto 0);
          fifo_MEMWADDR             : in    std_logic_vector(12 downto 0);
          fifo_MEMRADDR             : in    std_logic_vector(12 downto 0);
          fifo_MEMWE                : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          fifo_MEMRE                : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_2;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_2 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component RAM1K18
    generic (MEMORYFILE:string := "");

    port( A_DOUT        : out   std_logic_vector(17 downto 0);
          B_DOUT        : out   std_logic_vector(17 downto 0);
          BUSY          : out   std_logic;
          A_CLK         : in    std_logic := 'U';
          A_DOUT_CLK    : in    std_logic := 'U';
          A_ARST_N      : in    std_logic := 'U';
          A_DOUT_EN     : in    std_logic := 'U';
          A_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_DOUT_ARST_N : in    std_logic := 'U';
          A_DOUT_SRST_N : in    std_logic := 'U';
          A_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          A_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          A_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          B_CLK         : in    std_logic := 'U';
          B_DOUT_CLK    : in    std_logic := 'U';
          B_ARST_N      : in    std_logic := 'U';
          B_DOUT_EN     : in    std_logic := 'U';
          B_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_DOUT_ARST_N : in    std_logic := 'U';
          B_DOUT_SRST_N : in    std_logic := 'U';
          B_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          B_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          B_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          A_EN          : in    std_logic := 'U';
          A_DOUT_LAT    : in    std_logic := 'U';
          A_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_WMODE       : in    std_logic := 'U';
          B_EN          : in    std_logic := 'U';
          B_DOUT_LAT    : in    std_logic := 'U';
          B_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_WMODE       : in    std_logic := 'U';
          SII_LOCK      : in    std_logic := 'U'
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;
    signal nc151, nc23, nc58, nc116, nc74, nc133, nc167, nc84, 
        nc39, nc72, nc82, nc145, nc160, nc57, nc156, nc125, nc73, 
        nc107, nc66, nc83, nc9, nc171, nc54, nc135, nc41, nc100, 
        nc52, nc29, nc118, nc60, nc141, nc45, nc53, nc121, nc158, 
        nc162, nc11, nc131, nc96, nc79, nc146, nc89, nc119, nc48, 
        nc126, nc15, nc102, nc3, nc47, nc90, nc159, nc136, nc59, 
        nc18, nc44, nc117, nc164, nc148, nc42, nc17, nc2, nc110, 
        nc128, nc43, nc157, nc36, nc61, nc104, nc138, nc14, nc150, 
        nc149, nc12, nc30, nc65, nc7, nc129, nc8, nc13, nc26, 
        nc139, nc163, nc112, nc68, nc49, nc170, nc91, nc5, nc20, 
        nc147, nc67, nc152, nc127, nc103, nc76, nc140, nc86, nc95, 
        nc120, nc165, nc137, nc64, nc19, nc70, nc62, nc80, nc130, 
        nc98, nc114, nc56, nc105, nc63, nc97, nc161, nc31, nc154, 
        nc50, nc142, nc94, nc122, nc35, nc4, nc92, nc101, nc166, 
        nc132, nc21, nc93, nc69, nc38, nc113, nc106, nc25, nc1, 
        nc37, nc144, nc153, nc46, nc71, nc124, nc81, nc168, nc34, 
        nc28, nc115, nc134, nc32, nc40, nc99, nc75, nc85, nc27, 
        nc108, nc16, nc155, nc51, nc33, nc169, nc78, nc24, nc88, 
        nc111, nc55, nc10, nc22, nc143, nc77, nc6, nc109, nc87, 
        nc123 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C2 : RAM1K18
      port map(A_DOUT(17) => nc151, A_DOUT(16) => nc23, 
        A_DOUT(15) => nc58, A_DOUT(14) => nc116, A_DOUT(13) => 
        nc74, A_DOUT(12) => nc133, A_DOUT(11) => nc167, 
        A_DOUT(10) => nc84, A_DOUT(9) => nc39, A_DOUT(8) => nc72, 
        A_DOUT(7) => nc82, A_DOUT(6) => nc145, A_DOUT(5) => nc160, 
        A_DOUT(4) => nc57, A_DOUT(3) => nc156, A_DOUT(2) => nc125, 
        A_DOUT(1) => RDATA_int(5), A_DOUT(0) => RDATA_int(4), 
        B_DOUT(17) => nc73, B_DOUT(16) => nc107, B_DOUT(15) => 
        nc66, B_DOUT(14) => nc83, B_DOUT(13) => nc9, B_DOUT(12)
         => nc171, B_DOUT(11) => nc54, B_DOUT(10) => nc135, 
        B_DOUT(9) => nc41, B_DOUT(8) => nc100, B_DOUT(7) => nc52, 
        B_DOUT(6) => nc29, B_DOUT(5) => nc118, B_DOUT(4) => nc60, 
        B_DOUT(3) => nc141, B_DOUT(2) => nc45, B_DOUT(1) => nc53, 
        B_DOUT(0) => nc121, BUSY => OPEN, A_CLK => 
        m2s010_som_sb_0_CCC_71MHz, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => fifo_MEMRE, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => fifo_MEMRADDR(12), A_ADDR(12) => fifo_MEMRADDR(11), 
        A_ADDR(11) => fifo_MEMRADDR(10), A_ADDR(10) => 
        fifo_MEMRADDR(9), A_ADDR(9) => fifo_MEMRADDR(8), 
        A_ADDR(8) => fifo_MEMRADDR(7), A_ADDR(7) => 
        fifo_MEMRADDR(6), A_ADDR(6) => fifo_MEMRADDR(5), 
        A_ADDR(5) => fifo_MEMRADDR(4), A_ADDR(4) => 
        fifo_MEMRADDR(3), A_ADDR(3) => fifo_MEMRADDR(2), 
        A_ADDR(2) => fifo_MEMRADDR(1), A_ADDR(1) => 
        fifo_MEMRADDR(0), A_ADDR(0) => GND_net_1, A_WEN(1) => 
        GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => GND_net_1, B_DIN(2) => GND_net_1, B_DIN(1)
         => RX_FIFO_DIN_pipe(5), B_DIN(0) => RX_FIFO_DIN_pipe(4), 
        B_ADDR(13) => fifo_MEMWADDR(12), B_ADDR(12) => 
        fifo_MEMWADDR(11), B_ADDR(11) => fifo_MEMWADDR(10), 
        B_ADDR(10) => fifo_MEMWADDR(9), B_ADDR(9) => 
        fifo_MEMWADDR(8), B_ADDR(8) => fifo_MEMWADDR(7), 
        B_ADDR(7) => fifo_MEMWADDR(6), B_ADDR(6) => 
        fifo_MEMWADDR(5), B_ADDR(5) => fifo_MEMWADDR(4), 
        B_ADDR(4) => fifo_MEMWADDR(3), B_ADDR(3) => 
        fifo_MEMWADDR(2), B_ADDR(2) => fifo_MEMWADDR(1), 
        B_ADDR(1) => fifo_MEMWADDR(0), B_ADDR(0) => GND_net_1, 
        B_WEN(1) => GND_net_1, B_WEN(0) => VCC_net_1, A_EN => 
        VCC_net_1, A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => 
        GND_net_1, A_WIDTH(1) => GND_net_1, A_WIDTH(0) => 
        VCC_net_1, A_WMODE => GND_net_1, B_EN => VCC_net_1, 
        B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => GND_net_1, 
        B_WIDTH(1) => GND_net_1, B_WIDTH(0) => VCC_net_1, B_WMODE
         => GND_net_1, SII_LOCK => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C1 : RAM1K18
      port map(A_DOUT(17) => nc158, A_DOUT(16) => nc162, 
        A_DOUT(15) => nc11, A_DOUT(14) => nc131, A_DOUT(13) => 
        nc96, A_DOUT(12) => nc79, A_DOUT(11) => nc146, A_DOUT(10)
         => nc89, A_DOUT(9) => nc119, A_DOUT(8) => nc48, 
        A_DOUT(7) => nc126, A_DOUT(6) => nc15, A_DOUT(5) => nc102, 
        A_DOUT(4) => nc3, A_DOUT(3) => nc47, A_DOUT(2) => nc90, 
        A_DOUT(1) => RDATA_int(3), A_DOUT(0) => RDATA_int(2), 
        B_DOUT(17) => nc159, B_DOUT(16) => nc136, B_DOUT(15) => 
        nc59, B_DOUT(14) => nc18, B_DOUT(13) => nc44, B_DOUT(12)
         => nc117, B_DOUT(11) => nc164, B_DOUT(10) => nc148, 
        B_DOUT(9) => nc42, B_DOUT(8) => nc17, B_DOUT(7) => nc2, 
        B_DOUT(6) => nc110, B_DOUT(5) => nc128, B_DOUT(4) => nc43, 
        B_DOUT(3) => nc157, B_DOUT(2) => nc36, B_DOUT(1) => nc61, 
        B_DOUT(0) => nc104, BUSY => OPEN, A_CLK => 
        m2s010_som_sb_0_CCC_71MHz, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => fifo_MEMRE, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => fifo_MEMRADDR(12), A_ADDR(12) => fifo_MEMRADDR(11), 
        A_ADDR(11) => fifo_MEMRADDR(10), A_ADDR(10) => 
        fifo_MEMRADDR(9), A_ADDR(9) => fifo_MEMRADDR(8), 
        A_ADDR(8) => fifo_MEMRADDR(7), A_ADDR(7) => 
        fifo_MEMRADDR(6), A_ADDR(6) => fifo_MEMRADDR(5), 
        A_ADDR(5) => fifo_MEMRADDR(4), A_ADDR(4) => 
        fifo_MEMRADDR(3), A_ADDR(3) => fifo_MEMRADDR(2), 
        A_ADDR(2) => fifo_MEMRADDR(1), A_ADDR(1) => 
        fifo_MEMRADDR(0), A_ADDR(0) => GND_net_1, A_WEN(1) => 
        GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => GND_net_1, B_DIN(2) => GND_net_1, B_DIN(1)
         => RX_FIFO_DIN_pipe(3), B_DIN(0) => RX_FIFO_DIN_pipe(2), 
        B_ADDR(13) => fifo_MEMWADDR(12), B_ADDR(12) => 
        fifo_MEMWADDR(11), B_ADDR(11) => fifo_MEMWADDR(10), 
        B_ADDR(10) => fifo_MEMWADDR(9), B_ADDR(9) => 
        fifo_MEMWADDR(8), B_ADDR(8) => fifo_MEMWADDR(7), 
        B_ADDR(7) => fifo_MEMWADDR(6), B_ADDR(6) => 
        fifo_MEMWADDR(5), B_ADDR(5) => fifo_MEMWADDR(4), 
        B_ADDR(4) => fifo_MEMWADDR(3), B_ADDR(3) => 
        fifo_MEMWADDR(2), B_ADDR(2) => fifo_MEMWADDR(1), 
        B_ADDR(1) => fifo_MEMWADDR(0), B_ADDR(0) => GND_net_1, 
        B_WEN(1) => GND_net_1, B_WEN(0) => VCC_net_1, A_EN => 
        VCC_net_1, A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => 
        GND_net_1, A_WIDTH(1) => GND_net_1, A_WIDTH(0) => 
        VCC_net_1, A_WMODE => GND_net_1, B_EN => VCC_net_1, 
        B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => GND_net_1, 
        B_WIDTH(1) => GND_net_1, B_WIDTH(0) => VCC_net_1, B_WMODE
         => GND_net_1, SII_LOCK => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C4 : RAM1K18
      port map(A_DOUT(17) => nc138, A_DOUT(16) => nc14, 
        A_DOUT(15) => nc150, A_DOUT(14) => nc149, A_DOUT(13) => 
        nc12, A_DOUT(12) => nc30, A_DOUT(11) => nc65, A_DOUT(10)
         => nc7, A_DOUT(9) => nc129, A_DOUT(8) => nc8, A_DOUT(7)
         => nc13, A_DOUT(6) => nc26, A_DOUT(5) => nc139, 
        A_DOUT(4) => nc163, A_DOUT(3) => nc112, A_DOUT(2) => nc68, 
        A_DOUT(1) => nc49, A_DOUT(0) => RDATA_int(8), B_DOUT(17)
         => nc170, B_DOUT(16) => nc91, B_DOUT(15) => nc5, 
        B_DOUT(14) => nc20, B_DOUT(13) => nc147, B_DOUT(12) => 
        nc67, B_DOUT(11) => nc152, B_DOUT(10) => nc127, B_DOUT(9)
         => nc103, B_DOUT(8) => nc76, B_DOUT(7) => nc140, 
        B_DOUT(6) => nc86, B_DOUT(5) => nc95, B_DOUT(4) => nc120, 
        B_DOUT(3) => nc165, B_DOUT(2) => nc137, B_DOUT(1) => nc64, 
        B_DOUT(0) => nc19, BUSY => OPEN, A_CLK => 
        m2s010_som_sb_0_CCC_71MHz, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => fifo_MEMRE, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => fifo_MEMRADDR(12), A_ADDR(12) => fifo_MEMRADDR(11), 
        A_ADDR(11) => fifo_MEMRADDR(10), A_ADDR(10) => 
        fifo_MEMRADDR(9), A_ADDR(9) => fifo_MEMRADDR(8), 
        A_ADDR(8) => fifo_MEMRADDR(7), A_ADDR(7) => 
        fifo_MEMRADDR(6), A_ADDR(6) => fifo_MEMRADDR(5), 
        A_ADDR(5) => fifo_MEMRADDR(4), A_ADDR(4) => 
        fifo_MEMRADDR(3), A_ADDR(3) => fifo_MEMRADDR(2), 
        A_ADDR(2) => fifo_MEMRADDR(1), A_ADDR(1) => 
        fifo_MEMRADDR(0), A_ADDR(0) => GND_net_1, A_WEN(1) => 
        GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => GND_net_1, B_DIN(2) => GND_net_1, B_DIN(1)
         => GND_net_1, B_DIN(0) => RX_FIFO_DIN_pipe(8), 
        B_ADDR(13) => fifo_MEMWADDR(12), B_ADDR(12) => 
        fifo_MEMWADDR(11), B_ADDR(11) => fifo_MEMWADDR(10), 
        B_ADDR(10) => fifo_MEMWADDR(9), B_ADDR(9) => 
        fifo_MEMWADDR(8), B_ADDR(8) => fifo_MEMWADDR(7), 
        B_ADDR(7) => fifo_MEMWADDR(6), B_ADDR(6) => 
        fifo_MEMWADDR(5), B_ADDR(5) => fifo_MEMWADDR(4), 
        B_ADDR(4) => fifo_MEMWADDR(3), B_ADDR(3) => 
        fifo_MEMWADDR(2), B_ADDR(2) => fifo_MEMWADDR(1), 
        B_ADDR(1) => fifo_MEMWADDR(0), B_ADDR(0) => GND_net_1, 
        B_WEN(1) => GND_net_1, B_WEN(0) => VCC_net_1, A_EN => 
        VCC_net_1, A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => 
        GND_net_1, A_WIDTH(1) => GND_net_1, A_WIDTH(0) => 
        VCC_net_1, A_WMODE => GND_net_1, B_EN => VCC_net_1, 
        B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => GND_net_1, 
        B_WIDTH(1) => GND_net_1, B_WIDTH(0) => VCC_net_1, B_WMODE
         => GND_net_1, SII_LOCK => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C3 : RAM1K18
      port map(A_DOUT(17) => nc70, A_DOUT(16) => nc62, A_DOUT(15)
         => nc80, A_DOUT(14) => nc130, A_DOUT(13) => nc98, 
        A_DOUT(12) => nc114, A_DOUT(11) => nc56, A_DOUT(10) => 
        nc105, A_DOUT(9) => nc63, A_DOUT(8) => nc97, A_DOUT(7)
         => nc161, A_DOUT(6) => nc31, A_DOUT(5) => nc154, 
        A_DOUT(4) => nc50, A_DOUT(3) => nc142, A_DOUT(2) => nc94, 
        A_DOUT(1) => RDATA_int(7), A_DOUT(0) => RDATA_int(6), 
        B_DOUT(17) => nc122, B_DOUT(16) => nc35, B_DOUT(15) => 
        nc4, B_DOUT(14) => nc92, B_DOUT(13) => nc101, B_DOUT(12)
         => nc166, B_DOUT(11) => nc132, B_DOUT(10) => nc21, 
        B_DOUT(9) => nc93, B_DOUT(8) => nc69, B_DOUT(7) => nc38, 
        B_DOUT(6) => nc113, B_DOUT(5) => nc106, B_DOUT(4) => nc25, 
        B_DOUT(3) => nc1, B_DOUT(2) => nc37, B_DOUT(1) => nc144, 
        B_DOUT(0) => nc153, BUSY => OPEN, A_CLK => 
        m2s010_som_sb_0_CCC_71MHz, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => fifo_MEMRE, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => fifo_MEMRADDR(12), A_ADDR(12) => fifo_MEMRADDR(11), 
        A_ADDR(11) => fifo_MEMRADDR(10), A_ADDR(10) => 
        fifo_MEMRADDR(9), A_ADDR(9) => fifo_MEMRADDR(8), 
        A_ADDR(8) => fifo_MEMRADDR(7), A_ADDR(7) => 
        fifo_MEMRADDR(6), A_ADDR(6) => fifo_MEMRADDR(5), 
        A_ADDR(5) => fifo_MEMRADDR(4), A_ADDR(4) => 
        fifo_MEMRADDR(3), A_ADDR(3) => fifo_MEMRADDR(2), 
        A_ADDR(2) => fifo_MEMRADDR(1), A_ADDR(1) => 
        fifo_MEMRADDR(0), A_ADDR(0) => GND_net_1, A_WEN(1) => 
        GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => GND_net_1, B_DIN(2) => GND_net_1, B_DIN(1)
         => RX_FIFO_DIN_pipe(7), B_DIN(0) => RX_FIFO_DIN_pipe(6), 
        B_ADDR(13) => fifo_MEMWADDR(12), B_ADDR(12) => 
        fifo_MEMWADDR(11), B_ADDR(11) => fifo_MEMWADDR(10), 
        B_ADDR(10) => fifo_MEMWADDR(9), B_ADDR(9) => 
        fifo_MEMWADDR(8), B_ADDR(8) => fifo_MEMWADDR(7), 
        B_ADDR(7) => fifo_MEMWADDR(6), B_ADDR(6) => 
        fifo_MEMWADDR(5), B_ADDR(5) => fifo_MEMWADDR(4), 
        B_ADDR(4) => fifo_MEMWADDR(3), B_ADDR(3) => 
        fifo_MEMWADDR(2), B_ADDR(2) => fifo_MEMWADDR(1), 
        B_ADDR(1) => fifo_MEMWADDR(0), B_ADDR(0) => GND_net_1, 
        B_WEN(1) => GND_net_1, B_WEN(0) => VCC_net_1, A_EN => 
        VCC_net_1, A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => 
        GND_net_1, A_WIDTH(1) => GND_net_1, A_WIDTH(0) => 
        VCC_net_1, A_WMODE => GND_net_1, B_EN => VCC_net_1, 
        B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => GND_net_1, 
        B_WIDTH(1) => GND_net_1, B_WIDTH(0) => VCC_net_1, B_WMODE
         => GND_net_1, SII_LOCK => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C0 : RAM1K18
      port map(A_DOUT(17) => nc46, A_DOUT(16) => nc71, A_DOUT(15)
         => nc124, A_DOUT(14) => nc81, A_DOUT(13) => nc168, 
        A_DOUT(12) => nc34, A_DOUT(11) => nc28, A_DOUT(10) => 
        nc115, A_DOUT(9) => nc134, A_DOUT(8) => nc32, A_DOUT(7)
         => nc40, A_DOUT(6) => nc99, A_DOUT(5) => nc75, A_DOUT(4)
         => nc85, A_DOUT(3) => nc27, A_DOUT(2) => nc108, 
        A_DOUT(1) => RDATA_int(1), A_DOUT(0) => RDATA_int(0), 
        B_DOUT(17) => nc16, B_DOUT(16) => nc155, B_DOUT(15) => 
        nc51, B_DOUT(14) => nc33, B_DOUT(13) => nc169, B_DOUT(12)
         => nc78, B_DOUT(11) => nc24, B_DOUT(10) => nc88, 
        B_DOUT(9) => nc111, B_DOUT(8) => nc55, B_DOUT(7) => nc10, 
        B_DOUT(6) => nc22, B_DOUT(5) => nc143, B_DOUT(4) => nc77, 
        B_DOUT(3) => nc6, B_DOUT(2) => nc109, B_DOUT(1) => nc87, 
        B_DOUT(0) => nc123, BUSY => OPEN, A_CLK => 
        m2s010_som_sb_0_CCC_71MHz, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => fifo_MEMRE, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => fifo_MEMRADDR(12), A_ADDR(12) => fifo_MEMRADDR(11), 
        A_ADDR(11) => fifo_MEMRADDR(10), A_ADDR(10) => 
        fifo_MEMRADDR(9), A_ADDR(9) => fifo_MEMRADDR(8), 
        A_ADDR(8) => fifo_MEMRADDR(7), A_ADDR(7) => 
        fifo_MEMRADDR(6), A_ADDR(6) => fifo_MEMRADDR(5), 
        A_ADDR(5) => fifo_MEMRADDR(4), A_ADDR(4) => 
        fifo_MEMRADDR(3), A_ADDR(3) => fifo_MEMRADDR(2), 
        A_ADDR(2) => fifo_MEMRADDR(1), A_ADDR(1) => 
        fifo_MEMRADDR(0), A_ADDR(0) => GND_net_1, A_WEN(1) => 
        GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => GND_net_1, B_DIN(2) => GND_net_1, B_DIN(1)
         => RX_FIFO_DIN_pipe(1), B_DIN(0) => RX_FIFO_DIN_pipe(0), 
        B_ADDR(13) => fifo_MEMWADDR(12), B_ADDR(12) => 
        fifo_MEMWADDR(11), B_ADDR(11) => fifo_MEMWADDR(10), 
        B_ADDR(10) => fifo_MEMWADDR(9), B_ADDR(9) => 
        fifo_MEMWADDR(8), B_ADDR(8) => fifo_MEMWADDR(7), 
        B_ADDR(7) => fifo_MEMWADDR(6), B_ADDR(6) => 
        fifo_MEMWADDR(5), B_ADDR(5) => fifo_MEMWADDR(4), 
        B_ADDR(4) => fifo_MEMWADDR(3), B_ADDR(3) => 
        fifo_MEMWADDR(2), B_ADDR(2) => fifo_MEMWADDR(1), 
        B_ADDR(1) => fifo_MEMWADDR(0), B_ADDR(0) => GND_net_1, 
        B_WEN(1) => GND_net_1, B_WEN(0) => VCC_net_1, A_EN => 
        VCC_net_1, A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => 
        GND_net_1, A_WIDTH(1) => GND_net_1, A_WIDTH(0) => 
        VCC_net_1, A_WMODE => GND_net_1, B_EN => VCC_net_1, 
        B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => GND_net_1, 
        B_WIDTH(1) => GND_net_1, B_WIDTH(0) => VCC_net_1, B_WMODE
         => GND_net_1, SII_LOCK => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_2 is

    port( fifo_MEMRADDR             : in    std_logic_vector(12 downto 0);
          fifo_MEMWADDR             : in    std_logic_vector(12 downto 0);
          RDATA_int                 : out   std_logic_vector(8 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          fifo_MEMRE                : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          fifo_MEMWE                : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_2;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_2 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_2
    port( RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          RDATA_int                 : out   std_logic_vector(8 downto 0);
          fifo_MEMWADDR             : in    std_logic_vector(12 downto 0) := (others => 'U');
          fifo_MEMRADDR             : in    std_logic_vector(12 downto 0) := (others => 'U');
          fifo_MEMWE                : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          fifo_MEMRE                : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_2
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_2(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    L1_asyncnonpipe : FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_2
      port map(RX_FIFO_DIN_pipe(8) => RX_FIFO_DIN_pipe(8), 
        RX_FIFO_DIN_pipe(7) => RX_FIFO_DIN_pipe(7), 
        RX_FIFO_DIN_pipe(6) => RX_FIFO_DIN_pipe(6), 
        RX_FIFO_DIN_pipe(5) => RX_FIFO_DIN_pipe(5), 
        RX_FIFO_DIN_pipe(4) => RX_FIFO_DIN_pipe(4), 
        RX_FIFO_DIN_pipe(3) => RX_FIFO_DIN_pipe(3), 
        RX_FIFO_DIN_pipe(2) => RX_FIFO_DIN_pipe(2), 
        RX_FIFO_DIN_pipe(1) => RX_FIFO_DIN_pipe(1), 
        RX_FIFO_DIN_pipe(0) => RX_FIFO_DIN_pipe(0), RDATA_int(8)
         => RDATA_int(8), RDATA_int(7) => RDATA_int(7), 
        RDATA_int(6) => RDATA_int(6), RDATA_int(5) => 
        RDATA_int(5), RDATA_int(4) => RDATA_int(4), RDATA_int(3)
         => RDATA_int(3), RDATA_int(2) => RDATA_int(2), 
        RDATA_int(1) => RDATA_int(1), RDATA_int(0) => 
        RDATA_int(0), fifo_MEMWADDR(12) => fifo_MEMWADDR(12), 
        fifo_MEMWADDR(11) => fifo_MEMWADDR(11), fifo_MEMWADDR(10)
         => fifo_MEMWADDR(10), fifo_MEMWADDR(9) => 
        fifo_MEMWADDR(9), fifo_MEMWADDR(8) => fifo_MEMWADDR(8), 
        fifo_MEMWADDR(7) => fifo_MEMWADDR(7), fifo_MEMWADDR(6)
         => fifo_MEMWADDR(6), fifo_MEMWADDR(5) => 
        fifo_MEMWADDR(5), fifo_MEMWADDR(4) => fifo_MEMWADDR(4), 
        fifo_MEMWADDR(3) => fifo_MEMWADDR(3), fifo_MEMWADDR(2)
         => fifo_MEMWADDR(2), fifo_MEMWADDR(1) => 
        fifo_MEMWADDR(1), fifo_MEMWADDR(0) => fifo_MEMWADDR(0), 
        fifo_MEMRADDR(12) => fifo_MEMRADDR(12), fifo_MEMRADDR(11)
         => fifo_MEMRADDR(11), fifo_MEMRADDR(10) => 
        fifo_MEMRADDR(10), fifo_MEMRADDR(9) => fifo_MEMRADDR(9), 
        fifo_MEMRADDR(8) => fifo_MEMRADDR(8), fifo_MEMRADDR(7)
         => fifo_MEMRADDR(7), fifo_MEMRADDR(6) => 
        fifo_MEMRADDR(6), fifo_MEMRADDR(5) => fifo_MEMRADDR(5), 
        fifo_MEMRADDR(4) => fifo_MEMRADDR(4), fifo_MEMRADDR(3)
         => fifo_MEMRADDR(3), fifo_MEMRADDR(2) => 
        fifo_MEMRADDR(2), fifo_MEMRADDR(1) => fifo_MEMRADDR(1), 
        fifo_MEMRADDR(0) => fifo_MEMRADDR(0), fifo_MEMWE => 
        fifo_MEMWE, CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, 
        fifo_MEMRE => fifo_MEMRE, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_6 is

    port( wptr_bin_sync  : inout std_logic_vector(13 downto 0) := (others => 'Z');
          wptr_gray_sync : in    std_logic_vector(12 downto 0)
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_6;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_6 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    \bin_out_xhdl1_0_a2[1]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(3), B => wptr_gray_sync(1), C
         => wptr_bin_sync(4), D => wptr_gray_sync(2), Y => 
        wptr_bin_sync(1));
    
    \bin_out_xhdl1_0_a2[10]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(12), B => wptr_gray_sync(11), 
        C => wptr_gray_sync(10), D => wptr_bin_sync(13), Y => 
        wptr_bin_sync(10));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \bin_out_xhdl1_0_a2[5]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(7), B => wptr_gray_sync(6), C
         => wptr_gray_sync(5), D => wptr_bin_sync(8), Y => 
        wptr_bin_sync(5));
    
    \bin_out_xhdl1_0_a2[2]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(4), B => wptr_gray_sync(3), C
         => wptr_gray_sync(2), D => wptr_bin_sync(5), Y => 
        wptr_bin_sync(2));
    
    \bin_out_xhdl1_0_a2[0]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(2), B => wptr_bin_sync(3), C
         => wptr_gray_sync(0), D => wptr_gray_sync(1), Y => 
        wptr_bin_sync(0));
    
    \bin_out_xhdl1_0_a2[9]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(11), B => wptr_gray_sync(10), 
        C => wptr_gray_sync(9), D => wptr_bin_sync(12), Y => 
        wptr_bin_sync(9));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \bin_out_xhdl1_i_o2[12]\ : CFG2
      generic map(INIT => x"6")

      port map(A => wptr_bin_sync(13), B => wptr_gray_sync(12), Y
         => wptr_bin_sync(12));
    
    \bin_out_xhdl1_0_a2[6]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(8), B => wptr_gray_sync(7), C
         => wptr_gray_sync(6), D => wptr_bin_sync(9), Y => 
        wptr_bin_sync(6));
    
    \bin_out_xhdl1_0_a2[4]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(6), B => wptr_gray_sync(5), C
         => wptr_gray_sync(4), D => wptr_bin_sync(7), Y => 
        wptr_bin_sync(4));
    
    \bin_out_xhdl1_i_o2[11]\ : CFG3
      generic map(INIT => x"96")

      port map(A => wptr_gray_sync(12), B => wptr_gray_sync(11), 
        C => wptr_bin_sync(13), Y => wptr_bin_sync(11));
    
    \bin_out_xhdl1_0_a2[8]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(10), B => wptr_gray_sync(9), C
         => wptr_gray_sync(8), D => wptr_bin_sync(11), Y => 
        wptr_bin_sync(8));
    
    \bin_out_xhdl1_0_a2[7]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(9), B => wptr_gray_sync(8), C
         => wptr_gray_sync(7), D => wptr_bin_sync(10), Y => 
        wptr_bin_sync(7));
    
    \bin_out_xhdl1_0_a2[3]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(5), B => wptr_gray_sync(4), C
         => wptr_gray_sync(3), D => wptr_bin_sync(6), Y => 
        wptr_bin_sync(3));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_3 is

    port( wptr_gray                 : in    std_logic_vector(13 downto 0);
          wptr_gray_sync            : out   std_logic_vector(12 downto 0);
          wptr_bin_sync_0           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          irx_fifo_rst_i            : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_3;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_3 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \sync_int[11]_net_1\, GND_net_1, 
        \sync_int[12]_net_1\, \sync_int[13]_net_1\, 
        \sync_int[10]_net_1\, \sync_int[0]_net_1\, 
        \sync_int[1]_net_1\, \sync_int[2]_net_1\, 
        \sync_int[3]_net_1\, \sync_int[4]_net_1\, 
        \sync_int[5]_net_1\, \sync_int[6]_net_1\, 
        \sync_int[7]_net_1\, \sync_int[8]_net_1\, 
        \sync_int[9]_net_1\ : std_logic;

begin 


    \sync_int[9]\ : SLE
      port map(D => wptr_gray(9), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[9]_net_1\);
    
    \sync_int[4]\ : SLE
      port map(D => wptr_gray(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[4]_net_1\);
    
    \sync_out_xhdl1[10]\ : SLE
      port map(D => \sync_int[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(10));
    
    \sync_int[1]\ : SLE
      port map(D => wptr_gray(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[1]_net_1\);
    
    \sync_int[11]\ : SLE
      port map(D => wptr_gray(11), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[11]_net_1\);
    
    \sync_out_xhdl1[6]\ : SLE
      port map(D => \sync_int[6]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(6));
    
    \sync_out_xhdl1[3]\ : SLE
      port map(D => \sync_int[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(3));
    
    \sync_int[6]\ : SLE
      port map(D => wptr_gray(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[6]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \sync_out_xhdl1[11]\ : SLE
      port map(D => \sync_int[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(11));
    
    \sync_int[13]\ : SLE
      port map(D => wptr_gray(13), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[13]_net_1\);
    
    \sync_int[3]\ : SLE
      port map(D => wptr_gray(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[3]_net_1\);
    
    \sync_int[12]\ : SLE
      port map(D => wptr_gray(12), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[12]_net_1\);
    
    \sync_out_xhdl1[4]\ : SLE
      port map(D => \sync_int[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(4));
    
    \sync_int[0]\ : SLE
      port map(D => wptr_gray(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[0]_net_1\);
    
    \sync_out_xhdl1[1]\ : SLE
      port map(D => \sync_int[1]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(1));
    
    \sync_int[5]\ : SLE
      port map(D => wptr_gray(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[5]_net_1\);
    
    \sync_int[2]\ : SLE
      port map(D => wptr_gray(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[2]_net_1\);
    
    \sync_out_xhdl1[12]\ : SLE
      port map(D => \sync_int[12]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(12));
    
    \sync_out_xhdl1[9]\ : SLE
      port map(D => \sync_int[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(9));
    
    \sync_out_xhdl1[2]\ : SLE
      port map(D => \sync_int[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(2));
    
    \sync_int[8]\ : SLE
      port map(D => wptr_gray(8), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[8]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sync_out_xhdl1[7]\ : SLE
      port map(D => \sync_int[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(7));
    
    \sync_out_xhdl1[5]\ : SLE
      port map(D => \sync_int[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(5));
    
    \sync_out_xhdl1[0]\ : SLE
      port map(D => \sync_int[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(0));
    
    \sync_out_xhdl1[8]\ : SLE
      port map(D => \sync_int[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(8));
    
    \sync_int[7]\ : SLE
      port map(D => wptr_gray(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[7]_net_1\);
    
    \sync_int[10]\ : SLE
      port map(D => wptr_gray(10), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[10]_net_1\);
    
    \sync_out_xhdl1[13]\ : SLE
      port map(D => \sync_int[13]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_bin_sync_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_2 is

    port( rptr_gray           : in    std_logic_vector(13 downto 0);
          rptr_gray_sync      : out   std_logic_vector(12 downto 0);
          rptr_bin_sync_0     : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          irx_fifo_rst_i      : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_2;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_2 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \sync_int[13]_net_1\, GND_net_1, 
        \sync_int[12]_net_1\, \sync_int[0]_net_1\, 
        \sync_int[1]_net_1\, \sync_int[2]_net_1\, 
        \sync_int[3]_net_1\, \sync_int[4]_net_1\, 
        \sync_int[5]_net_1\, \sync_int[6]_net_1\, 
        \sync_int[7]_net_1\, \sync_int[8]_net_1\, 
        \sync_int[9]_net_1\, \sync_int[10]_net_1\, 
        \sync_int[11]_net_1\ : std_logic;

begin 


    \sync_int[9]\ : SLE
      port map(D => rptr_gray(9), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[9]_net_1\);
    
    \sync_int[4]\ : SLE
      port map(D => rptr_gray(4), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[4]_net_1\);
    
    \sync_out_xhdl1[10]\ : SLE
      port map(D => \sync_int[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(10));
    
    \sync_int[1]\ : SLE
      port map(D => rptr_gray(1), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[1]_net_1\);
    
    \sync_int[11]\ : SLE
      port map(D => rptr_gray(11), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[11]_net_1\);
    
    \sync_out_xhdl1[6]\ : SLE
      port map(D => \sync_int[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(6));
    
    \sync_out_xhdl1[3]\ : SLE
      port map(D => \sync_int[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(3));
    
    \sync_int[6]\ : SLE
      port map(D => rptr_gray(6), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[6]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \sync_out_xhdl1[11]\ : SLE
      port map(D => \sync_int[11]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(11));
    
    \sync_int[13]\ : SLE
      port map(D => rptr_gray(13), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[13]_net_1\);
    
    \sync_int[3]\ : SLE
      port map(D => rptr_gray(3), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[3]_net_1\);
    
    \sync_int[12]\ : SLE
      port map(D => rptr_gray(12), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[12]_net_1\);
    
    \sync_out_xhdl1[4]\ : SLE
      port map(D => \sync_int[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(4));
    
    \sync_int[0]\ : SLE
      port map(D => rptr_gray(0), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[0]_net_1\);
    
    \sync_out_xhdl1[1]\ : SLE
      port map(D => \sync_int[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(1));
    
    \sync_int[5]\ : SLE
      port map(D => rptr_gray(5), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[5]_net_1\);
    
    \sync_int[2]\ : SLE
      port map(D => rptr_gray(2), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[2]_net_1\);
    
    \sync_out_xhdl1[12]\ : SLE
      port map(D => \sync_int[12]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(12));
    
    \sync_out_xhdl1[9]\ : SLE
      port map(D => \sync_int[9]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(9));
    
    \sync_out_xhdl1[2]\ : SLE
      port map(D => \sync_int[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(2));
    
    \sync_int[8]\ : SLE
      port map(D => rptr_gray(8), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[8]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sync_out_xhdl1[7]\ : SLE
      port map(D => \sync_int[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(7));
    
    \sync_out_xhdl1[5]\ : SLE
      port map(D => \sync_int[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(5));
    
    \sync_out_xhdl1[0]\ : SLE
      port map(D => \sync_int[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(0));
    
    \sync_out_xhdl1[8]\ : SLE
      port map(D => \sync_int[8]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(8));
    
    \sync_int[7]\ : SLE
      port map(D => rptr_gray(7), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[7]_net_1\);
    
    \sync_int[10]\ : SLE
      port map(D => rptr_gray(10), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[10]_net_1\);
    
    \sync_out_xhdl1[13]\ : SLE
      port map(D => \sync_int[13]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_bin_sync_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_5 is

    port( rptr_bin_sync  : inout std_logic_vector(13 downto 0) := (others => 'Z');
          rptr_gray_sync : in    std_logic_vector(12 downto 0);
          bin_N_6_i      : out   std_logic;
          bin_N_4_0_i    : out   std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_5;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_5 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \bin_m5_5\, \bin_m5_4\, \bin_m3_0_3\, \bin_N_4_0_i\, 
        GND_net_1, VCC_net_1 : std_logic;

begin 

    bin_N_4_0_i <= \bin_N_4_0_i\;

    bin_m5_4 : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(4), B => rptr_gray_sync(6), C
         => rptr_gray_sync(5), D => rptr_gray_sync(10), Y => 
        \bin_m5_4\);
    
    \bin_out_xhdl1_0_a2[10]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(12), B => rptr_gray_sync(10), 
        C => rptr_gray_sync(11), D => rptr_bin_sync(13), Y => 
        rptr_bin_sync(10));
    
    \bin_out_xhdl1_0_a2[8]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(8), B => rptr_gray_sync(9), C
         => rptr_bin_sync(10), Y => rptr_bin_sync(8));
    
    bin_m5_5 : CFG4
      generic map(INIT => x"9669")

      port map(A => rptr_gray_sync(8), B => rptr_gray_sync(9), C
         => rptr_gray_sync(7), D => rptr_gray_sync(11), Y => 
        \bin_m5_5\);
    
    bin_m3_0_3 : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(7), B => rptr_gray_sync(9), C
         => rptr_gray_sync(6), D => rptr_gray_sync(10), Y => 
        \bin_m3_0_3\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \bin_out_xhdl1_0_a2[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(3), B => rptr_gray_sync(2), Y
         => rptr_bin_sync(2));
    
    \bin_out_xhdl1_0_a2[1]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(1), B => rptr_gray_sync(2), C
         => rptr_bin_sync(3), Y => rptr_bin_sync(1));
    
    \bin_out_xhdl1_0_a2[0]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(1), B => rptr_gray_sync(0), C
         => rptr_bin_sync(3), D => rptr_gray_sync(2), Y => 
        rptr_bin_sync(0));
    
    \bin_out_xhdl1_i_o2_RNIO8EI1[12]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(8), B => rptr_gray_sync(11), C
         => rptr_bin_sync(12), D => \bin_m3_0_3\, Y => 
        \bin_N_4_0_i\);
    
    \bin_out_xhdl1_i_o2[11]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(11), B => rptr_bin_sync(13), C
         => rptr_gray_sync(12), Y => rptr_bin_sync(11));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \bin_out_xhdl1_0_a2[7]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(9), B => rptr_bin_sync(10), C
         => rptr_gray_sync(7), D => rptr_gray_sync(8), Y => 
        rptr_bin_sync(7));
    
    \bin_out_xhdl1_0_a2[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \bin_N_4_0_i\, B => rptr_gray_sync(5), Y => 
        rptr_bin_sync(5));
    
    \bin_out_xhdl1_i_o2_RNIBP3N1[12]\ : CFG3
      generic map(INIT => x"69")

      port map(A => \bin_m5_5\, B => \bin_m5_4\, C => 
        rptr_bin_sync(12), Y => bin_N_6_i);
    
    \bin_out_xhdl1_i_o2[12]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(13), B => rptr_gray_sync(12), Y
         => rptr_bin_sync(12));
    
    \bin_out_xhdl1_0_a2[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(10), B => rptr_gray_sync(9), Y
         => rptr_bin_sync(9));
    
    \bin_out_xhdl1_0_a2[3]\ : CFG4
      generic map(INIT => x"9669")

      port map(A => rptr_bin_sync(12), B => \bin_m5_5\, C => 
        rptr_gray_sync(3), D => \bin_m5_4\, Y => rptr_bin_sync(3));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_2 is

    port( fifo_MEMRADDR             : out   std_logic_vector(12 downto 0);
          fifo_MEMWADDR             : out   std_logic_vector(12 downto 0);
          iRX_FIFO_wr_en_0_0        : in    std_logic;
          iRX_FIFO_rd_en_0          : in    std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          RX_FIFO_TxColDetDis_wr_en : in    std_logic;
          fifo_MEMRE                : out   std_logic;
          fifo_MEMWE                : out   std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          irx_fifo_rst_i            : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_2;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_2 is 

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_6
    port( wptr_bin_sync  : inout   std_logic_vector(13 downto 0);
          wptr_gray_sync : in    std_logic_vector(12 downto 0) := (others => 'U')
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_3
    port( wptr_gray                 : in    std_logic_vector(13 downto 0) := (others => 'U');
          wptr_gray_sync            : out   std_logic_vector(12 downto 0);
          wptr_bin_sync_0           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          irx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_2
    port( rptr_gray           : in    std_logic_vector(13 downto 0) := (others => 'U');
          rptr_gray_sync      : out   std_logic_vector(12 downto 0);
          rptr_bin_sync_0     : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          irx_fifo_rst_i      : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_5
    port( rptr_bin_sync  : inout   std_logic_vector(13 downto 0);
          rptr_gray_sync : in    std_logic_vector(12 downto 0) := (others => 'U');
          bin_N_6_i      : out   std_logic;
          bin_N_4_0_i    : out   std_logic
        );
  end component;

    signal \rptr[0]_net_1\, \rptr_s[0]\, \wptr[0]_net_1\, 
        \wptr_s[0]\, \fifo_MEMRADDR[0]\, \fifo_MEMRADDR_i[0]\, 
        \fifo_MEMWADDR[0]\, \fifo_MEMWADDR_i[0]\, 
        \rptr_gray[1]_net_1\, VCC_net_1, \rptr_gray_1[1]_net_1\, 
        GND_net_1, \rptr_gray[2]_net_1\, \rptr_gray_1[2]_net_1\, 
        \rptr_gray[3]_net_1\, \rptr_gray_1[3]_net_1\, 
        \rptr_gray[4]_net_1\, \rptr_gray_1[4]_net_1\, 
        \rptr_gray[5]_net_1\, \rptr_gray_1[5]_net_1\, 
        \rptr_gray[6]_net_1\, \rptr_gray_1[6]_net_1\, 
        \rptr_gray[7]_net_1\, \rptr_gray_1[7]_net_1\, 
        \rptr_gray[8]_net_1\, \rptr_gray_1[8]_net_1\, 
        \rptr_gray[9]_net_1\, \rptr_gray_1[9]_net_1\, 
        \rptr_gray[10]_net_1\, \rptr_gray_1[10]_net_1\, 
        \rptr_gray[11]_net_1\, \rptr_gray_1[11]_net_1\, 
        \rptr_gray[12]_net_1\, \rptr_gray_1[12]_net_1\, 
        \rptr_gray[13]_net_1\, \rptr[13]_net_1\, 
        \wptr_gray[0]_net_1\, \wptr_gray_1[0]_net_1\, 
        \wptr_gray[1]_net_1\, \wptr_gray_1[1]_net_1\, 
        \wptr_gray[2]_net_1\, \wptr_gray_1[2]_net_1\, 
        \wptr_gray[3]_net_1\, \wptr_gray_1[3]_net_1\, 
        \wptr_gray[4]_net_1\, \wptr_gray_1[4]_net_1\, 
        \wptr_gray[5]_net_1\, \wptr_gray_1[5]_net_1\, 
        \wptr_gray[6]_net_1\, \wptr_gray_1[6]_net_1\, 
        \wptr_gray[7]_net_1\, \wptr_gray_1[7]_net_1\, 
        \wptr_gray[8]_net_1\, \wptr_gray_1[8]_net_1\, 
        \wptr_gray[9]_net_1\, \wptr_gray_1[9]_net_1\, 
        \wptr_gray[10]_net_1\, \wptr_gray_1[10]_net_1\, 
        \wptr_gray[11]_net_1\, \wptr_gray_1[11]_net_1\, 
        \wptr_gray[12]_net_1\, \wptr_gray_1[12]_net_1\, 
        \wptr_gray[13]_net_1\, \wptr[13]_net_1\, 
        \rptr_gray[0]_net_1\, \rptr_gray_1[0]_net_1\, rdiff_bus, 
        \wptr_bin_sync[0]\, \wptr_bin_sync2[1]_net_1\, 
        \wptr_bin_sync[1]\, \wptr_bin_sync2[2]_net_1\, 
        \wptr_bin_sync[2]\, \wptr_bin_sync2[3]_net_1\, 
        \wptr_bin_sync[3]\, \wptr_bin_sync2[4]_net_1\, 
        \wptr_bin_sync[4]\, \wptr_bin_sync2[5]_net_1\, 
        \wptr_bin_sync[5]\, \wptr_bin_sync2[6]_net_1\, 
        \wptr_bin_sync[6]\, \wptr_bin_sync2[7]_net_1\, 
        \wptr_bin_sync[7]\, \wptr_bin_sync2[8]_net_1\, 
        \wptr_bin_sync[8]\, \wptr_bin_sync2[9]_net_1\, 
        \wptr_bin_sync[9]\, \wptr_bin_sync2[10]_net_1\, 
        \wptr_bin_sync[10]\, \wptr_bin_sync2[11]_net_1\, 
        \wptr_bin_sync[11]\, \wptr_bin_sync2[12]_net_1\, 
        \wptr_bin_sync[12]\, \wptr_bin_sync2[13]_net_1\, 
        \wptr_bin_sync[13]\, \rptr_bin_sync2[9]_net_1\, 
        \rptr_bin_sync[9]\, \rptr_bin_sync2[10]_net_1\, 
        \rptr_bin_sync[10]\, \rptr_bin_sync2[11]_net_1\, 
        \rptr_bin_sync[11]\, \rptr_bin_sync2[12]_net_1\, 
        \rptr_bin_sync[12]\, \rptr_bin_sync2[13]_net_1\, 
        \rptr_bin_sync[13]\, \fifo_MEMWADDR[7]\, 
        \memwaddr_r_2[7]_net_1\, \fifo_MEMWE\, \fifo_MEMWADDR[8]\, 
        \memwaddr_r_2[8]_net_1\, \fifo_MEMWADDR[9]\, 
        \memwaddr_r_2[9]_net_1\, \fifo_MEMWADDR[10]\, 
        \memwaddr_r_2[10]_net_1\, \fifo_MEMWADDR[11]\, 
        \memwaddr_r_2[11]_net_1\, \fifo_MEMWADDR[12]\, 
        \memwaddr_r_2[12]_net_1\, \rptr_bin_sync2[0]_net_1\, 
        \rptr_bin_sync[0]\, \rptr_bin_sync2[1]_net_1\, 
        \rptr_bin_sync[1]\, \rptr_bin_sync2[2]_net_1\, 
        \rptr_bin_sync[2]\, \rptr_bin_sync2[3]_net_1\, 
        \rptr_bin_sync[3]\, \rptr_bin_sync2[4]_net_1\, bin_N_6_i, 
        \rptr_bin_sync2[5]_net_1\, \rptr_bin_sync[5]\, 
        \rptr_bin_sync2[6]_net_1\, bin_N_4_0_i, 
        \rptr_bin_sync2[7]_net_1\, \rptr_bin_sync[7]\, 
        \rptr_bin_sync2[8]_net_1\, \rptr_bin_sync[8]\, 
        \fifo_MEMRADDR[5]\, \memraddr_r_2[5]_net_1\, \fifo_MEMRE\, 
        \fifo_MEMRADDR[6]\, un1_memraddr_r_cry_6_S_2, 
        \fifo_MEMRADDR[7]\, \memraddr_r_2[7]_net_1\, 
        \fifo_MEMRADDR[8]\, \memraddr_r_2[8]_net_1\, 
        \fifo_MEMRADDR[9]\, \memraddr_r_2[9]_net_1\, 
        \fifo_MEMRADDR[10]\, \memraddr_r_2[10]_net_1\, 
        \fifo_MEMRADDR[11]\, \memraddr_r_2[11]_net_1\, 
        \fifo_MEMRADDR[12]\, \memraddr_r_2[12]_net_1\, 
        \fifo_MEMWADDR[1]\, un1_memwaddr_r_cry_1_S_2, 
        \fifo_MEMWADDR[2]\, un1_memwaddr_r_cry_2_S_2, 
        \fifo_MEMWADDR[3]\, un1_memwaddr_r_cry_3_S_2, 
        \fifo_MEMWADDR[4]\, un1_memwaddr_r_cry_4_S_2, 
        \fifo_MEMWADDR[5]\, \memwaddr_r_2[5]_net_1\, 
        \fifo_MEMWADDR[6]\, un1_memwaddr_r_cry_6_S_2, 
        \fifo_MEMRADDR[1]\, un1_memraddr_r_cry_1_S_2, 
        \fifo_MEMRADDR[2]\, un1_memraddr_r_cry_2_S_2, 
        \fifo_MEMRADDR[3]\, un1_memraddr_r_cry_3_S_2, 
        \fifo_MEMRADDR[4]\, un1_memraddr_r_cry_4_S_2, 
        \iRX_FIFO_Full_0\, fulli, N_6_i, N_5_i, 
        \iRX_FIFO_Empty_0\, empty_r_3, \wptr[1]_net_1\, 
        \wptr_s[1]\, \wptr[2]_net_1\, \wptr_s[2]\, 
        \wptr[3]_net_1\, \wptr_s[3]\, \wptr[4]_net_1\, 
        \wptr_s[4]\, \wptr[5]_net_1\, \wptr_s[5]\, 
        \wptr[6]_net_1\, \wptr_s[6]\, \wptr[7]_net_1\, 
        \wptr_s[7]\, \wptr[8]_net_1\, \wptr_s[8]\, 
        \wptr[9]_net_1\, \wptr_s[9]\, \wptr[10]_net_1\, 
        \wptr_s[10]\, \wptr[11]_net_1\, \wptr_s[11]\, 
        \wptr[12]_net_1\, \wptr_s[12]\, \wptr_s[13]_net_1\, 
        \rptr[1]_net_1\, \rptr_s[1]\, \rptr[2]_net_1\, 
        \rptr_s[2]\, \rptr[3]_net_1\, \rptr_s[3]\, 
        \rptr[4]_net_1\, \rptr_s[4]\, \rptr[5]_net_1\, 
        \rptr_s[5]\, \rptr[6]_net_1\, \rptr_s[6]\, 
        \rptr[7]_net_1\, \rptr_s[7]\, \rptr[8]_net_1\, 
        \rptr_s[8]\, \rptr[9]_net_1\, \rptr_s[9]\, 
        \rptr[10]_net_1\, \rptr_s[10]\, \rptr[11]_net_1\, 
        \rptr_s[11]\, \rptr[12]_net_1\, \rptr_s[12]\, 
        \rptr_s[13]_net_1\, \rdiff_bus_cry_0\, 
        rdiff_bus_cry_0_Y_3, \rdiff_bus_cry_1\, \rdiff_bus[1]\, 
        \rdiff_bus_cry_2\, \rdiff_bus[2]\, \rdiff_bus_cry_3\, 
        \rdiff_bus[3]\, \rdiff_bus_cry_4\, \rdiff_bus[4]\, 
        \rdiff_bus_cry_5\, \rdiff_bus[5]\, \rdiff_bus_cry_6\, 
        \rdiff_bus[6]\, \rdiff_bus_cry_7\, \rdiff_bus[7]\, 
        \rdiff_bus_cry_8\, \rdiff_bus[8]\, \rdiff_bus_cry_9\, 
        \rdiff_bus[9]\, \rdiff_bus_cry_10\, \rdiff_bus[10]\, 
        \rdiff_bus_cry_11\, \rdiff_bus[11]\, \rdiff_bus[13]\, 
        \rdiff_bus_cry_12\, \rdiff_bus[12]\, \wdiff_bus_cry_0\, 
        wdiff_bus_cry_0_Y_3, \wdiff_bus_cry_1\, \wdiff_bus[1]\, 
        \wdiff_bus_cry_2\, \wdiff_bus[2]\, \wdiff_bus_cry_3\, 
        \wdiff_bus[3]\, \wdiff_bus_cry_4\, \wdiff_bus[4]\, 
        \wdiff_bus_cry_5\, \wdiff_bus[5]\, \wdiff_bus_cry_6\, 
        \wdiff_bus[6]\, \wdiff_bus_cry_7\, \wdiff_bus[7]\, 
        \wdiff_bus_cry_8\, \wdiff_bus[8]\, \wdiff_bus_cry_9\, 
        \wdiff_bus[9]\, \wdiff_bus_cry_10\, \wdiff_bus[10]\, 
        \wdiff_bus_cry_11\, \wdiff_bus[11]\, \wdiff_bus[13]\, 
        \wdiff_bus_cry_12\, \wdiff_bus[12]\, rptr_s_902_FCO, 
        \rptr_cry[1]_net_1\, \rptr_cry[2]_net_1\, 
        \rptr_cry[3]_net_1\, \rptr_cry[4]_net_1\, 
        \rptr_cry[5]_net_1\, \rptr_cry[6]_net_1\, 
        \rptr_cry[7]_net_1\, \rptr_cry[8]_net_1\, 
        \rptr_cry[9]_net_1\, \rptr_cry[10]_net_1\, 
        \rptr_cry[11]_net_1\, \rptr_cry[12]_net_1\, 
        wptr_s_903_FCO, \wptr_cry[1]_net_1\, \wptr_cry[2]_net_1\, 
        \wptr_cry[3]_net_1\, \wptr_cry[4]_net_1\, 
        \wptr_cry[5]_net_1\, \wptr_cry[6]_net_1\, 
        \wptr_cry[7]_net_1\, \wptr_cry[8]_net_1\, 
        \wptr_cry[9]_net_1\, \wptr_cry[10]_net_1\, 
        \wptr_cry[11]_net_1\, \wptr_cry[12]_net_1\, 
        un1_memraddr_r_s_1_929_FCO, \un1_memraddr_r_cry_1\, 
        \un1_memraddr_r_cry_2\, \un1_memraddr_r_cry_3\, 
        \un1_memraddr_r_cry_4\, \un1_memraddr_r_cry_5\, 
        un1_memraddr_r_cry_5_S_2, \un1_memraddr_r_cry_6\, 
        \un1_memraddr_r_cry_7\, un1_memraddr_r_cry_7_S_2, 
        \un1_memraddr_r_cry_8\, un1_memraddr_r_cry_8_S_2, 
        \un1_memraddr_r_cry_9\, un1_memraddr_r_cry_9_S_2, 
        \un1_memraddr_r_cry_10\, un1_memraddr_r_cry_10_S_2, 
        un1_memraddr_r_s_12_S_2, \un1_memraddr_r_cry_11\, 
        un1_memraddr_r_cry_11_S_2, un1_memwaddr_r_s_1_930_FCO, 
        \un1_memwaddr_r_cry_1\, \un1_memwaddr_r_cry_2\, 
        \un1_memwaddr_r_cry_3\, \un1_memwaddr_r_cry_4\, 
        \un1_memwaddr_r_cry_5\, un1_memwaddr_r_cry_5_S_2, 
        \un1_memwaddr_r_cry_6\, \un1_memwaddr_r_cry_7\, 
        un1_memwaddr_r_cry_7_S_2, \un1_memwaddr_r_cry_8\, 
        un1_memwaddr_r_cry_8_S_2, \un1_memwaddr_r_cry_9\, 
        un1_memwaddr_r_cry_9_S_2, \un1_memwaddr_r_cry_10\, 
        un1_memwaddr_r_cry_10_S_2, un1_memwaddr_r_s_12_S_2, 
        \un1_memwaddr_r_cry_11\, un1_memwaddr_r_cry_11_S_2, 
        \fulli_0_1\, N_12, \fulli_0_a3_3\, un4_re_i_0, un4_we_i_0, 
        empty_r_3_0_a2_9, empty_r_3_0_a2_8, empty_r_3_0_a2_7, 
        un4_re_i_8, un4_re_i_7, un4_we_i_8, un4_we_i_7, 
        un4_re_i_9, un4_we_i_9, empty_r_3_0_a2_6, 
        \fulli_0_a3_0_3\, \wptr_gray_sync[0]\, 
        \wptr_gray_sync[1]\, \wptr_gray_sync[2]\, 
        \wptr_gray_sync[3]\, \wptr_gray_sync[4]\, 
        \wptr_gray_sync[5]\, \wptr_gray_sync[6]\, 
        \wptr_gray_sync[7]\, \wptr_gray_sync[8]\, 
        \wptr_gray_sync[9]\, \wptr_gray_sync[10]\, 
        \wptr_gray_sync[11]\, \wptr_gray_sync[12]\, 
        \rptr_gray_sync[0]\, \rptr_gray_sync[1]\, 
        \rptr_gray_sync[2]\, \rptr_gray_sync[3]\, 
        \rptr_gray_sync[4]\, \rptr_gray_sync[5]\, 
        \rptr_gray_sync[6]\, \rptr_gray_sync[7]\, 
        \rptr_gray_sync[8]\, \rptr_gray_sync[9]\, 
        \rptr_gray_sync[10]\, \rptr_gray_sync[11]\, 
        \rptr_gray_sync[12]\ : std_logic;
    signal nc2, nc1 : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_6
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_6(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_3
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_3(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_2
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_2(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_5
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_5(DEF_ARCH);
begin 

    fifo_MEMRADDR(12) <= \fifo_MEMRADDR[12]\;
    fifo_MEMRADDR(11) <= \fifo_MEMRADDR[11]\;
    fifo_MEMRADDR(10) <= \fifo_MEMRADDR[10]\;
    fifo_MEMRADDR(9) <= \fifo_MEMRADDR[9]\;
    fifo_MEMRADDR(8) <= \fifo_MEMRADDR[8]\;
    fifo_MEMRADDR(7) <= \fifo_MEMRADDR[7]\;
    fifo_MEMRADDR(6) <= \fifo_MEMRADDR[6]\;
    fifo_MEMRADDR(5) <= \fifo_MEMRADDR[5]\;
    fifo_MEMRADDR(4) <= \fifo_MEMRADDR[4]\;
    fifo_MEMRADDR(3) <= \fifo_MEMRADDR[3]\;
    fifo_MEMRADDR(2) <= \fifo_MEMRADDR[2]\;
    fifo_MEMRADDR(1) <= \fifo_MEMRADDR[1]\;
    fifo_MEMRADDR(0) <= \fifo_MEMRADDR[0]\;
    fifo_MEMWADDR(12) <= \fifo_MEMWADDR[12]\;
    fifo_MEMWADDR(11) <= \fifo_MEMWADDR[11]\;
    fifo_MEMWADDR(10) <= \fifo_MEMWADDR[10]\;
    fifo_MEMWADDR(9) <= \fifo_MEMWADDR[9]\;
    fifo_MEMWADDR(8) <= \fifo_MEMWADDR[8]\;
    fifo_MEMWADDR(7) <= \fifo_MEMWADDR[7]\;
    fifo_MEMWADDR(6) <= \fifo_MEMWADDR[6]\;
    fifo_MEMWADDR(5) <= \fifo_MEMWADDR[5]\;
    fifo_MEMWADDR(4) <= \fifo_MEMWADDR[4]\;
    fifo_MEMWADDR(3) <= \fifo_MEMWADDR[3]\;
    fifo_MEMWADDR(2) <= \fifo_MEMWADDR[2]\;
    fifo_MEMWADDR(1) <= \fifo_MEMWADDR[1]\;
    fifo_MEMWADDR(0) <= \fifo_MEMWADDR[0]\;
    iRX_FIFO_Empty_0 <= \iRX_FIFO_Empty_0\;
    iRX_FIFO_Full_0 <= \iRX_FIFO_Full_0\;
    fifo_MEMRE <= \fifo_MEMRE\;
    fifo_MEMWE <= \fifo_MEMWE\;

    \rptr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[4]_net_1\, S
         => \rptr_s[5]\, Y => OPEN, FCO => \rptr_cry[5]_net_1\);
    
    \memwaddr_r_2[9]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_9_S_2, D => un4_we_i_9, Y => 
        \memwaddr_r_2[9]_net_1\);
    
    wdiff_bus_cry_8 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[8]_net_1\, B => 
        \rptr_bin_sync2[8]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_7\, S => \wdiff_bus[8]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_8\);
    
    \wptr_bin_sync2[12]\ : SLE
      port map(D => \wptr_bin_sync[12]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[12]_net_1\);
    
    wdiff_bus_cry_11 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[11]_net_1\, B => 
        \rptr_bin_sync2[11]_net_1\, C => GND_net_1, D => 
        GND_net_1, FCI => \wdiff_bus_cry_10\, S => 
        \wdiff_bus[11]\, Y => OPEN, FCO => \wdiff_bus_cry_11\);
    
    \wptr_gray[4]\ : SLE
      port map(D => \wptr_gray_1[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[4]_net_1\);
    
    \rptr_gray_1[3]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[3]_net_1\, B => \rptr[4]_net_1\, Y => 
        \rptr_gray_1[3]_net_1\);
    
    \rptr_bin_sync2[6]\ : SLE
      port map(D => bin_N_4_0_i, CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_bin_sync2[6]_net_1\);
    
    \rptr[1]\ : SLE
      port map(D => \rptr_s[1]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[1]_net_1\);
    
    fulli_0_a3_0_3 : CFG4
      generic map(INIT => x"8000")

      port map(A => \wdiff_bus[2]\, B => 
        RX_FIFO_TxColDetDis_wr_en, C => iRX_FIFO_wr_en_0_0, D => 
        \wdiff_bus[3]\, Y => \fulli_0_a3_0_3\);
    
    \wptr_gray_1[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[9]_net_1\, B => \wptr[10]_net_1\, Y => 
        \wptr_gray_1[9]_net_1\);
    
    \rptr_gray_1[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[5]_net_1\, B => \rptr[6]_net_1\, Y => 
        \rptr_gray_1[5]_net_1\);
    
    \rptr_gray[9]\ : SLE
      port map(D => \rptr_gray_1[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[9]_net_1\);
    
    un1_memwaddr_r_cry_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_6\, 
        S => un1_memwaddr_r_cry_7_S_2, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_7\);
    
    \rptr_gray[8]\ : SLE
      port map(D => \rptr_gray_1[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[8]_net_1\);
    
    un1_memraddr_r_cry_11 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[11]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_10\, 
        S => un1_memraddr_r_cry_11_S_2, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_11\);
    
    \rptr_gray_1[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[2]_net_1\, B => \rptr[3]_net_1\, Y => 
        \rptr_gray_1[2]_net_1\);
    
    \rptr_bin_sync2[7]\ : SLE
      port map(D => \rptr_bin_sync[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[7]_net_1\);
    
    \memwaddr_r[1]\ : SLE
      port map(D => un1_memwaddr_r_cry_1_S_2, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[1]\);
    
    \wptr_gray_1[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[7]_net_1\, B => \wptr[8]_net_1\, Y => 
        \wptr_gray_1[7]_net_1\);
    
    \rptr_gray[13]\ : SLE
      port map(D => \rptr[13]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[13]_net_1\);
    
    \memraddr_r[0]\ : SLE
      port map(D => \fifo_MEMRADDR_i[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[0]\);
    
    \memraddr_r_2[9]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => 
        un1_memraddr_r_cry_9_S_2, D => un4_re_i_9, Y => 
        \memraddr_r_2[9]_net_1\);
    
    \wptr[0]\ : SLE
      port map(D => \wptr_s[0]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[0]_net_1\);
    
    \rptr_bin_sync2[8]\ : SLE
      port map(D => \rptr_bin_sync[8]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[8]_net_1\);
    
    \rptr_gray_1[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[1]_net_1\, B => \rptr[2]_net_1\, Y => 
        \rptr_gray_1[1]_net_1\);
    
    \rptr_gray[10]\ : SLE
      port map(D => \rptr_gray_1[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[10]_net_1\);
    
    \wptr_gray_1[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[0]_net_1\, B => \wptr[1]_net_1\, Y => 
        \wptr_gray_1[0]_net_1\);
    
    wdiff_bus_cry_9 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[9]_net_1\, B => 
        \rptr_bin_sync2[9]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_8\, S => \wdiff_bus[9]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_9\);
    
    \rptr[5]\ : SLE
      port map(D => \rptr_s[5]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[5]_net_1\);
    
    \rptr_gray[3]\ : SLE
      port map(D => \rptr_gray_1[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[3]_net_1\);
    
    \rptr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[5]_net_1\, S
         => \rptr_s[6]\, Y => OPEN, FCO => \rptr_cry[6]_net_1\);
    
    \wptr_gray[3]\ : SLE
      port map(D => \wptr_gray_1[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[3]_net_1\);
    
    \rptr_gray_1[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[10]_net_1\, B => \rptr[11]_net_1\, Y
         => \rptr_gray_1[10]_net_1\);
    
    un1_memraddr_r_cry_10 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_9\, 
        S => un1_memraddr_r_cry_10_S_2, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_10\);
    
    \rptr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[7]_net_1\, S
         => \rptr_s[8]\, Y => OPEN, FCO => \rptr_cry[8]_net_1\);
    
    \rptr[7]\ : SLE
      port map(D => \rptr_s[7]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[7]_net_1\);
    
    rdiff_bus_cry_4 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[4]_net_1\, B => 
        \rptr[4]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_3\, S => \rdiff_bus[4]\, Y => OPEN, FCO
         => \rdiff_bus_cry_4\);
    
    \rptr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[9]_net_1\, S
         => \rptr_s[10]\, Y => OPEN, FCO => \rptr_cry[10]_net_1\);
    
    \rptr_bin_sync2[12]\ : SLE
      port map(D => \rptr_bin_sync[12]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[12]_net_1\);
    
    memwe_0_a3 : CFG3
      generic map(INIT => x"20")

      port map(A => RX_FIFO_TxColDetDis_wr_en, B => 
        \iRX_FIFO_Full_0\, C => iRX_FIFO_wr_en_0_0, Y => 
        \fifo_MEMWE\);
    
    \rptr_bin_sync2[0]\ : SLE
      port map(D => \rptr_bin_sync[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[0]_net_1\);
    
    \L1.empty_r_3_0_a2_7\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \rdiff_bus[1]\, B => \rdiff_bus[4]\, C => 
        \rdiff_bus[3]\, D => \rdiff_bus[2]\, Y => 
        empty_r_3_0_a2_7);
    
    \wptr[11]\ : SLE
      port map(D => \wptr_s[11]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[11]_net_1\);
    
    un1_memwaddr_r_s_1_930 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[0]\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => un1_memwaddr_r_s_1_930_FCO);
    
    rdiff_bus_cry_1 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[1]_net_1\, B => 
        \rptr[1]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_0\, S => \rdiff_bus[1]\, Y => OPEN, FCO
         => \rdiff_bus_cry_1\);
    
    \memraddr_r[1]\ : SLE
      port map(D => un1_memraddr_r_cry_1_S_2, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[1]\);
    
    \L1.empty_r_3_0_a2_9\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \rdiff_bus[9]\, B => \rdiff_bus[10]\, C => 
        \rdiff_bus[11]\, D => \rdiff_bus[12]\, Y => 
        empty_r_3_0_a2_9);
    
    \rptr_bin_sync2[2]\ : SLE
      port map(D => \rptr_bin_sync[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[2]_net_1\);
    
    \memraddr_r_2[7]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => 
        un1_memraddr_r_cry_7_S_2, D => un4_re_i_9, Y => 
        \memraddr_r_2[7]_net_1\);
    
    un1_memwaddr_r_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_5\, 
        S => un1_memwaddr_r_cry_6_S_2, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_6\);
    
    rdiff_bus_cry_6 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[6]_net_1\, B => 
        \rptr[6]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_5\, S => \rdiff_bus[6]\, Y => OPEN, FCO
         => \rdiff_bus_cry_6\);
    
    \memwaddr_r_2[10]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_10_S_2, D => un4_we_i_9, Y => 
        \memwaddr_r_2[10]_net_1\);
    
    \memraddr_r_2[5]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => 
        un1_memraddr_r_cry_5_S_2, D => un4_re_i_9, Y => 
        \memraddr_r_2[5]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    un1_memwaddr_r_cry_9 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[9]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_8\, 
        S => un1_memwaddr_r_cry_9_S_2, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_9\);
    
    \rptr_gray[1]\ : SLE
      port map(D => \rptr_gray_1[1]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[1]_net_1\);
    
    \memwaddr_r[7]\ : SLE
      port map(D => \memwaddr_r_2[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[7]\);
    
    \wptr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[3]_net_1\, S
         => \wptr_s[4]\, Y => OPEN, FCO => \wptr_cry[4]_net_1\);
    
    \wptr_gray_1[12]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[13]_net_1\, B => \wptr[12]_net_1\, Y
         => \wptr_gray_1[12]_net_1\);
    
    \wptr[12]\ : SLE
      port map(D => \wptr_s[12]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[12]_net_1\);
    
    \wptr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[9]_net_1\, S
         => \wptr_s[10]\, Y => OPEN, FCO => \wptr_cry[10]_net_1\);
    
    wdiff_bus_cry_5 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[5]_net_1\, B => 
        \rptr_bin_sync2[5]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_4\, S => \wdiff_bus[5]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_5\);
    
    \rptr_gray[12]\ : SLE
      port map(D => \rptr_gray_1[12]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[12]_net_1\);
    
    \memwaddr_r[4]\ : SLE
      port map(D => un1_memwaddr_r_cry_4_S_2, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[4]\);
    
    \wptr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[1]_net_1\, S
         => \wptr_s[2]\, Y => OPEN, FCO => \wptr_cry[2]_net_1\);
    
    \memraddr_r_2[10]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => 
        un1_memraddr_r_cry_10_S_2, D => un4_re_i_9, Y => 
        \memraddr_r_2[10]_net_1\);
    
    rdiff_bus_cry_11 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[11]_net_1\, B => 
        \rptr[11]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_10\, S => \rdiff_bus[11]\, Y => OPEN, FCO
         => \rdiff_bus_cry_11\);
    
    wdiff_bus_cry_0 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[0]_net_1\, B => 
        \rptr_bin_sync2[0]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => VCC_net_1, S => OPEN, Y => wdiff_bus_cry_0_Y_3, 
        FCO => \wdiff_bus_cry_0\);
    
    \wptr[1]\ : SLE
      port map(D => \wptr_s[1]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[1]_net_1\);
    
    \rptr_bin_sync2[4]\ : SLE
      port map(D => bin_N_6_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[4]_net_1\);
    
    \wptr_bin_sync2[6]\ : SLE
      port map(D => \wptr_bin_sync[6]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[6]_net_1\);
    
    \rptr[3]\ : SLE
      port map(D => \rptr_s[3]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[3]_net_1\);
    
    \wptr_gray[13]\ : SLE
      port map(D => \wptr[13]_net_1\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr_gray[13]_net_1\);
    
    \wptr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[2]_net_1\, S
         => \wptr_s[3]\, Y => OPEN, FCO => \wptr_cry[3]_net_1\);
    
    \L1.empty_r_3_0_a2_8\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \rdiff_bus[5]\, B => \rdiff_bus[6]\, C => 
        \rdiff_bus[7]\, D => \rdiff_bus[8]\, Y => 
        empty_r_3_0_a2_8);
    
    \rptr[6]\ : SLE
      port map(D => \rptr_s[6]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[6]_net_1\);
    
    rdiff_bus_cry_8 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[8]_net_1\, B => 
        \rptr[8]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_7\, S => \rdiff_bus[8]\, Y => OPEN, FCO
         => \rdiff_bus_cry_8\);
    
    \wptr_gray[10]\ : SLE
      port map(D => \wptr_gray_1[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[10]_net_1\);
    
    rdiff_bus_cry_7 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[7]_net_1\, B => 
        \rptr[7]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_6\, S => \rdiff_bus[7]\, Y => OPEN, FCO
         => \rdiff_bus_cry_7\);
    
    \wptr_bin_sync2[7]\ : SLE
      port map(D => \wptr_bin_sync[7]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[7]_net_1\);
    
    \rptr_gray_1[11]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[11]_net_1\, B => \rptr[12]_net_1\, Y
         => \rptr_gray_1[11]_net_1\);
    
    \rptr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[8]_net_1\, S
         => \rptr_s[9]\, Y => OPEN, FCO => \rptr_cry[9]_net_1\);
    
    un1_memwaddr_r_cry_1 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[1]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        un1_memwaddr_r_s_1_930_FCO, S => un1_memwaddr_r_cry_1_S_2, 
        Y => OPEN, FCO => \un1_memwaddr_r_cry_1\);
    
    \rptr_gray[5]\ : SLE
      port map(D => \rptr_gray_1[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[5]_net_1\);
    
    un1_memwaddr_r_s_12 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[12]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_11\, 
        S => un1_memwaddr_r_s_12_S_2, Y => OPEN, FCO => OPEN);
    
    \wptr_gray_1[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[2]_net_1\, B => \wptr[3]_net_1\, Y => 
        \wptr_gray_1[2]_net_1\);
    
    \wptr[5]\ : SLE
      port map(D => \wptr_s[5]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[5]_net_1\);
    
    rdiff_bus_cry_5 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[5]_net_1\, B => 
        \rptr[5]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_4\, S => \rdiff_bus[5]\, Y => OPEN, FCO
         => \rdiff_bus_cry_5\);
    
    \wptr_bin_sync2[8]\ : SLE
      port map(D => \wptr_bin_sync[8]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[8]_net_1\);
    
    fulli_0_a3_3 : CFG4
      generic map(INIT => x"8000")

      port map(A => \wdiff_bus[7]\, B => \wdiff_bus[8]\, C => 
        \wdiff_bus[9]\, D => \wdiff_bus[10]\, Y => \fulli_0_a3_3\);
    
    \wptr[7]\ : SLE
      port map(D => \wptr_s[7]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[7]_net_1\);
    
    un1_memwaddr_r_cry_2 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[2]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_1\, 
        S => un1_memwaddr_r_cry_2_S_2, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_2\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \wptr_gray[1]\ : SLE
      port map(D => \wptr_gray_1[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[1]_net_1\);
    
    \rptr_gray_1[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[9]_net_1\, B => \rptr[10]_net_1\, Y => 
        \rptr_gray_1[9]_net_1\);
    
    \rptr_bin_sync2[5]\ : SLE
      port map(D => \rptr_bin_sync[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[5]_net_1\);
    
    \rptr_bin_sync2[1]\ : SLE
      port map(D => \rptr_bin_sync[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[1]_net_1\);
    
    \memwaddr_r[10]\ : SLE
      port map(D => \memwaddr_r_2[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[10]\);
    
    wdiff_bus_cry_7 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[7]_net_1\, B => 
        \rptr_bin_sync2[7]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_6\, S => \wdiff_bus[7]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_7\);
    
    \wptr_bin_sync2[0]\ : SLE
      port map(D => \wptr_bin_sync[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rdiff_bus);
    
    un1_memwaddr_r_cry_8 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[8]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_7\, 
        S => un1_memwaddr_r_cry_8_S_2, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_8\);
    
    \wptr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => wptr_s_903_FCO, S => 
        \wptr_s[1]\, Y => OPEN, FCO => \wptr_cry[1]_net_1\);
    
    un1_memwaddr_r_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_3\, 
        S => un1_memwaddr_r_cry_4_S_2, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_4\);
    
    un1_memwaddr_r_cry_3 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[3]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_2\, 
        S => un1_memwaddr_r_cry_3_S_2, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_3\);
    
    \memraddr_r[8]\ : SLE
      port map(D => \memraddr_r_2[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[8]\);
    
    \rptr[9]\ : SLE
      port map(D => \rptr_s[9]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[9]_net_1\);
    
    \wptr_gray_1[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[6]_net_1\, B => \wptr[7]_net_1\, Y => 
        \wptr_gray_1[6]_net_1\);
    
    \wptr_gray[12]\ : SLE
      port map(D => \wptr_gray_1[12]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[12]_net_1\);
    
    \wptr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[6]_net_1\, S
         => \wptr_s[7]\, Y => OPEN, FCO => \wptr_cry[7]_net_1\);
    
    \wptr_bin_sync2[2]\ : SLE
      port map(D => \wptr_bin_sync[2]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[2]_net_1\);
    
    fulli_0_1 : CFG4
      generic map(INIT => x"01FF")

      port map(A => \wdiff_bus[6]\, B => \wdiff_bus[5]\, C => 
        N_12, D => \fulli_0_a3_3\, Y => \fulli_0_1\);
    
    \L1.un4_re_i_9\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \fifo_MEMRADDR[4]\, B => \fifo_MEMRADDR[3]\, 
        C => \fifo_MEMRADDR[0]\, D => un4_re_i_0, Y => un4_re_i_9);
    
    un1_memraddr_r_cry_3 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[3]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_2\, 
        S => un1_memraddr_r_cry_3_S_2, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_3\);
    
    \rptr_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \rptr[0]_net_1\, Y => \rptr_s[0]\);
    
    un1_memraddr_r_cry_1 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[1]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        un1_memraddr_r_s_1_929_FCO, S => un1_memraddr_r_cry_1_S_2, 
        Y => OPEN, FCO => \un1_memraddr_r_cry_1\);
    
    \rptr[4]\ : SLE
      port map(D => \rptr_s[4]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[4]_net_1\);
    
    \memwaddr_r_2[5]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_5_S_2, D => un4_we_i_9, Y => 
        \memwaddr_r_2[5]_net_1\);
    
    \wptr_gray[6]\ : SLE
      port map(D => \wptr_gray_1[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[6]_net_1\);
    
    \wptr_gray_1[3]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[3]_net_1\, B => \wptr[4]_net_1\, Y => 
        \wptr_gray_1[3]_net_1\);
    
    \wptr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[4]_net_1\, S
         => \wptr_s[5]\, Y => OPEN, FCO => \wptr_cry[5]_net_1\);
    
    un1_memraddr_r_cry_9 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[9]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_8\, 
        S => un1_memraddr_r_cry_9_S_2, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_9\);
    
    fulli_0_a3_0 : CFG4
      generic map(INIT => x"4000")

      port map(A => wdiff_bus_cry_0_Y_3, B => \wdiff_bus[1]\, C
         => \wdiff_bus[4]\, D => \fulli_0_a3_0_3\, Y => N_12);
    
    \rptr_gray[4]\ : SLE
      port map(D => \rptr_gray_1[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[4]_net_1\);
    
    un1_memraddr_r_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_4\, 
        S => un1_memraddr_r_cry_5_S_2, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_5\);
    
    \wptr_bin_sync2[4]\ : SLE
      port map(D => \wptr_bin_sync[4]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[4]_net_1\);
    
    \L1.empty_r_3_0_a2_6\ : CFG3
      generic map(INIT => x"0E")

      port map(A => iRX_FIFO_rd_en_0, B => rdiff_bus_cry_0_Y_3, C
         => \rdiff_bus[13]\, Y => empty_r_3_0_a2_6);
    
    \wptr[3]\ : SLE
      port map(D => \wptr_s[3]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[3]_net_1\);
    
    \L1.un4_we_i_9\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \fifo_MEMWADDR[4]\, B => \fifo_MEMWADDR[3]\, 
        C => \fifo_MEMWADDR[0]\, D => un4_we_i_0, Y => un4_we_i_9);
    
    \memwaddr_r[6]\ : SLE
      port map(D => un1_memwaddr_r_cry_6_S_2, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[6]\);
    
    \wptr[6]\ : SLE
      port map(D => \wptr_s[6]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[6]_net_1\);
    
    \memwaddr_r[9]\ : SLE
      port map(D => \memwaddr_r_2[9]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[9]\);
    
    un1_memraddr_r_s_1_929 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[0]\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => un1_memraddr_r_s_1_929_FCO);
    
    \memraddr_r[10]\ : SLE
      port map(D => \memraddr_r_2[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[10]\);
    
    \L1.un4_re_i_8\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \fifo_MEMRADDR[10]\, B => \fifo_MEMRADDR[9]\, 
        C => \fifo_MEMRADDR[8]\, D => \fifo_MEMRADDR[7]\, Y => 
        un4_re_i_8);
    
    \memwaddr_r[3]\ : SLE
      port map(D => un1_memwaddr_r_cry_3_S_2, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[3]\);
    
    \rptr_gray_1[12]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[13]_net_1\, B => \rptr[12]_net_1\, Y
         => \rptr_gray_1[12]_net_1\);
    
    wptr_s_903 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => wptr_s_903_FCO);
    
    full_r : SLE
      port map(D => fulli, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \iRX_FIFO_Full_0\);
    
    \rptr_bin_sync2[3]\ : SLE
      port map(D => \rptr_bin_sync[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[3]_net_1\);
    
    \wptr_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \wptr[0]_net_1\, Y => \wptr_s[0]\);
    
    \rptr[2]\ : SLE
      port map(D => \rptr_s[2]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[2]_net_1\);
    
    \memraddr_r[3]\ : SLE
      port map(D => un1_memraddr_r_cry_3_S_2, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[3]\);
    
    \wptr[13]\ : SLE
      port map(D => \wptr_s[13]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \wptr[13]_net_1\);
    
    \rptr_bin_sync2[9]\ : SLE
      port map(D => \rptr_bin_sync[9]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[9]_net_1\);
    
    \wptr_bin_sync2[13]\ : SLE
      port map(D => \wptr_bin_sync[13]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[13]_net_1\);
    
    \rptr[11]\ : SLE
      port map(D => \rptr_s[11]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rptr[11]_net_1\);
    
    \wptr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[5]_net_1\, S
         => \wptr_s[6]\, Y => OPEN, FCO => \wptr_cry[6]_net_1\);
    
    \rptr_bin_sync2[11]\ : SLE
      port map(D => \rptr_bin_sync[11]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[11]_net_1\);
    
    \wptr_bin_sync2[5]\ : SLE
      port map(D => \wptr_bin_sync[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[5]_net_1\);
    
    \L1.un4_we_i_8\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \fifo_MEMWADDR[10]\, B => \fifo_MEMWADDR[9]\, 
        C => \fifo_MEMWADDR[8]\, D => \fifo_MEMWADDR[7]\, Y => 
        un4_we_i_8);
    
    \wptr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[7]_net_1\, S
         => \wptr_s[8]\, Y => OPEN, FCO => \wptr_cry[8]_net_1\);
    
    \wptr_bin_sync2[1]\ : SLE
      port map(D => \wptr_bin_sync[1]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[1]_net_1\);
    
    Wr_corefifo_grayToBinConv : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_6
      port map(wptr_bin_sync(13) => \wptr_bin_sync[13]\, 
        wptr_bin_sync(12) => \wptr_bin_sync[12]\, 
        wptr_bin_sync(11) => \wptr_bin_sync[11]\, 
        wptr_bin_sync(10) => \wptr_bin_sync[10]\, 
        wptr_bin_sync(9) => \wptr_bin_sync[9]\, wptr_bin_sync(8)
         => \wptr_bin_sync[8]\, wptr_bin_sync(7) => 
        \wptr_bin_sync[7]\, wptr_bin_sync(6) => 
        \wptr_bin_sync[6]\, wptr_bin_sync(5) => 
        \wptr_bin_sync[5]\, wptr_bin_sync(4) => 
        \wptr_bin_sync[4]\, wptr_bin_sync(3) => 
        \wptr_bin_sync[3]\, wptr_bin_sync(2) => 
        \wptr_bin_sync[2]\, wptr_bin_sync(1) => 
        \wptr_bin_sync[1]\, wptr_bin_sync(0) => 
        \wptr_bin_sync[0]\, wptr_gray_sync(12) => 
        \wptr_gray_sync[12]\, wptr_gray_sync(11) => 
        \wptr_gray_sync[11]\, wptr_gray_sync(10) => 
        \wptr_gray_sync[10]\, wptr_gray_sync(9) => 
        \wptr_gray_sync[9]\, wptr_gray_sync(8) => 
        \wptr_gray_sync[8]\, wptr_gray_sync(7) => 
        \wptr_gray_sync[7]\, wptr_gray_sync(6) => 
        \wptr_gray_sync[6]\, wptr_gray_sync(5) => 
        \wptr_gray_sync[5]\, wptr_gray_sync(4) => 
        \wptr_gray_sync[4]\, wptr_gray_sync(3) => 
        \wptr_gray_sync[3]\, wptr_gray_sync(2) => 
        \wptr_gray_sync[2]\, wptr_gray_sync(1) => 
        \wptr_gray_sync[1]\, wptr_gray_sync(0) => 
        \wptr_gray_sync[0]\);
    
    \wptr_gray_1[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[4]_net_1\, B => \wptr[5]_net_1\, Y => 
        \wptr_gray_1[4]_net_1\);
    
    \rptr_bin_sync2[13]\ : SLE
      port map(D => \rptr_bin_sync[13]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[13]_net_1\);
    
    \L1.un4_re_i_7\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \fifo_MEMRADDR[12]\, B => \fifo_MEMRADDR[11]\, 
        C => \fifo_MEMRADDR[6]\, D => \fifo_MEMRADDR[5]\, Y => 
        un4_re_i_7);
    
    overflow_r : SLE
      port map(D => N_6_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        iRX_FIFO_OVERFLOW_0);
    
    fulli_0 : CFG4
      generic map(INIT => x"BAAA")

      port map(A => \wdiff_bus[13]\, B => \fulli_0_1\, C => 
        \wdiff_bus[11]\, D => \wdiff_bus[12]\, Y => fulli);
    
    \memraddr_r_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \fifo_MEMRADDR[0]\, Y => \fifo_MEMRADDR_i[0]\);
    
    \memraddr_r_2[8]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => 
        un1_memraddr_r_cry_8_S_2, D => un4_re_i_9, Y => 
        \memraddr_r_2[8]_net_1\);
    
    \rptr_gray[11]\ : SLE
      port map(D => \rptr_gray_1[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[11]_net_1\);
    
    \wptr_bin_sync2[10]\ : SLE
      port map(D => \wptr_bin_sync[10]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[10]_net_1\);
    
    \rptr[10]\ : SLE
      port map(D => \rptr_s[10]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rptr[10]_net_1\);
    
    \wptr[9]\ : SLE
      port map(D => \wptr_s[9]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[9]_net_1\);
    
    Wr_corefifo_doubleSync : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_3
      port map(wptr_gray(13) => \wptr_gray[13]_net_1\, 
        wptr_gray(12) => \wptr_gray[12]_net_1\, wptr_gray(11) => 
        \wptr_gray[11]_net_1\, wptr_gray(10) => 
        \wptr_gray[10]_net_1\, wptr_gray(9) => 
        \wptr_gray[9]_net_1\, wptr_gray(8) => 
        \wptr_gray[8]_net_1\, wptr_gray(7) => 
        \wptr_gray[7]_net_1\, wptr_gray(6) => 
        \wptr_gray[6]_net_1\, wptr_gray(5) => 
        \wptr_gray[5]_net_1\, wptr_gray(4) => 
        \wptr_gray[4]_net_1\, wptr_gray(3) => 
        \wptr_gray[3]_net_1\, wptr_gray(2) => 
        \wptr_gray[2]_net_1\, wptr_gray(1) => 
        \wptr_gray[1]_net_1\, wptr_gray(0) => 
        \wptr_gray[0]_net_1\, wptr_gray_sync(12) => 
        \wptr_gray_sync[12]\, wptr_gray_sync(11) => 
        \wptr_gray_sync[11]\, wptr_gray_sync(10) => 
        \wptr_gray_sync[10]\, wptr_gray_sync(9) => 
        \wptr_gray_sync[9]\, wptr_gray_sync(8) => 
        \wptr_gray_sync[8]\, wptr_gray_sync(7) => 
        \wptr_gray_sync[7]\, wptr_gray_sync(6) => 
        \wptr_gray_sync[6]\, wptr_gray_sync(5) => 
        \wptr_gray_sync[5]\, wptr_gray_sync(4) => 
        \wptr_gray_sync[4]\, wptr_gray_sync(3) => 
        \wptr_gray_sync[3]\, wptr_gray_sync(2) => 
        \wptr_gray_sync[2]\, wptr_gray_sync(1) => 
        \wptr_gray_sync[1]\, wptr_gray_sync(0) => 
        \wptr_gray_sync[0]\, wptr_bin_sync_0 => 
        \wptr_bin_sync[13]\, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, irx_fifo_rst_i => 
        irx_fifo_rst_i);
    
    un1_memwaddr_r_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_4\, 
        S => un1_memwaddr_r_cry_5_S_2, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_5\);
    
    \rptr_gray[0]\ : SLE
      port map(D => \rptr_gray_1[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[0]_net_1\);
    
    empty_r : SLE
      port map(D => empty_r_3, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \iRX_FIFO_Empty_0\);
    
    \memwaddr_r_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \fifo_MEMWADDR[0]\, Y => \fifo_MEMWADDR_i[0]\);
    
    \memwaddr_r_2[12]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_s_12_S_2, D => un4_we_i_9, Y => 
        \memwaddr_r_2[12]_net_1\);
    
    \rptr_gray_1[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[7]_net_1\, B => \rptr[8]_net_1\, Y => 
        \rptr_gray_1[7]_net_1\);
    
    un1_memraddr_r_cry_2 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[2]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_1\, 
        S => un1_memraddr_r_cry_2_S_2, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_2\);
    
    wdiff_bus_cry_12 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[12]_net_1\, B => 
        \rptr_bin_sync2[12]_net_1\, C => GND_net_1, D => 
        GND_net_1, FCI => \wdiff_bus_cry_11\, S => 
        \wdiff_bus[12]\, Y => OPEN, FCO => \wdiff_bus_cry_12\);
    
    \wptr[4]\ : SLE
      port map(D => \wptr_s[4]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[4]_net_1\);
    
    rptr_s_902 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => rptr_s_902_FCO);
    
    un1_memraddr_r_cry_8 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[8]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_7\, 
        S => un1_memraddr_r_cry_8_S_2, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_8\);
    
    \rptr_s[13]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[13]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[12]_net_1\, S
         => \rptr_s[13]_net_1\, Y => OPEN, FCO => OPEN);
    
    \memwaddr_r[8]\ : SLE
      port map(D => \memwaddr_r_2[8]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[8]\);
    
    \memwaddr_r[2]\ : SLE
      port map(D => un1_memwaddr_r_cry_2_S_2, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[2]\);
    
    \wptr_bin_sync2[11]\ : SLE
      port map(D => \wptr_bin_sync[11]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[11]_net_1\);
    
    \L1.un4_we_i_7\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \fifo_MEMWADDR[12]\, B => \fifo_MEMWADDR[11]\, 
        C => \fifo_MEMWADDR[6]\, D => \fifo_MEMWADDR[5]\, Y => 
        un4_we_i_7);
    
    \wptr_gray_1[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[1]_net_1\, B => \wptr[2]_net_1\, Y => 
        \wptr_gray_1[1]_net_1\);
    
    underflow_r : SLE
      port map(D => N_5_i, CLK => m2s010_som_sb_0_CCC_71MHz, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => iRX_FIFO_UNDERRUN_0);
    
    \memwaddr_r_2[11]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_11_S_2, D => un4_we_i_9, Y => 
        \memwaddr_r_2[11]_net_1\);
    
    \memraddr_r_2[12]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => 
        un1_memraddr_r_s_12_S_2, D => un4_re_i_9, Y => 
        \memraddr_r_2[12]_net_1\);
    
    \wptr_gray[5]\ : SLE
      port map(D => \wptr_gray_1[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[5]_net_1\);
    
    overflow_r_RNO : CFG3
      generic map(INIT => x"80")

      port map(A => RX_FIFO_TxColDetDis_wr_en, B => 
        \iRX_FIFO_Full_0\, C => iRX_FIFO_wr_en_0_0, Y => N_6_i);
    
    \memraddr_r[7]\ : SLE
      port map(D => \memraddr_r_2[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[7]\);
    
    un1_memraddr_r_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_5\, 
        S => un1_memraddr_r_cry_6_S_2, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_6\);
    
    \rptr_bin_sync2[10]\ : SLE
      port map(D => \rptr_bin_sync[10]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[10]_net_1\);
    
    wdiff_bus_s_13 : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \rptr_bin_sync2[13]_net_1\, C
         => \wptr[13]_net_1\, D => GND_net_1, FCI => 
        \wdiff_bus_cry_12\, S => \wdiff_bus[13]\, Y => OPEN, FCO
         => OPEN);
    
    wdiff_bus_cry_10 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[10]_net_1\, B => 
        \rptr_bin_sync2[10]_net_1\, C => GND_net_1, D => 
        GND_net_1, FCI => \wdiff_bus_cry_9\, S => \wdiff_bus[10]\, 
        Y => OPEN, FCO => \wdiff_bus_cry_10\);
    
    \memwaddr_r[11]\ : SLE
      port map(D => \memwaddr_r_2[11]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[11]\);
    
    \wptr_gray[8]\ : SLE
      port map(D => \wptr_gray_1[8]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[8]_net_1\);
    
    \memraddr_r_2[11]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => 
        un1_memraddr_r_cry_11_S_2, D => un4_re_i_9, Y => 
        \memraddr_r_2[11]_net_1\);
    
    un1_memraddr_r_s_12 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[12]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_11\, 
        S => un1_memraddr_r_s_12_S_2, Y => OPEN, FCO => OPEN);
    
    \wptr_gray[7]\ : SLE
      port map(D => \wptr_gray_1[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[7]_net_1\);
    
    \wptr_gray_1[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[5]_net_1\, B => \wptr[6]_net_1\, Y => 
        \wptr_gray_1[5]_net_1\);
    
    \memwaddr_r[5]\ : SLE
      port map(D => \memwaddr_r_2[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[5]\);
    
    \L1.empty_r_3_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => empty_r_3_0_a2_6, B => empty_r_3_0_a2_7, C
         => empty_r_3_0_a2_9, D => empty_r_3_0_a2_8, Y => 
        empty_r_3);
    
    un1_memraddr_r_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_3\, 
        S => un1_memraddr_r_cry_4_S_2, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_4\);
    
    \rptr[8]\ : SLE
      port map(D => \rptr_s[8]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[8]_net_1\);
    
    Rd_corefifo_doubleSync : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0_2
      port map(rptr_gray(13) => \rptr_gray[13]_net_1\, 
        rptr_gray(12) => \rptr_gray[12]_net_1\, rptr_gray(11) => 
        \rptr_gray[11]_net_1\, rptr_gray(10) => 
        \rptr_gray[10]_net_1\, rptr_gray(9) => 
        \rptr_gray[9]_net_1\, rptr_gray(8) => 
        \rptr_gray[8]_net_1\, rptr_gray(7) => 
        \rptr_gray[7]_net_1\, rptr_gray(6) => 
        \rptr_gray[6]_net_1\, rptr_gray(5) => 
        \rptr_gray[5]_net_1\, rptr_gray(4) => 
        \rptr_gray[4]_net_1\, rptr_gray(3) => 
        \rptr_gray[3]_net_1\, rptr_gray(2) => 
        \rptr_gray[2]_net_1\, rptr_gray(1) => 
        \rptr_gray[1]_net_1\, rptr_gray(0) => 
        \rptr_gray[0]_net_1\, rptr_gray_sync(12) => 
        \rptr_gray_sync[12]\, rptr_gray_sync(11) => 
        \rptr_gray_sync[11]\, rptr_gray_sync(10) => 
        \rptr_gray_sync[10]\, rptr_gray_sync(9) => 
        \rptr_gray_sync[9]\, rptr_gray_sync(8) => 
        \rptr_gray_sync[8]\, rptr_gray_sync(7) => 
        \rptr_gray_sync[7]\, rptr_gray_sync(6) => 
        \rptr_gray_sync[6]\, rptr_gray_sync(5) => 
        \rptr_gray_sync[5]\, rptr_gray_sync(4) => 
        \rptr_gray_sync[4]\, rptr_gray_sync(3) => 
        \rptr_gray_sync[3]\, rptr_gray_sync(2) => 
        \rptr_gray_sync[2]\, rptr_gray_sync(1) => 
        \rptr_gray_sync[1]\, rptr_gray_sync(0) => 
        \rptr_gray_sync[0]\, rptr_bin_sync_0 => 
        \rptr_bin_sync[13]\, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, irx_fifo_rst_i => irx_fifo_rst_i);
    
    underflow_r_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => iRX_FIFO_rd_en_0, B => \iRX_FIFO_Empty_0\, Y
         => N_5_i);
    
    \rptr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[3]_net_1\, S
         => \rptr_s[4]\, Y => OPEN, FCO => \rptr_cry[4]_net_1\);
    
    wdiff_bus_cry_2 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[2]_net_1\, B => 
        \rptr_bin_sync2[2]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_1\, S => \wdiff_bus[2]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_2\);
    
    \rptr_gray[2]\ : SLE
      port map(D => \rptr_gray_1[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[2]_net_1\);
    
    \wptr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[8]_net_1\, S
         => \wptr_s[9]\, Y => OPEN, FCO => \wptr_cry[9]_net_1\);
    
    \wptr_bin_sync2[3]\ : SLE
      port map(D => \wptr_bin_sync[3]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[3]_net_1\);
    
    \rptr[12]\ : SLE
      port map(D => \rptr_s[12]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rptr[12]_net_1\);
    
    \wptr[2]\ : SLE
      port map(D => \wptr_s[2]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[2]_net_1\);
    
    \rptr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[1]_net_1\, S
         => \rptr_s[2]\, Y => OPEN, FCO => \rptr_cry[2]_net_1\);
    
    rdiff_bus_cry_9 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[9]_net_1\, B => 
        \rptr[9]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_8\, S => \rdiff_bus[9]\, Y => OPEN, FCO
         => \rdiff_bus_cry_9\);
    
    \memwaddr_r[0]\ : SLE
      port map(D => \fifo_MEMWADDR_i[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[0]\);
    
    \wptr_gray[2]\ : SLE
      port map(D => \wptr_gray_1[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[2]_net_1\);
    
    \wptr_cry[12]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[12]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[11]_net_1\, S
         => \wptr_s[12]\, Y => OPEN, FCO => \wptr_cry[12]_net_1\);
    
    \memwaddr_r_2[7]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_7_S_2, D => un4_we_i_9, Y => 
        \memwaddr_r_2[7]_net_1\);
    
    wdiff_bus_cry_4 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[4]_net_1\, B => 
        \rptr_bin_sync2[4]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_3\, S => \wdiff_bus[4]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_4\);
    
    un1_memraddr_r_cry_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_6\, 
        S => un1_memraddr_r_cry_7_S_2, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_7\);
    
    \wptr_s[13]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[13]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[12]_net_1\, S
         => \wptr_s[13]_net_1\, Y => OPEN, FCO => OPEN);
    
    \wptr_gray[11]\ : SLE
      port map(D => \wptr_gray_1[11]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[11]_net_1\);
    
    \wptr_bin_sync2[9]\ : SLE
      port map(D => \wptr_bin_sync[9]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[9]_net_1\);
    
    \rptr_gray_1[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[6]_net_1\, B => \rptr[7]_net_1\, Y => 
        \rptr_gray_1[6]_net_1\);
    
    \wptr_gray_1[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[10]_net_1\, B => \wptr[11]_net_1\, Y
         => \wptr_gray_1[10]_net_1\);
    
    wdiff_bus_cry_6 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[6]_net_1\, B => 
        \rptr_bin_sync2[6]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_5\, S => \wdiff_bus[6]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_6\);
    
    \rptr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[2]_net_1\, S
         => \rptr_s[3]\, Y => OPEN, FCO => \rptr_cry[3]_net_1\);
    
    \memraddr_r[4]\ : SLE
      port map(D => un1_memraddr_r_cry_4_S_2, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[4]\);
    
    \rptr[13]\ : SLE
      port map(D => \rptr_s[13]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rptr[13]_net_1\);
    
    \wptr_cry[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[10]_net_1\, S
         => \wptr_s[11]\, Y => OPEN, FCO => \wptr_cry[11]_net_1\);
    
    \memwaddr_r_2[8]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_8_S_2, D => un4_we_i_9, Y => 
        \memwaddr_r_2[8]_net_1\);
    
    \memwaddr_r[12]\ : SLE
      port map(D => \memwaddr_r_2[12]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[12]\);
    
    \L1.un4_re_i_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => \fifo_MEMRADDR[1]\, B => \fifo_MEMRADDR[2]\, 
        Y => un4_re_i_0);
    
    \rptr_cry[12]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[12]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[11]_net_1\, S
         => \rptr_s[12]\, Y => OPEN, FCO => \rptr_cry[12]_net_1\);
    
    memre_0_a2 : CFG2
      generic map(INIT => x"2")

      port map(A => iRX_FIFO_rd_en_0, B => \iRX_FIFO_Empty_0\, Y
         => \fifo_MEMRE\);
    
    \memraddr_r[11]\ : SLE
      port map(D => \memraddr_r_2[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[11]\);
    
    rdiff_bus_cry_12 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[12]_net_1\, B => 
        \rptr[12]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_11\, S => \rdiff_bus[12]\, Y => OPEN, FCO
         => \rdiff_bus_cry_12\);
    
    \memraddr_r[5]\ : SLE
      port map(D => \memraddr_r_2[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[5]\);
    
    \rptr_gray[6]\ : SLE
      port map(D => \rptr_gray_1[6]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[6]_net_1\);
    
    \memraddr_r[9]\ : SLE
      port map(D => \memraddr_r_2[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[9]\);
    
    \rptr[0]\ : SLE
      port map(D => \rptr_s[0]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[0]_net_1\);
    
    \wptr[10]\ : SLE
      port map(D => \wptr_s[10]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[10]_net_1\);
    
    \L1.un4_we_i_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => \fifo_MEMWADDR[1]\, B => \fifo_MEMWADDR[2]\, 
        Y => un4_we_i_0);
    
    wdiff_bus_cry_1 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[1]_net_1\, B => 
        \rptr_bin_sync2[1]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_0\, S => \wdiff_bus[1]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_1\);
    
    rdiff_bus_cry_2 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[2]_net_1\, B => 
        \rptr[2]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_1\, S => \rdiff_bus[2]\, Y => OPEN, FCO
         => \rdiff_bus_cry_2\);
    
    \wptr_gray[9]\ : SLE
      port map(D => \wptr_gray_1[9]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[9]_net_1\);
    
    \rptr_gray_1[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[4]_net_1\, B => \rptr[5]_net_1\, Y => 
        \rptr_gray_1[4]_net_1\);
    
    \wptr_gray_1[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[8]_net_1\, B => \wptr[9]_net_1\, Y => 
        \wptr_gray_1[8]_net_1\);
    
    Rd_corefifo_grayToBinConv : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_5
      port map(rptr_bin_sync(13) => \rptr_bin_sync[13]\, 
        rptr_bin_sync(12) => \rptr_bin_sync[12]\, 
        rptr_bin_sync(11) => \rptr_bin_sync[11]\, 
        rptr_bin_sync(10) => \rptr_bin_sync[10]\, 
        rptr_bin_sync(9) => \rptr_bin_sync[9]\, rptr_bin_sync(8)
         => \rptr_bin_sync[8]\, rptr_bin_sync(7) => 
        \rptr_bin_sync[7]\, rptr_bin_sync(6) => nc2, 
        rptr_bin_sync(5) => \rptr_bin_sync[5]\, rptr_bin_sync(4)
         => nc1, rptr_bin_sync(3) => \rptr_bin_sync[3]\, 
        rptr_bin_sync(2) => \rptr_bin_sync[2]\, rptr_bin_sync(1)
         => \rptr_bin_sync[1]\, rptr_bin_sync(0) => 
        \rptr_bin_sync[0]\, rptr_gray_sync(12) => 
        \rptr_gray_sync[12]\, rptr_gray_sync(11) => 
        \rptr_gray_sync[11]\, rptr_gray_sync(10) => 
        \rptr_gray_sync[10]\, rptr_gray_sync(9) => 
        \rptr_gray_sync[9]\, rptr_gray_sync(8) => 
        \rptr_gray_sync[8]\, rptr_gray_sync(7) => 
        \rptr_gray_sync[7]\, rptr_gray_sync(6) => 
        \rptr_gray_sync[6]\, rptr_gray_sync(5) => 
        \rptr_gray_sync[5]\, rptr_gray_sync(4) => 
        \rptr_gray_sync[4]\, rptr_gray_sync(3) => 
        \rptr_gray_sync[3]\, rptr_gray_sync(2) => 
        \rptr_gray_sync[2]\, rptr_gray_sync(1) => 
        \rptr_gray_sync[1]\, rptr_gray_sync(0) => 
        \rptr_gray_sync[0]\, bin_N_6_i => bin_N_6_i, bin_N_4_0_i
         => bin_N_4_0_i);
    
    \rptr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => rptr_s_902_FCO, S => 
        \rptr_s[1]\, Y => OPEN, FCO => \rptr_cry[1]_net_1\);
    
    \rptr_cry[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[10]_net_1\, S
         => \rptr_s[11]\, Y => OPEN, FCO => \rptr_cry[11]_net_1\);
    
    rdiff_bus_cry_3 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[3]_net_1\, B => 
        \rptr[3]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_2\, S => \rdiff_bus[3]\, Y => OPEN, FCO
         => \rdiff_bus_cry_3\);
    
    rdiff_bus_cry_10 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[10]_net_1\, B => 
        \rptr[10]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_9\, S => \rdiff_bus[10]\, Y => OPEN, FCO
         => \rdiff_bus_cry_10\);
    
    un1_memwaddr_r_cry_11 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[11]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_10\, 
        S => un1_memwaddr_r_cry_11_S_2, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_11\);
    
    \memraddr_r[6]\ : SLE
      port map(D => un1_memraddr_r_cry_6_S_2, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[6]\);
    
    \rptr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[6]_net_1\, S
         => \rptr_s[7]\, Y => OPEN, FCO => \rptr_cry[7]_net_1\);
    
    rdiff_bus_cry_0 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => rdiff_bus, B => \rptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => rdiff_bus_cry_0_Y_3, FCO => \rdiff_bus_cry_0\);
    
    \memraddr_r[2]\ : SLE
      port map(D => un1_memraddr_r_cry_2_S_2, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[2]\);
    
    \wptr[8]\ : SLE
      port map(D => \wptr_s[8]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[8]_net_1\);
    
    wdiff_bus_cry_3 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[3]_net_1\, B => 
        \rptr_bin_sync2[3]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_2\, S => \wdiff_bus[3]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_3\);
    
    rdiff_bus_s_13 : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \rptr[13]_net_1\, C => 
        \wptr_bin_sync2[13]_net_1\, D => GND_net_1, FCI => 
        \rdiff_bus_cry_12\, S => \rdiff_bus[13]\, Y => OPEN, FCO
         => OPEN);
    
    \memraddr_r[12]\ : SLE
      port map(D => \memraddr_r_2[12]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[12]\);
    
    \wptr_gray_1[11]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[11]_net_1\, B => \wptr[12]_net_1\, Y
         => \wptr_gray_1[11]_net_1\);
    
    \rptr_gray[7]\ : SLE
      port map(D => \rptr_gray_1[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[7]_net_1\);
    
    \wptr_gray[0]\ : SLE
      port map(D => \wptr_gray_1[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[0]_net_1\);
    
    \rptr_gray_1[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[0]_net_1\, B => \rptr[1]_net_1\, Y => 
        \rptr_gray_1[0]_net_1\);
    
    un1_memwaddr_r_cry_10 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_9\, 
        S => un1_memwaddr_r_cry_10_S_2, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_10\);
    
    \rptr_gray_1[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[8]_net_1\, B => \rptr[9]_net_1\, Y => 
        \rptr_gray_1[8]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_2 is

    port( RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          RX_FIFO_DOUT_3            : out   std_logic_vector(8 downto 0);
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_wr_en_0_0        : in    std_logic;
          iRX_FIFO_rd_en_0          : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          RX_FIFO_TxColDetDis_wr_en : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          irx_fifo_rst_i            : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_2;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_2 is 

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_2
    port( fifo_MEMRADDR             : in    std_logic_vector(12 downto 0) := (others => 'U');
          fifo_MEMWADDR             : in    std_logic_vector(12 downto 0) := (others => 'U');
          RDATA_int                 : out   std_logic_vector(8 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          fifo_MEMRE                : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          fifo_MEMWE                : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_2
    port( fifo_MEMRADDR             : out   std_logic_vector(12 downto 0);
          fifo_MEMWADDR             : out   std_logic_vector(12 downto 0);
          iRX_FIFO_wr_en_0_0        : in    std_logic := 'U';
          iRX_FIFO_rd_en_0          : in    std_logic := 'U';
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          RX_FIFO_TxColDetDis_wr_en : in    std_logic := 'U';
          fifo_MEMRE                : out   std_logic;
          fifo_MEMWE                : out   std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          irx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \RDATA_r[0]_net_1\, VCC_net_1, \RDATA_int[0]\, 
        un6_fifo_memre_2, GND_net_1, \RDATA_r[1]_net_1\, 
        \RDATA_int[1]\, \RDATA_r[2]_net_1\, \RDATA_int[2]\, 
        \RDATA_r[3]_net_1\, \RDATA_int[3]\, \RDATA_r[4]_net_1\, 
        \RDATA_int[4]\, \RDATA_r[5]_net_1\, \RDATA_int[5]\, 
        \RDATA_r[6]_net_1\, \RDATA_int[6]\, \RDATA_r[7]_net_1\, 
        \RDATA_int[7]\, \RDATA_r[8]_net_1\, \RDATA_int[8]\, 
        \re_set\, \REN_d1\, un9_fifo_memre_2, fifo_MEMRE, \RE_d1\, 
        \re_pulse_d1\, \re_pulse\, \fifo_MEMRADDR[0]\, 
        \fifo_MEMRADDR[1]\, \fifo_MEMRADDR[2]\, 
        \fifo_MEMRADDR[3]\, \fifo_MEMRADDR[4]\, 
        \fifo_MEMRADDR[5]\, \fifo_MEMRADDR[6]\, 
        \fifo_MEMRADDR[7]\, \fifo_MEMRADDR[8]\, 
        \fifo_MEMRADDR[9]\, \fifo_MEMRADDR[10]\, 
        \fifo_MEMRADDR[11]\, \fifo_MEMRADDR[12]\, 
        \fifo_MEMWADDR[0]\, \fifo_MEMWADDR[1]\, 
        \fifo_MEMWADDR[2]\, \fifo_MEMWADDR[3]\, 
        \fifo_MEMWADDR[4]\, \fifo_MEMWADDR[5]\, 
        \fifo_MEMWADDR[6]\, \fifo_MEMWADDR[7]\, 
        \fifo_MEMWADDR[8]\, \fifo_MEMWADDR[9]\, 
        \fifo_MEMWADDR[10]\, \fifo_MEMWADDR[11]\, 
        \fifo_MEMWADDR[12]\, fifo_MEMWE : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_2
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_2(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_2
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_2(DEF_ARCH);
begin 


    re_pulse : CFG3
      generic map(INIT => x"DC")

      port map(A => fifo_MEMRE, B => \re_set\, C => \REN_d1\, Y
         => \re_pulse\);
    
    \RDATA_r[3]\ : SLE
      port map(D => \RDATA_int[3]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un6_fifo_memre_2, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[3]_net_1\);
    
    \Q[6]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[6]_net_1\, C => 
        \RDATA_int[6]\, D => \RE_d1\, Y => RX_FIFO_DOUT_3(6));
    
    re_pulse_d1 : SLE
      port map(D => \re_pulse\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \re_pulse_d1\);
    
    \RDATA_r[5]\ : SLE
      port map(D => \RDATA_int[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un6_fifo_memre_2, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[5]_net_1\);
    
    un9_fifo_memre : CFG2
      generic map(INIT => x"6")

      port map(A => fifo_MEMRE, B => \REN_d1\, Y => 
        un9_fifo_memre_2);
    
    \RDATA_r[8]\ : SLE
      port map(D => \RDATA_int[8]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un6_fifo_memre_2, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[8]_net_1\);
    
    \Q[2]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[2]_net_1\, C => 
        \RDATA_int[2]\, D => \RE_d1\, Y => RX_FIFO_DOUT_3(2));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \RW1.UI_ram_wrapper_1\ : FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper_2
      port map(fifo_MEMRADDR(12) => \fifo_MEMRADDR[12]\, 
        fifo_MEMRADDR(11) => \fifo_MEMRADDR[11]\, 
        fifo_MEMRADDR(10) => \fifo_MEMRADDR[10]\, 
        fifo_MEMRADDR(9) => \fifo_MEMRADDR[9]\, fifo_MEMRADDR(8)
         => \fifo_MEMRADDR[8]\, fifo_MEMRADDR(7) => 
        \fifo_MEMRADDR[7]\, fifo_MEMRADDR(6) => 
        \fifo_MEMRADDR[6]\, fifo_MEMRADDR(5) => 
        \fifo_MEMRADDR[5]\, fifo_MEMRADDR(4) => 
        \fifo_MEMRADDR[4]\, fifo_MEMRADDR(3) => 
        \fifo_MEMRADDR[3]\, fifo_MEMRADDR(2) => 
        \fifo_MEMRADDR[2]\, fifo_MEMRADDR(1) => 
        \fifo_MEMRADDR[1]\, fifo_MEMRADDR(0) => 
        \fifo_MEMRADDR[0]\, fifo_MEMWADDR(12) => 
        \fifo_MEMWADDR[12]\, fifo_MEMWADDR(11) => 
        \fifo_MEMWADDR[11]\, fifo_MEMWADDR(10) => 
        \fifo_MEMWADDR[10]\, fifo_MEMWADDR(9) => 
        \fifo_MEMWADDR[9]\, fifo_MEMWADDR(8) => 
        \fifo_MEMWADDR[8]\, fifo_MEMWADDR(7) => 
        \fifo_MEMWADDR[7]\, fifo_MEMWADDR(6) => 
        \fifo_MEMWADDR[6]\, fifo_MEMWADDR(5) => 
        \fifo_MEMWADDR[5]\, fifo_MEMWADDR(4) => 
        \fifo_MEMWADDR[4]\, fifo_MEMWADDR(3) => 
        \fifo_MEMWADDR[3]\, fifo_MEMWADDR(2) => 
        \fifo_MEMWADDR[2]\, fifo_MEMWADDR(1) => 
        \fifo_MEMWADDR[1]\, fifo_MEMWADDR(0) => 
        \fifo_MEMWADDR[0]\, RDATA_int(8) => \RDATA_int[8]\, 
        RDATA_int(7) => \RDATA_int[7]\, RDATA_int(6) => 
        \RDATA_int[6]\, RDATA_int(5) => \RDATA_int[5]\, 
        RDATA_int(4) => \RDATA_int[4]\, RDATA_int(3) => 
        \RDATA_int[3]\, RDATA_int(2) => \RDATA_int[2]\, 
        RDATA_int(1) => \RDATA_int[1]\, RDATA_int(0) => 
        \RDATA_int[0]\, RX_FIFO_DIN_pipe(8) => 
        RX_FIFO_DIN_pipe(8), RX_FIFO_DIN_pipe(7) => 
        RX_FIFO_DIN_pipe(7), RX_FIFO_DIN_pipe(6) => 
        RX_FIFO_DIN_pipe(6), RX_FIFO_DIN_pipe(5) => 
        RX_FIFO_DIN_pipe(5), RX_FIFO_DIN_pipe(4) => 
        RX_FIFO_DIN_pipe(4), RX_FIFO_DIN_pipe(3) => 
        RX_FIFO_DIN_pipe(3), RX_FIFO_DIN_pipe(2) => 
        RX_FIFO_DIN_pipe(2), RX_FIFO_DIN_pipe(1) => 
        RX_FIFO_DIN_pipe(1), RX_FIFO_DIN_pipe(0) => 
        RX_FIFO_DIN_pipe(0), m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, fifo_MEMRE => fifo_MEMRE, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, fifo_MEMWE
         => fifo_MEMWE);
    
    \RDATA_r[0]\ : SLE
      port map(D => \RDATA_int[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un6_fifo_memre_2, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[0]_net_1\);
    
    \Q[4]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[4]_net_1\, C => 
        \RDATA_int[4]\, D => \RE_d1\, Y => RX_FIFO_DOUT_3(4));
    
    \RDATA_r[2]\ : SLE
      port map(D => \RDATA_int[2]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un6_fifo_memre_2, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[2]_net_1\);
    
    \RDATA_r[6]\ : SLE
      port map(D => \RDATA_int[6]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un6_fifo_memre_2, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[6]_net_1\);
    
    \L31.U_corefifo_async\ : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3_2
      port map(fifo_MEMRADDR(12) => \fifo_MEMRADDR[12]\, 
        fifo_MEMRADDR(11) => \fifo_MEMRADDR[11]\, 
        fifo_MEMRADDR(10) => \fifo_MEMRADDR[10]\, 
        fifo_MEMRADDR(9) => \fifo_MEMRADDR[9]\, fifo_MEMRADDR(8)
         => \fifo_MEMRADDR[8]\, fifo_MEMRADDR(7) => 
        \fifo_MEMRADDR[7]\, fifo_MEMRADDR(6) => 
        \fifo_MEMRADDR[6]\, fifo_MEMRADDR(5) => 
        \fifo_MEMRADDR[5]\, fifo_MEMRADDR(4) => 
        \fifo_MEMRADDR[4]\, fifo_MEMRADDR(3) => 
        \fifo_MEMRADDR[3]\, fifo_MEMRADDR(2) => 
        \fifo_MEMRADDR[2]\, fifo_MEMRADDR(1) => 
        \fifo_MEMRADDR[1]\, fifo_MEMRADDR(0) => 
        \fifo_MEMRADDR[0]\, fifo_MEMWADDR(12) => 
        \fifo_MEMWADDR[12]\, fifo_MEMWADDR(11) => 
        \fifo_MEMWADDR[11]\, fifo_MEMWADDR(10) => 
        \fifo_MEMWADDR[10]\, fifo_MEMWADDR(9) => 
        \fifo_MEMWADDR[9]\, fifo_MEMWADDR(8) => 
        \fifo_MEMWADDR[8]\, fifo_MEMWADDR(7) => 
        \fifo_MEMWADDR[7]\, fifo_MEMWADDR(6) => 
        \fifo_MEMWADDR[6]\, fifo_MEMWADDR(5) => 
        \fifo_MEMWADDR[5]\, fifo_MEMWADDR(4) => 
        \fifo_MEMWADDR[4]\, fifo_MEMWADDR(3) => 
        \fifo_MEMWADDR[3]\, fifo_MEMWADDR(2) => 
        \fifo_MEMWADDR[2]\, fifo_MEMWADDR(1) => 
        \fifo_MEMWADDR[1]\, fifo_MEMWADDR(0) => 
        \fifo_MEMWADDR[0]\, iRX_FIFO_wr_en_0_0 => 
        iRX_FIFO_wr_en_0_0, iRX_FIFO_rd_en_0 => iRX_FIFO_rd_en_0, 
        iRX_FIFO_Empty_0 => iRX_FIFO_Empty_0, iRX_FIFO_UNDERRUN_0
         => iRX_FIFO_UNDERRUN_0, iRX_FIFO_OVERFLOW_0 => 
        iRX_FIFO_OVERFLOW_0, iRX_FIFO_Full_0 => iRX_FIFO_Full_0, 
        RX_FIFO_TxColDetDis_wr_en => RX_FIFO_TxColDetDis_wr_en, 
        fifo_MEMRE => fifo_MEMRE, fifo_MEMWE => fifo_MEMWE, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz, 
        irx_fifo_rst_i => irx_fifo_rst_i);
    
    re_set : SLE
      port map(D => \REN_d1\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => un9_fifo_memre_2, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \re_set\);
    
    \Q[3]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[3]_net_1\, C => 
        \RDATA_int[3]\, D => \RE_d1\, Y => RX_FIFO_DOUT_3(3));
    
    \Q[7]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[7]_net_1\, C => 
        \RDATA_int[7]\, D => \RE_d1\, Y => RX_FIFO_DOUT_3(7));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \Q[8]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[8]_net_1\, C => 
        \RDATA_int[8]\, D => \RE_d1\, Y => RX_FIFO_DOUT_3(8));
    
    RE_d1 : SLE
      port map(D => iRX_FIFO_rd_en_0, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RE_d1\);
    
    \RDATA_r[7]\ : SLE
      port map(D => \RDATA_int[7]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un6_fifo_memre_2, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[7]_net_1\);
    
    \RDATA_r[4]\ : SLE
      port map(D => \RDATA_int[4]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un6_fifo_memre_2, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[4]_net_1\);
    
    \Q[1]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[1]_net_1\, C => 
        \RDATA_int[1]\, D => \RE_d1\, Y => RX_FIFO_DOUT_3(1));
    
    \Q[0]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[0]_net_1\, C => 
        \RDATA_int[0]\, D => \RE_d1\, Y => RX_FIFO_DOUT_3(0));
    
    REN_d1 : SLE
      port map(D => fifo_MEMRE, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \REN_d1\);
    
    \Q[5]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[5]_net_1\, C => 
        \RDATA_int[5]\, D => \RE_d1\, Y => RX_FIFO_DOUT_3(5));
    
    un6_fifo_memre : CFG2
      generic map(INIT => x"4")

      port map(A => fifo_MEMRE, B => \REN_d1\, Y => 
        un6_fifo_memre_2);
    
    \RDATA_r[1]\ : SLE
      port map(D => \RDATA_int[1]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un6_fifo_memre_2, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[1]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_2 is

    port( RX_FIFO_DOUT_3            : out   std_logic_vector(8 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          iRX_FIFO_rd_en_0          : in    std_logic;
          iRX_FIFO_wr_en_0_0        : in    std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          irx_fifo_rst_i            : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          RX_FIFO_TxColDetDis_wr_en : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic
        );

end FIFO_8Kx9_2;

architecture DEF_ARCH of FIFO_8Kx9_2 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_2
    port( RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          RX_FIFO_DOUT_3            : out   std_logic_vector(8 downto 0);
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_wr_en_0_0        : in    std_logic := 'U';
          iRX_FIFO_rd_en_0          : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          RX_FIFO_TxColDetDis_wr_en : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          irx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_2
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_2(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    FIFO_8Kx9_0 : FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO_2
      port map(RX_FIFO_DIN_pipe(8) => RX_FIFO_DIN_pipe(8), 
        RX_FIFO_DIN_pipe(7) => RX_FIFO_DIN_pipe(7), 
        RX_FIFO_DIN_pipe(6) => RX_FIFO_DIN_pipe(6), 
        RX_FIFO_DIN_pipe(5) => RX_FIFO_DIN_pipe(5), 
        RX_FIFO_DIN_pipe(4) => RX_FIFO_DIN_pipe(4), 
        RX_FIFO_DIN_pipe(3) => RX_FIFO_DIN_pipe(3), 
        RX_FIFO_DIN_pipe(2) => RX_FIFO_DIN_pipe(2), 
        RX_FIFO_DIN_pipe(1) => RX_FIFO_DIN_pipe(1), 
        RX_FIFO_DIN_pipe(0) => RX_FIFO_DIN_pipe(0), 
        RX_FIFO_DOUT_3(8) => RX_FIFO_DOUT_3(8), RX_FIFO_DOUT_3(7)
         => RX_FIFO_DOUT_3(7), RX_FIFO_DOUT_3(6) => 
        RX_FIFO_DOUT_3(6), RX_FIFO_DOUT_3(5) => RX_FIFO_DOUT_3(5), 
        RX_FIFO_DOUT_3(4) => RX_FIFO_DOUT_3(4), RX_FIFO_DOUT_3(3)
         => RX_FIFO_DOUT_3(3), RX_FIFO_DOUT_3(2) => 
        RX_FIFO_DOUT_3(2), RX_FIFO_DOUT_3(1) => RX_FIFO_DOUT_3(1), 
        RX_FIFO_DOUT_3(0) => RX_FIFO_DOUT_3(0), iRX_FIFO_Full_0
         => iRX_FIFO_Full_0, iRX_FIFO_OVERFLOW_0 => 
        iRX_FIFO_OVERFLOW_0, iRX_FIFO_UNDERRUN_0 => 
        iRX_FIFO_UNDERRUN_0, iRX_FIFO_Empty_0 => iRX_FIFO_Empty_0, 
        iRX_FIFO_wr_en_0_0 => iRX_FIFO_wr_en_0_0, 
        iRX_FIFO_rd_en_0 => iRX_FIFO_rd_en_0, CommsFPGA_CCC_0_GL0
         => CommsFPGA_CCC_0_GL0, RX_FIFO_TxColDetDis_wr_en => 
        RX_FIFO_TxColDetDis_wr_en, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, irx_fifo_rst_i => 
        irx_fifo_rst_i);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top is

    port( RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          RDATA_int                 : out   std_logic_vector(8 downto 0);
          fifo_MEMWADDR             : in    std_logic_vector(12 downto 0);
          fifo_MEMRADDR             : in    std_logic_vector(12 downto 0);
          fifo_MEMWE                : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          fifo_MEMRE                : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component RAM1K18
    generic (MEMORYFILE:string := "");

    port( A_DOUT        : out   std_logic_vector(17 downto 0);
          B_DOUT        : out   std_logic_vector(17 downto 0);
          BUSY          : out   std_logic;
          A_CLK         : in    std_logic := 'U';
          A_DOUT_CLK    : in    std_logic := 'U';
          A_ARST_N      : in    std_logic := 'U';
          A_DOUT_EN     : in    std_logic := 'U';
          A_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_DOUT_ARST_N : in    std_logic := 'U';
          A_DOUT_SRST_N : in    std_logic := 'U';
          A_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          A_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          A_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          B_CLK         : in    std_logic := 'U';
          B_DOUT_CLK    : in    std_logic := 'U';
          B_ARST_N      : in    std_logic := 'U';
          B_DOUT_EN     : in    std_logic := 'U';
          B_BLK         : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_DOUT_ARST_N : in    std_logic := 'U';
          B_DOUT_SRST_N : in    std_logic := 'U';
          B_DIN         : in    std_logic_vector(17 downto 0) := (others => 'U');
          B_ADDR        : in    std_logic_vector(13 downto 0) := (others => 'U');
          B_WEN         : in    std_logic_vector(1 downto 0) := (others => 'U');
          A_EN          : in    std_logic := 'U';
          A_DOUT_LAT    : in    std_logic := 'U';
          A_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          A_WMODE       : in    std_logic := 'U';
          B_EN          : in    std_logic := 'U';
          B_DOUT_LAT    : in    std_logic := 'U';
          B_WIDTH       : in    std_logic_vector(2 downto 0) := (others => 'U');
          B_WMODE       : in    std_logic := 'U';
          SII_LOCK      : in    std_logic := 'U'
        );
  end component;

    signal VCC_net_1, GND_net_1 : std_logic;
    signal nc151, nc23, nc58, nc116, nc74, nc133, nc167, nc84, 
        nc39, nc72, nc82, nc145, nc160, nc57, nc156, nc125, nc73, 
        nc107, nc66, nc83, nc9, nc171, nc54, nc135, nc41, nc100, 
        nc52, nc29, nc118, nc60, nc141, nc45, nc53, nc121, nc158, 
        nc162, nc11, nc131, nc96, nc79, nc146, nc89, nc119, nc48, 
        nc126, nc15, nc102, nc3, nc47, nc90, nc159, nc136, nc59, 
        nc18, nc44, nc117, nc164, nc148, nc42, nc17, nc2, nc110, 
        nc128, nc43, nc157, nc36, nc61, nc104, nc138, nc14, nc150, 
        nc149, nc12, nc30, nc65, nc7, nc129, nc8, nc13, nc26, 
        nc139, nc163, nc112, nc68, nc49, nc170, nc91, nc5, nc20, 
        nc147, nc67, nc152, nc127, nc103, nc76, nc140, nc86, nc95, 
        nc120, nc165, nc137, nc64, nc19, nc70, nc62, nc80, nc130, 
        nc98, nc114, nc56, nc105, nc63, nc97, nc161, nc31, nc154, 
        nc50, nc142, nc94, nc122, nc35, nc4, nc92, nc101, nc166, 
        nc132, nc21, nc93, nc69, nc38, nc113, nc106, nc25, nc1, 
        nc37, nc144, nc153, nc46, nc71, nc124, nc81, nc168, nc34, 
        nc28, nc115, nc134, nc32, nc40, nc99, nc75, nc85, nc27, 
        nc108, nc16, nc155, nc51, nc33, nc169, nc78, nc24, nc88, 
        nc111, nc55, nc10, nc22, nc143, nc77, nc6, nc109, nc87, 
        nc123 : std_logic;

begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C2 : RAM1K18
      port map(A_DOUT(17) => nc151, A_DOUT(16) => nc23, 
        A_DOUT(15) => nc58, A_DOUT(14) => nc116, A_DOUT(13) => 
        nc74, A_DOUT(12) => nc133, A_DOUT(11) => nc167, 
        A_DOUT(10) => nc84, A_DOUT(9) => nc39, A_DOUT(8) => nc72, 
        A_DOUT(7) => nc82, A_DOUT(6) => nc145, A_DOUT(5) => nc160, 
        A_DOUT(4) => nc57, A_DOUT(3) => nc156, A_DOUT(2) => nc125, 
        A_DOUT(1) => RDATA_int(5), A_DOUT(0) => RDATA_int(4), 
        B_DOUT(17) => nc73, B_DOUT(16) => nc107, B_DOUT(15) => 
        nc66, B_DOUT(14) => nc83, B_DOUT(13) => nc9, B_DOUT(12)
         => nc171, B_DOUT(11) => nc54, B_DOUT(10) => nc135, 
        B_DOUT(9) => nc41, B_DOUT(8) => nc100, B_DOUT(7) => nc52, 
        B_DOUT(6) => nc29, B_DOUT(5) => nc118, B_DOUT(4) => nc60, 
        B_DOUT(3) => nc141, B_DOUT(2) => nc45, B_DOUT(1) => nc53, 
        B_DOUT(0) => nc121, BUSY => OPEN, A_CLK => 
        m2s010_som_sb_0_CCC_71MHz, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => fifo_MEMRE, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => fifo_MEMRADDR(12), A_ADDR(12) => fifo_MEMRADDR(11), 
        A_ADDR(11) => fifo_MEMRADDR(10), A_ADDR(10) => 
        fifo_MEMRADDR(9), A_ADDR(9) => fifo_MEMRADDR(8), 
        A_ADDR(8) => fifo_MEMRADDR(7), A_ADDR(7) => 
        fifo_MEMRADDR(6), A_ADDR(6) => fifo_MEMRADDR(5), 
        A_ADDR(5) => fifo_MEMRADDR(4), A_ADDR(4) => 
        fifo_MEMRADDR(3), A_ADDR(3) => fifo_MEMRADDR(2), 
        A_ADDR(2) => fifo_MEMRADDR(1), A_ADDR(1) => 
        fifo_MEMRADDR(0), A_ADDR(0) => GND_net_1, A_WEN(1) => 
        GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => GND_net_1, B_DIN(2) => GND_net_1, B_DIN(1)
         => RX_FIFO_DIN_pipe(5), B_DIN(0) => RX_FIFO_DIN_pipe(4), 
        B_ADDR(13) => fifo_MEMWADDR(12), B_ADDR(12) => 
        fifo_MEMWADDR(11), B_ADDR(11) => fifo_MEMWADDR(10), 
        B_ADDR(10) => fifo_MEMWADDR(9), B_ADDR(9) => 
        fifo_MEMWADDR(8), B_ADDR(8) => fifo_MEMWADDR(7), 
        B_ADDR(7) => fifo_MEMWADDR(6), B_ADDR(6) => 
        fifo_MEMWADDR(5), B_ADDR(5) => fifo_MEMWADDR(4), 
        B_ADDR(4) => fifo_MEMWADDR(3), B_ADDR(3) => 
        fifo_MEMWADDR(2), B_ADDR(2) => fifo_MEMWADDR(1), 
        B_ADDR(1) => fifo_MEMWADDR(0), B_ADDR(0) => GND_net_1, 
        B_WEN(1) => GND_net_1, B_WEN(0) => VCC_net_1, A_EN => 
        VCC_net_1, A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => 
        GND_net_1, A_WIDTH(1) => GND_net_1, A_WIDTH(0) => 
        VCC_net_1, A_WMODE => GND_net_1, B_EN => VCC_net_1, 
        B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => GND_net_1, 
        B_WIDTH(1) => GND_net_1, B_WIDTH(0) => VCC_net_1, B_WMODE
         => GND_net_1, SII_LOCK => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C1 : RAM1K18
      port map(A_DOUT(17) => nc158, A_DOUT(16) => nc162, 
        A_DOUT(15) => nc11, A_DOUT(14) => nc131, A_DOUT(13) => 
        nc96, A_DOUT(12) => nc79, A_DOUT(11) => nc146, A_DOUT(10)
         => nc89, A_DOUT(9) => nc119, A_DOUT(8) => nc48, 
        A_DOUT(7) => nc126, A_DOUT(6) => nc15, A_DOUT(5) => nc102, 
        A_DOUT(4) => nc3, A_DOUT(3) => nc47, A_DOUT(2) => nc90, 
        A_DOUT(1) => RDATA_int(3), A_DOUT(0) => RDATA_int(2), 
        B_DOUT(17) => nc159, B_DOUT(16) => nc136, B_DOUT(15) => 
        nc59, B_DOUT(14) => nc18, B_DOUT(13) => nc44, B_DOUT(12)
         => nc117, B_DOUT(11) => nc164, B_DOUT(10) => nc148, 
        B_DOUT(9) => nc42, B_DOUT(8) => nc17, B_DOUT(7) => nc2, 
        B_DOUT(6) => nc110, B_DOUT(5) => nc128, B_DOUT(4) => nc43, 
        B_DOUT(3) => nc157, B_DOUT(2) => nc36, B_DOUT(1) => nc61, 
        B_DOUT(0) => nc104, BUSY => OPEN, A_CLK => 
        m2s010_som_sb_0_CCC_71MHz, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => fifo_MEMRE, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => fifo_MEMRADDR(12), A_ADDR(12) => fifo_MEMRADDR(11), 
        A_ADDR(11) => fifo_MEMRADDR(10), A_ADDR(10) => 
        fifo_MEMRADDR(9), A_ADDR(9) => fifo_MEMRADDR(8), 
        A_ADDR(8) => fifo_MEMRADDR(7), A_ADDR(7) => 
        fifo_MEMRADDR(6), A_ADDR(6) => fifo_MEMRADDR(5), 
        A_ADDR(5) => fifo_MEMRADDR(4), A_ADDR(4) => 
        fifo_MEMRADDR(3), A_ADDR(3) => fifo_MEMRADDR(2), 
        A_ADDR(2) => fifo_MEMRADDR(1), A_ADDR(1) => 
        fifo_MEMRADDR(0), A_ADDR(0) => GND_net_1, A_WEN(1) => 
        GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => GND_net_1, B_DIN(2) => GND_net_1, B_DIN(1)
         => RX_FIFO_DIN_pipe(3), B_DIN(0) => RX_FIFO_DIN_pipe(2), 
        B_ADDR(13) => fifo_MEMWADDR(12), B_ADDR(12) => 
        fifo_MEMWADDR(11), B_ADDR(11) => fifo_MEMWADDR(10), 
        B_ADDR(10) => fifo_MEMWADDR(9), B_ADDR(9) => 
        fifo_MEMWADDR(8), B_ADDR(8) => fifo_MEMWADDR(7), 
        B_ADDR(7) => fifo_MEMWADDR(6), B_ADDR(6) => 
        fifo_MEMWADDR(5), B_ADDR(5) => fifo_MEMWADDR(4), 
        B_ADDR(4) => fifo_MEMWADDR(3), B_ADDR(3) => 
        fifo_MEMWADDR(2), B_ADDR(2) => fifo_MEMWADDR(1), 
        B_ADDR(1) => fifo_MEMWADDR(0), B_ADDR(0) => GND_net_1, 
        B_WEN(1) => GND_net_1, B_WEN(0) => VCC_net_1, A_EN => 
        VCC_net_1, A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => 
        GND_net_1, A_WIDTH(1) => GND_net_1, A_WIDTH(0) => 
        VCC_net_1, A_WMODE => GND_net_1, B_EN => VCC_net_1, 
        B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => GND_net_1, 
        B_WIDTH(1) => GND_net_1, B_WIDTH(0) => VCC_net_1, B_WMODE
         => GND_net_1, SII_LOCK => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C4 : RAM1K18
      port map(A_DOUT(17) => nc138, A_DOUT(16) => nc14, 
        A_DOUT(15) => nc150, A_DOUT(14) => nc149, A_DOUT(13) => 
        nc12, A_DOUT(12) => nc30, A_DOUT(11) => nc65, A_DOUT(10)
         => nc7, A_DOUT(9) => nc129, A_DOUT(8) => nc8, A_DOUT(7)
         => nc13, A_DOUT(6) => nc26, A_DOUT(5) => nc139, 
        A_DOUT(4) => nc163, A_DOUT(3) => nc112, A_DOUT(2) => nc68, 
        A_DOUT(1) => nc49, A_DOUT(0) => RDATA_int(8), B_DOUT(17)
         => nc170, B_DOUT(16) => nc91, B_DOUT(15) => nc5, 
        B_DOUT(14) => nc20, B_DOUT(13) => nc147, B_DOUT(12) => 
        nc67, B_DOUT(11) => nc152, B_DOUT(10) => nc127, B_DOUT(9)
         => nc103, B_DOUT(8) => nc76, B_DOUT(7) => nc140, 
        B_DOUT(6) => nc86, B_DOUT(5) => nc95, B_DOUT(4) => nc120, 
        B_DOUT(3) => nc165, B_DOUT(2) => nc137, B_DOUT(1) => nc64, 
        B_DOUT(0) => nc19, BUSY => OPEN, A_CLK => 
        m2s010_som_sb_0_CCC_71MHz, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => fifo_MEMRE, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => fifo_MEMRADDR(12), A_ADDR(12) => fifo_MEMRADDR(11), 
        A_ADDR(11) => fifo_MEMRADDR(10), A_ADDR(10) => 
        fifo_MEMRADDR(9), A_ADDR(9) => fifo_MEMRADDR(8), 
        A_ADDR(8) => fifo_MEMRADDR(7), A_ADDR(7) => 
        fifo_MEMRADDR(6), A_ADDR(6) => fifo_MEMRADDR(5), 
        A_ADDR(5) => fifo_MEMRADDR(4), A_ADDR(4) => 
        fifo_MEMRADDR(3), A_ADDR(3) => fifo_MEMRADDR(2), 
        A_ADDR(2) => fifo_MEMRADDR(1), A_ADDR(1) => 
        fifo_MEMRADDR(0), A_ADDR(0) => GND_net_1, A_WEN(1) => 
        GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => GND_net_1, B_DIN(2) => GND_net_1, B_DIN(1)
         => GND_net_1, B_DIN(0) => RX_FIFO_DIN_pipe(8), 
        B_ADDR(13) => fifo_MEMWADDR(12), B_ADDR(12) => 
        fifo_MEMWADDR(11), B_ADDR(11) => fifo_MEMWADDR(10), 
        B_ADDR(10) => fifo_MEMWADDR(9), B_ADDR(9) => 
        fifo_MEMWADDR(8), B_ADDR(8) => fifo_MEMWADDR(7), 
        B_ADDR(7) => fifo_MEMWADDR(6), B_ADDR(6) => 
        fifo_MEMWADDR(5), B_ADDR(5) => fifo_MEMWADDR(4), 
        B_ADDR(4) => fifo_MEMWADDR(3), B_ADDR(3) => 
        fifo_MEMWADDR(2), B_ADDR(2) => fifo_MEMWADDR(1), 
        B_ADDR(1) => fifo_MEMWADDR(0), B_ADDR(0) => GND_net_1, 
        B_WEN(1) => GND_net_1, B_WEN(0) => VCC_net_1, A_EN => 
        VCC_net_1, A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => 
        GND_net_1, A_WIDTH(1) => GND_net_1, A_WIDTH(0) => 
        VCC_net_1, A_WMODE => GND_net_1, B_EN => VCC_net_1, 
        B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => GND_net_1, 
        B_WIDTH(1) => GND_net_1, B_WIDTH(0) => VCC_net_1, B_WMODE
         => GND_net_1, SII_LOCK => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C3 : RAM1K18
      port map(A_DOUT(17) => nc70, A_DOUT(16) => nc62, A_DOUT(15)
         => nc80, A_DOUT(14) => nc130, A_DOUT(13) => nc98, 
        A_DOUT(12) => nc114, A_DOUT(11) => nc56, A_DOUT(10) => 
        nc105, A_DOUT(9) => nc63, A_DOUT(8) => nc97, A_DOUT(7)
         => nc161, A_DOUT(6) => nc31, A_DOUT(5) => nc154, 
        A_DOUT(4) => nc50, A_DOUT(3) => nc142, A_DOUT(2) => nc94, 
        A_DOUT(1) => RDATA_int(7), A_DOUT(0) => RDATA_int(6), 
        B_DOUT(17) => nc122, B_DOUT(16) => nc35, B_DOUT(15) => 
        nc4, B_DOUT(14) => nc92, B_DOUT(13) => nc101, B_DOUT(12)
         => nc166, B_DOUT(11) => nc132, B_DOUT(10) => nc21, 
        B_DOUT(9) => nc93, B_DOUT(8) => nc69, B_DOUT(7) => nc38, 
        B_DOUT(6) => nc113, B_DOUT(5) => nc106, B_DOUT(4) => nc25, 
        B_DOUT(3) => nc1, B_DOUT(2) => nc37, B_DOUT(1) => nc144, 
        B_DOUT(0) => nc153, BUSY => OPEN, A_CLK => 
        m2s010_som_sb_0_CCC_71MHz, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => fifo_MEMRE, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => fifo_MEMRADDR(12), A_ADDR(12) => fifo_MEMRADDR(11), 
        A_ADDR(11) => fifo_MEMRADDR(10), A_ADDR(10) => 
        fifo_MEMRADDR(9), A_ADDR(9) => fifo_MEMRADDR(8), 
        A_ADDR(8) => fifo_MEMRADDR(7), A_ADDR(7) => 
        fifo_MEMRADDR(6), A_ADDR(6) => fifo_MEMRADDR(5), 
        A_ADDR(5) => fifo_MEMRADDR(4), A_ADDR(4) => 
        fifo_MEMRADDR(3), A_ADDR(3) => fifo_MEMRADDR(2), 
        A_ADDR(2) => fifo_MEMRADDR(1), A_ADDR(1) => 
        fifo_MEMRADDR(0), A_ADDR(0) => GND_net_1, A_WEN(1) => 
        GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => GND_net_1, B_DIN(2) => GND_net_1, B_DIN(1)
         => RX_FIFO_DIN_pipe(7), B_DIN(0) => RX_FIFO_DIN_pipe(6), 
        B_ADDR(13) => fifo_MEMWADDR(12), B_ADDR(12) => 
        fifo_MEMWADDR(11), B_ADDR(11) => fifo_MEMWADDR(10), 
        B_ADDR(10) => fifo_MEMWADDR(9), B_ADDR(9) => 
        fifo_MEMWADDR(8), B_ADDR(8) => fifo_MEMWADDR(7), 
        B_ADDR(7) => fifo_MEMWADDR(6), B_ADDR(6) => 
        fifo_MEMWADDR(5), B_ADDR(5) => fifo_MEMWADDR(4), 
        B_ADDR(4) => fifo_MEMWADDR(3), B_ADDR(3) => 
        fifo_MEMWADDR(2), B_ADDR(2) => fifo_MEMWADDR(1), 
        B_ADDR(1) => fifo_MEMWADDR(0), B_ADDR(0) => GND_net_1, 
        B_WEN(1) => GND_net_1, B_WEN(0) => VCC_net_1, A_EN => 
        VCC_net_1, A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => 
        GND_net_1, A_WIDTH(1) => GND_net_1, A_WIDTH(0) => 
        VCC_net_1, A_WMODE => GND_net_1, B_EN => VCC_net_1, 
        B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => GND_net_1, 
        B_WIDTH(1) => GND_net_1, B_WIDTH(0) => VCC_net_1, B_WMODE
         => GND_net_1, SII_LOCK => GND_net_1);
    
    FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top_R0C0 : RAM1K18
      port map(A_DOUT(17) => nc46, A_DOUT(16) => nc71, A_DOUT(15)
         => nc124, A_DOUT(14) => nc81, A_DOUT(13) => nc168, 
        A_DOUT(12) => nc34, A_DOUT(11) => nc28, A_DOUT(10) => 
        nc115, A_DOUT(9) => nc134, A_DOUT(8) => nc32, A_DOUT(7)
         => nc40, A_DOUT(6) => nc99, A_DOUT(5) => nc75, A_DOUT(4)
         => nc85, A_DOUT(3) => nc27, A_DOUT(2) => nc108, 
        A_DOUT(1) => RDATA_int(1), A_DOUT(0) => RDATA_int(0), 
        B_DOUT(17) => nc16, B_DOUT(16) => nc155, B_DOUT(15) => 
        nc51, B_DOUT(14) => nc33, B_DOUT(13) => nc169, B_DOUT(12)
         => nc78, B_DOUT(11) => nc24, B_DOUT(10) => nc88, 
        B_DOUT(9) => nc111, B_DOUT(8) => nc55, B_DOUT(7) => nc10, 
        B_DOUT(6) => nc22, B_DOUT(5) => nc143, B_DOUT(4) => nc77, 
        B_DOUT(3) => nc6, B_DOUT(2) => nc109, B_DOUT(1) => nc87, 
        B_DOUT(0) => nc123, BUSY => OPEN, A_CLK => 
        m2s010_som_sb_0_CCC_71MHz, A_DOUT_CLK => VCC_net_1, 
        A_ARST_N => VCC_net_1, A_DOUT_EN => VCC_net_1, A_BLK(2)
         => fifo_MEMRE, A_BLK(1) => VCC_net_1, A_BLK(0) => 
        VCC_net_1, A_DOUT_ARST_N => VCC_net_1, A_DOUT_SRST_N => 
        VCC_net_1, A_DIN(17) => GND_net_1, A_DIN(16) => GND_net_1, 
        A_DIN(15) => GND_net_1, A_DIN(14) => GND_net_1, A_DIN(13)
         => GND_net_1, A_DIN(12) => GND_net_1, A_DIN(11) => 
        GND_net_1, A_DIN(10) => GND_net_1, A_DIN(9) => GND_net_1, 
        A_DIN(8) => GND_net_1, A_DIN(7) => GND_net_1, A_DIN(6)
         => GND_net_1, A_DIN(5) => GND_net_1, A_DIN(4) => 
        GND_net_1, A_DIN(3) => GND_net_1, A_DIN(2) => GND_net_1, 
        A_DIN(1) => GND_net_1, A_DIN(0) => GND_net_1, A_ADDR(13)
         => fifo_MEMRADDR(12), A_ADDR(12) => fifo_MEMRADDR(11), 
        A_ADDR(11) => fifo_MEMRADDR(10), A_ADDR(10) => 
        fifo_MEMRADDR(9), A_ADDR(9) => fifo_MEMRADDR(8), 
        A_ADDR(8) => fifo_MEMRADDR(7), A_ADDR(7) => 
        fifo_MEMRADDR(6), A_ADDR(6) => fifo_MEMRADDR(5), 
        A_ADDR(5) => fifo_MEMRADDR(4), A_ADDR(4) => 
        fifo_MEMRADDR(3), A_ADDR(3) => fifo_MEMRADDR(2), 
        A_ADDR(2) => fifo_MEMRADDR(1), A_ADDR(1) => 
        fifo_MEMRADDR(0), A_ADDR(0) => GND_net_1, A_WEN(1) => 
        GND_net_1, A_WEN(0) => GND_net_1, B_CLK => 
        CommsFPGA_CCC_0_GL0, B_DOUT_CLK => VCC_net_1, B_ARST_N
         => VCC_net_1, B_DOUT_EN => VCC_net_1, B_BLK(2) => 
        fifo_MEMWE, B_BLK(1) => VCC_net_1, B_BLK(0) => VCC_net_1, 
        B_DOUT_ARST_N => GND_net_1, B_DOUT_SRST_N => VCC_net_1, 
        B_DIN(17) => GND_net_1, B_DIN(16) => GND_net_1, B_DIN(15)
         => GND_net_1, B_DIN(14) => GND_net_1, B_DIN(13) => 
        GND_net_1, B_DIN(12) => GND_net_1, B_DIN(11) => GND_net_1, 
        B_DIN(10) => GND_net_1, B_DIN(9) => GND_net_1, B_DIN(8)
         => GND_net_1, B_DIN(7) => GND_net_1, B_DIN(6) => 
        GND_net_1, B_DIN(5) => GND_net_1, B_DIN(4) => GND_net_1, 
        B_DIN(3) => GND_net_1, B_DIN(2) => GND_net_1, B_DIN(1)
         => RX_FIFO_DIN_pipe(1), B_DIN(0) => RX_FIFO_DIN_pipe(0), 
        B_ADDR(13) => fifo_MEMWADDR(12), B_ADDR(12) => 
        fifo_MEMWADDR(11), B_ADDR(11) => fifo_MEMWADDR(10), 
        B_ADDR(10) => fifo_MEMWADDR(9), B_ADDR(9) => 
        fifo_MEMWADDR(8), B_ADDR(8) => fifo_MEMWADDR(7), 
        B_ADDR(7) => fifo_MEMWADDR(6), B_ADDR(6) => 
        fifo_MEMWADDR(5), B_ADDR(5) => fifo_MEMWADDR(4), 
        B_ADDR(4) => fifo_MEMWADDR(3), B_ADDR(3) => 
        fifo_MEMWADDR(2), B_ADDR(2) => fifo_MEMWADDR(1), 
        B_ADDR(1) => fifo_MEMWADDR(0), B_ADDR(0) => GND_net_1, 
        B_WEN(1) => GND_net_1, B_WEN(0) => VCC_net_1, A_EN => 
        VCC_net_1, A_DOUT_LAT => VCC_net_1, A_WIDTH(2) => 
        GND_net_1, A_WIDTH(1) => GND_net_1, A_WIDTH(0) => 
        VCC_net_1, A_WMODE => GND_net_1, B_EN => VCC_net_1, 
        B_DOUT_LAT => VCC_net_1, B_WIDTH(2) => GND_net_1, 
        B_WIDTH(1) => GND_net_1, B_WIDTH(0) => VCC_net_1, B_WMODE
         => GND_net_1, SII_LOCK => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper is

    port( fifo_MEMRADDR             : in    std_logic_vector(12 downto 0);
          fifo_MEMWADDR             : in    std_logic_vector(12 downto 0);
          RDATA_int                 : out   std_logic_vector(8 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          fifo_MEMRE                : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          fifo_MEMWE                : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top
    port( RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          RDATA_int                 : out   std_logic_vector(8 downto 0);
          fifo_MEMWADDR             : in    std_logic_vector(12 downto 0) := (others => 'U');
          fifo_MEMRADDR             : in    std_logic_vector(12 downto 0) := (others => 'U');
          fifo_MEMWE                : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          fifo_MEMRE                : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    L1_asyncnonpipe : FIFO_8Kx9_FIFO_8Kx9_0_LSRAM_top
      port map(RX_FIFO_DIN_pipe(8) => RX_FIFO_DIN_pipe(8), 
        RX_FIFO_DIN_pipe(7) => RX_FIFO_DIN_pipe(7), 
        RX_FIFO_DIN_pipe(6) => RX_FIFO_DIN_pipe(6), 
        RX_FIFO_DIN_pipe(5) => RX_FIFO_DIN_pipe(5), 
        RX_FIFO_DIN_pipe(4) => RX_FIFO_DIN_pipe(4), 
        RX_FIFO_DIN_pipe(3) => RX_FIFO_DIN_pipe(3), 
        RX_FIFO_DIN_pipe(2) => RX_FIFO_DIN_pipe(2), 
        RX_FIFO_DIN_pipe(1) => RX_FIFO_DIN_pipe(1), 
        RX_FIFO_DIN_pipe(0) => RX_FIFO_DIN_pipe(0), RDATA_int(8)
         => RDATA_int(8), RDATA_int(7) => RDATA_int(7), 
        RDATA_int(6) => RDATA_int(6), RDATA_int(5) => 
        RDATA_int(5), RDATA_int(4) => RDATA_int(4), RDATA_int(3)
         => RDATA_int(3), RDATA_int(2) => RDATA_int(2), 
        RDATA_int(1) => RDATA_int(1), RDATA_int(0) => 
        RDATA_int(0), fifo_MEMWADDR(12) => fifo_MEMWADDR(12), 
        fifo_MEMWADDR(11) => fifo_MEMWADDR(11), fifo_MEMWADDR(10)
         => fifo_MEMWADDR(10), fifo_MEMWADDR(9) => 
        fifo_MEMWADDR(9), fifo_MEMWADDR(8) => fifo_MEMWADDR(8), 
        fifo_MEMWADDR(7) => fifo_MEMWADDR(7), fifo_MEMWADDR(6)
         => fifo_MEMWADDR(6), fifo_MEMWADDR(5) => 
        fifo_MEMWADDR(5), fifo_MEMWADDR(4) => fifo_MEMWADDR(4), 
        fifo_MEMWADDR(3) => fifo_MEMWADDR(3), fifo_MEMWADDR(2)
         => fifo_MEMWADDR(2), fifo_MEMWADDR(1) => 
        fifo_MEMWADDR(1), fifo_MEMWADDR(0) => fifo_MEMWADDR(0), 
        fifo_MEMRADDR(12) => fifo_MEMRADDR(12), fifo_MEMRADDR(11)
         => fifo_MEMRADDR(11), fifo_MEMRADDR(10) => 
        fifo_MEMRADDR(10), fifo_MEMRADDR(9) => fifo_MEMRADDR(9), 
        fifo_MEMRADDR(8) => fifo_MEMRADDR(8), fifo_MEMRADDR(7)
         => fifo_MEMRADDR(7), fifo_MEMRADDR(6) => 
        fifo_MEMRADDR(6), fifo_MEMRADDR(5) => fifo_MEMRADDR(5), 
        fifo_MEMRADDR(4) => fifo_MEMRADDR(4), fifo_MEMRADDR(3)
         => fifo_MEMRADDR(3), fifo_MEMRADDR(2) => 
        fifo_MEMRADDR(2), fifo_MEMRADDR(1) => fifo_MEMRADDR(1), 
        fifo_MEMRADDR(0) => fifo_MEMRADDR(0), fifo_MEMWE => 
        fifo_MEMWE, CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, 
        fifo_MEMRE => fifo_MEMRE, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_0 is

    port( wptr_bin_sync  : inout std_logic_vector(13 downto 0) := (others => 'Z');
          wptr_gray_sync : in    std_logic_vector(12 downto 0)
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_0;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_0 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

begin 


    \bin_out_xhdl1_0_a2[1]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(3), B => wptr_gray_sync(1), C
         => wptr_bin_sync(4), D => wptr_gray_sync(2), Y => 
        wptr_bin_sync(1));
    
    \bin_out_xhdl1_0_a2[10]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(12), B => wptr_gray_sync(11), 
        C => wptr_gray_sync(10), D => wptr_bin_sync(13), Y => 
        wptr_bin_sync(10));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \bin_out_xhdl1_0_a2[5]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(7), B => wptr_gray_sync(6), C
         => wptr_gray_sync(5), D => wptr_bin_sync(8), Y => 
        wptr_bin_sync(5));
    
    \bin_out_xhdl1_0_a2[2]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(4), B => wptr_gray_sync(3), C
         => wptr_gray_sync(2), D => wptr_bin_sync(5), Y => 
        wptr_bin_sync(2));
    
    \bin_out_xhdl1_0_a2[0]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(2), B => wptr_bin_sync(3), C
         => wptr_gray_sync(0), D => wptr_gray_sync(1), Y => 
        wptr_bin_sync(0));
    
    \bin_out_xhdl1_0_a2[9]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(11), B => wptr_gray_sync(10), 
        C => wptr_gray_sync(9), D => wptr_bin_sync(12), Y => 
        wptr_bin_sync(9));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \bin_out_xhdl1_i_o2[12]\ : CFG2
      generic map(INIT => x"6")

      port map(A => wptr_bin_sync(13), B => wptr_gray_sync(12), Y
         => wptr_bin_sync(12));
    
    \bin_out_xhdl1_0_a2[6]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(8), B => wptr_gray_sync(7), C
         => wptr_gray_sync(6), D => wptr_bin_sync(9), Y => 
        wptr_bin_sync(6));
    
    \bin_out_xhdl1_0_a2[4]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(6), B => wptr_gray_sync(5), C
         => wptr_gray_sync(4), D => wptr_bin_sync(7), Y => 
        wptr_bin_sync(4));
    
    \bin_out_xhdl1_i_o2[11]\ : CFG3
      generic map(INIT => x"96")

      port map(A => wptr_gray_sync(12), B => wptr_gray_sync(11), 
        C => wptr_bin_sync(13), Y => wptr_bin_sync(11));
    
    \bin_out_xhdl1_0_a2[8]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(10), B => wptr_gray_sync(9), C
         => wptr_gray_sync(8), D => wptr_bin_sync(11), Y => 
        wptr_bin_sync(8));
    
    \bin_out_xhdl1_0_a2[7]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(9), B => wptr_gray_sync(8), C
         => wptr_gray_sync(7), D => wptr_bin_sync(10), Y => 
        wptr_bin_sync(7));
    
    \bin_out_xhdl1_0_a2[3]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => wptr_gray_sync(5), B => wptr_gray_sync(4), C
         => wptr_gray_sync(3), D => wptr_bin_sync(6), Y => 
        wptr_bin_sync(3));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync is

    port( wptr_gray                 : in    std_logic_vector(13 downto 0);
          wptr_gray_sync            : out   std_logic_vector(12 downto 0);
          wptr_bin_sync_0           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          irx_fifo_rst_i            : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \sync_int[11]_net_1\, GND_net_1, 
        \sync_int[12]_net_1\, \sync_int[13]_net_1\, 
        \sync_int[10]_net_1\, \sync_int[0]_net_1\, 
        \sync_int[1]_net_1\, \sync_int[2]_net_1\, 
        \sync_int[3]_net_1\, \sync_int[4]_net_1\, 
        \sync_int[5]_net_1\, \sync_int[6]_net_1\, 
        \sync_int[7]_net_1\, \sync_int[8]_net_1\, 
        \sync_int[9]_net_1\ : std_logic;

begin 


    \sync_int[9]\ : SLE
      port map(D => wptr_gray(9), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[9]_net_1\);
    
    \sync_int[4]\ : SLE
      port map(D => wptr_gray(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[4]_net_1\);
    
    \sync_out_xhdl1[10]\ : SLE
      port map(D => \sync_int[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(10));
    
    \sync_int[1]\ : SLE
      port map(D => wptr_gray(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[1]_net_1\);
    
    \sync_int[11]\ : SLE
      port map(D => wptr_gray(11), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[11]_net_1\);
    
    \sync_out_xhdl1[6]\ : SLE
      port map(D => \sync_int[6]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(6));
    
    \sync_out_xhdl1[3]\ : SLE
      port map(D => \sync_int[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(3));
    
    \sync_int[6]\ : SLE
      port map(D => wptr_gray(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[6]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \sync_out_xhdl1[11]\ : SLE
      port map(D => \sync_int[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(11));
    
    \sync_int[13]\ : SLE
      port map(D => wptr_gray(13), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[13]_net_1\);
    
    \sync_int[3]\ : SLE
      port map(D => wptr_gray(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[3]_net_1\);
    
    \sync_int[12]\ : SLE
      port map(D => wptr_gray(12), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[12]_net_1\);
    
    \sync_out_xhdl1[4]\ : SLE
      port map(D => \sync_int[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(4));
    
    \sync_int[0]\ : SLE
      port map(D => wptr_gray(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[0]_net_1\);
    
    \sync_out_xhdl1[1]\ : SLE
      port map(D => \sync_int[1]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(1));
    
    \sync_int[5]\ : SLE
      port map(D => wptr_gray(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[5]_net_1\);
    
    \sync_int[2]\ : SLE
      port map(D => wptr_gray(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[2]_net_1\);
    
    \sync_out_xhdl1[12]\ : SLE
      port map(D => \sync_int[12]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(12));
    
    \sync_out_xhdl1[9]\ : SLE
      port map(D => \sync_int[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(9));
    
    \sync_out_xhdl1[2]\ : SLE
      port map(D => \sync_int[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(2));
    
    \sync_int[8]\ : SLE
      port map(D => wptr_gray(8), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[8]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sync_out_xhdl1[7]\ : SLE
      port map(D => \sync_int[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(7));
    
    \sync_out_xhdl1[5]\ : SLE
      port map(D => \sync_int[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(5));
    
    \sync_out_xhdl1[0]\ : SLE
      port map(D => \sync_int[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(0));
    
    \sync_out_xhdl1[8]\ : SLE
      port map(D => \sync_int[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_gray_sync(8));
    
    \sync_int[7]\ : SLE
      port map(D => wptr_gray(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \sync_int[7]_net_1\);
    
    \sync_int[10]\ : SLE
      port map(D => wptr_gray(10), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \sync_int[10]_net_1\);
    
    \sync_out_xhdl1[13]\ : SLE
      port map(D => \sync_int[13]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => wptr_bin_sync_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0 is

    port( rptr_gray           : in    std_logic_vector(13 downto 0);
          rptr_gray_sync      : out   std_logic_vector(12 downto 0);
          rptr_bin_sync_0     : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic;
          irx_fifo_rst_i      : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0 is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal VCC_net_1, \sync_int[13]_net_1\, GND_net_1, 
        \sync_int[12]_net_1\, \sync_int[0]_net_1\, 
        \sync_int[1]_net_1\, \sync_int[2]_net_1\, 
        \sync_int[3]_net_1\, \sync_int[4]_net_1\, 
        \sync_int[5]_net_1\, \sync_int[6]_net_1\, 
        \sync_int[7]_net_1\, \sync_int[8]_net_1\, 
        \sync_int[9]_net_1\, \sync_int[10]_net_1\, 
        \sync_int[11]_net_1\ : std_logic;

begin 


    \sync_int[9]\ : SLE
      port map(D => rptr_gray(9), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[9]_net_1\);
    
    \sync_int[4]\ : SLE
      port map(D => rptr_gray(4), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[4]_net_1\);
    
    \sync_out_xhdl1[10]\ : SLE
      port map(D => \sync_int[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(10));
    
    \sync_int[1]\ : SLE
      port map(D => rptr_gray(1), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[1]_net_1\);
    
    \sync_int[11]\ : SLE
      port map(D => rptr_gray(11), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[11]_net_1\);
    
    \sync_out_xhdl1[6]\ : SLE
      port map(D => \sync_int[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(6));
    
    \sync_out_xhdl1[3]\ : SLE
      port map(D => \sync_int[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(3));
    
    \sync_int[6]\ : SLE
      port map(D => rptr_gray(6), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[6]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \sync_out_xhdl1[11]\ : SLE
      port map(D => \sync_int[11]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(11));
    
    \sync_int[13]\ : SLE
      port map(D => rptr_gray(13), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[13]_net_1\);
    
    \sync_int[3]\ : SLE
      port map(D => rptr_gray(3), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[3]_net_1\);
    
    \sync_int[12]\ : SLE
      port map(D => rptr_gray(12), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[12]_net_1\);
    
    \sync_out_xhdl1[4]\ : SLE
      port map(D => \sync_int[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(4));
    
    \sync_int[0]\ : SLE
      port map(D => rptr_gray(0), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[0]_net_1\);
    
    \sync_out_xhdl1[1]\ : SLE
      port map(D => \sync_int[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(1));
    
    \sync_int[5]\ : SLE
      port map(D => rptr_gray(5), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[5]_net_1\);
    
    \sync_int[2]\ : SLE
      port map(D => rptr_gray(2), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[2]_net_1\);
    
    \sync_out_xhdl1[12]\ : SLE
      port map(D => \sync_int[12]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(12));
    
    \sync_out_xhdl1[9]\ : SLE
      port map(D => \sync_int[9]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(9));
    
    \sync_out_xhdl1[2]\ : SLE
      port map(D => \sync_int[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(2));
    
    \sync_int[8]\ : SLE
      port map(D => rptr_gray(8), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[8]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \sync_out_xhdl1[7]\ : SLE
      port map(D => \sync_int[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(7));
    
    \sync_out_xhdl1[5]\ : SLE
      port map(D => \sync_int[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(5));
    
    \sync_out_xhdl1[0]\ : SLE
      port map(D => \sync_int[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(0));
    
    \sync_out_xhdl1[8]\ : SLE
      port map(D => \sync_int[8]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_gray_sync(8));
    
    \sync_int[7]\ : SLE
      port map(D => rptr_gray(7), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[7]_net_1\);
    
    \sync_int[10]\ : SLE
      port map(D => rptr_gray(10), CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \sync_int[10]_net_1\);
    
    \sync_out_xhdl1[13]\ : SLE
      port map(D => \sync_int[13]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rptr_bin_sync_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3 is

    port( rptr_bin_sync  : inout std_logic_vector(13 downto 0) := (others => 'Z');
          rptr_gray_sync : in    std_logic_vector(12 downto 0);
          bin_N_6_i      : out   std_logic;
          bin_N_4_0_i    : out   std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3;

architecture DEF_ARCH of 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3 is 

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \bin_m5_5\, \bin_m5_4\, \bin_m3_0_3\, \bin_N_4_0_i\, 
        GND_net_1, VCC_net_1 : std_logic;

begin 

    bin_N_4_0_i <= \bin_N_4_0_i\;

    bin_m5_4 : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(4), B => rptr_gray_sync(6), C
         => rptr_gray_sync(5), D => rptr_gray_sync(10), Y => 
        \bin_m5_4\);
    
    \bin_out_xhdl1_0_a2[10]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(12), B => rptr_gray_sync(10), 
        C => rptr_gray_sync(11), D => rptr_bin_sync(13), Y => 
        rptr_bin_sync(10));
    
    \bin_out_xhdl1_0_a2[8]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(8), B => rptr_gray_sync(9), C
         => rptr_bin_sync(10), Y => rptr_bin_sync(8));
    
    bin_m5_5 : CFG4
      generic map(INIT => x"9669")

      port map(A => rptr_gray_sync(8), B => rptr_gray_sync(9), C
         => rptr_gray_sync(7), D => rptr_gray_sync(11), Y => 
        \bin_m5_5\);
    
    bin_m3_0_3 : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(7), B => rptr_gray_sync(9), C
         => rptr_gray_sync(6), D => rptr_gray_sync(10), Y => 
        \bin_m3_0_3\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \bin_out_xhdl1_i_o2_RNIGC583[12]\ : CFG3
      generic map(INIT => x"69")

      port map(A => \bin_m5_5\, B => \bin_m5_4\, C => 
        rptr_bin_sync(12), Y => bin_N_6_i);
    
    \bin_out_xhdl1_0_a2[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(3), B => rptr_gray_sync(2), Y
         => rptr_bin_sync(2));
    
    \bin_out_xhdl1_0_a2[1]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(1), B => rptr_gray_sync(2), C
         => rptr_bin_sync(3), Y => rptr_bin_sync(1));
    
    \bin_out_xhdl1_0_a2[0]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(1), B => rptr_gray_sync(0), C
         => rptr_bin_sync(3), D => rptr_gray_sync(2), Y => 
        rptr_bin_sync(0));
    
    \bin_out_xhdl1_i_o2_RNI3OBE2[12]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(8), B => rptr_gray_sync(11), C
         => rptr_bin_sync(12), D => \bin_m3_0_3\, Y => 
        \bin_N_4_0_i\);
    
    \bin_out_xhdl1_i_o2[11]\ : CFG3
      generic map(INIT => x"96")

      port map(A => rptr_gray_sync(11), B => rptr_bin_sync(13), C
         => rptr_gray_sync(12), Y => rptr_bin_sync(11));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \bin_out_xhdl1_0_a2[7]\ : CFG4
      generic map(INIT => x"6996")

      port map(A => rptr_gray_sync(9), B => rptr_bin_sync(10), C
         => rptr_gray_sync(7), D => rptr_gray_sync(8), Y => 
        rptr_bin_sync(7));
    
    \bin_out_xhdl1_0_a2[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \bin_N_4_0_i\, B => rptr_gray_sync(5), Y => 
        rptr_bin_sync(5));
    
    \bin_out_xhdl1_i_o2[12]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(13), B => rptr_gray_sync(12), Y
         => rptr_bin_sync(12));
    
    \bin_out_xhdl1_0_a2[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rptr_bin_sync(10), B => rptr_gray_sync(9), Y
         => rptr_bin_sync(9));
    
    \bin_out_xhdl1_0_a2[3]\ : CFG4
      generic map(INIT => x"9669")

      port map(A => rptr_bin_sync(12), B => \bin_m5_5\, C => 
        rptr_gray_sync(3), D => \bin_m5_4\, Y => rptr_bin_sync(3));
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3 is

    port( fifo_MEMRADDR             : out   std_logic_vector(12 downto 0);
          fifo_MEMWADDR             : out   std_logic_vector(12 downto 0);
          iRX_FIFO_wr_en_0_0        : in    std_logic;
          iRX_FIFO_rd_en_0          : in    std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          RX_FIFO_TxColDetDis_wr_en : in    std_logic;
          fifo_MEMRE                : out   std_logic;
          fifo_MEMWE                : out   std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          irx_fifo_rst_i            : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3 is 

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_0
    port( wptr_bin_sync  : inout   std_logic_vector(13 downto 0);
          wptr_gray_sync : in    std_logic_vector(12 downto 0) := (others => 'U')
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync
    port( wptr_gray                 : in    std_logic_vector(13 downto 0) := (others => 'U');
          wptr_gray_sync            : out   std_logic_vector(12 downto 0);
          wptr_bin_sync_0           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          irx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0
    port( rptr_gray           : in    std_logic_vector(13 downto 0) := (others => 'U');
          rptr_gray_sync      : out   std_logic_vector(12 downto 0);
          rptr_bin_sync_0     : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          irx_fifo_rst_i      : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3
    port( rptr_bin_sync  : inout   std_logic_vector(13 downto 0);
          rptr_gray_sync : in    std_logic_vector(12 downto 0) := (others => 'U');
          bin_N_6_i      : out   std_logic;
          bin_N_4_0_i    : out   std_logic
        );
  end component;

    signal \rptr[0]_net_1\, \rptr_s[0]\, \wptr[0]_net_1\, 
        \wptr_s[0]\, \fifo_MEMRADDR[0]\, \fifo_MEMRADDR_i[0]\, 
        \fifo_MEMWADDR[0]\, \fifo_MEMWADDR_i[0]\, 
        \rptr_gray[1]_net_1\, VCC_net_1, \rptr_gray_1[1]_net_1\, 
        GND_net_1, \rptr_gray[2]_net_1\, \rptr_gray_1[2]_net_1\, 
        \rptr_gray[3]_net_1\, \rptr_gray_1[3]_net_1\, 
        \rptr_gray[4]_net_1\, \rptr_gray_1[4]_net_1\, 
        \rptr_gray[5]_net_1\, \rptr_gray_1[5]_net_1\, 
        \rptr_gray[6]_net_1\, \rptr_gray_1[6]_net_1\, 
        \rptr_gray[7]_net_1\, \rptr_gray_1[7]_net_1\, 
        \rptr_gray[8]_net_1\, \rptr_gray_1[8]_net_1\, 
        \rptr_gray[9]_net_1\, \rptr_gray_1[9]_net_1\, 
        \rptr_gray[10]_net_1\, \rptr_gray_1[10]_net_1\, 
        \rptr_gray[11]_net_1\, \rptr_gray_1[11]_net_1\, 
        \rptr_gray[12]_net_1\, \rptr_gray_1[12]_net_1\, 
        \rptr_gray[13]_net_1\, \rptr[13]_net_1\, 
        \wptr_gray[0]_net_1\, \wptr_gray_1[0]_net_1\, 
        \wptr_gray[1]_net_1\, \wptr_gray_1[1]_net_1\, 
        \wptr_gray[2]_net_1\, \wptr_gray_1[2]_net_1\, 
        \wptr_gray[3]_net_1\, \wptr_gray_1[3]_net_1\, 
        \wptr_gray[4]_net_1\, \wptr_gray_1[4]_net_1\, 
        \wptr_gray[5]_net_1\, \wptr_gray_1[5]_net_1\, 
        \wptr_gray[6]_net_1\, \wptr_gray_1[6]_net_1\, 
        \wptr_gray[7]_net_1\, \wptr_gray_1[7]_net_1\, 
        \wptr_gray[8]_net_1\, \wptr_gray_1[8]_net_1\, 
        \wptr_gray[9]_net_1\, \wptr_gray_1[9]_net_1\, 
        \wptr_gray[10]_net_1\, \wptr_gray_1[10]_net_1\, 
        \wptr_gray[11]_net_1\, \wptr_gray_1[11]_net_1\, 
        \wptr_gray[12]_net_1\, \wptr_gray_1[12]_net_1\, 
        \wptr_gray[13]_net_1\, \wptr[13]_net_1\, 
        \rptr_gray[0]_net_1\, \rptr_gray_1[0]_net_1\, rdiff_bus, 
        \wptr_bin_sync[0]\, \wptr_bin_sync2[1]_net_1\, 
        \wptr_bin_sync[1]\, \wptr_bin_sync2[2]_net_1\, 
        \wptr_bin_sync[2]\, \wptr_bin_sync2[3]_net_1\, 
        \wptr_bin_sync[3]\, \wptr_bin_sync2[4]_net_1\, 
        \wptr_bin_sync[4]\, \wptr_bin_sync2[5]_net_1\, 
        \wptr_bin_sync[5]\, \wptr_bin_sync2[6]_net_1\, 
        \wptr_bin_sync[6]\, \wptr_bin_sync2[7]_net_1\, 
        \wptr_bin_sync[7]\, \wptr_bin_sync2[8]_net_1\, 
        \wptr_bin_sync[8]\, \wptr_bin_sync2[9]_net_1\, 
        \wptr_bin_sync[9]\, \wptr_bin_sync2[10]_net_1\, 
        \wptr_bin_sync[10]\, \wptr_bin_sync2[11]_net_1\, 
        \wptr_bin_sync[11]\, \wptr_bin_sync2[12]_net_1\, 
        \wptr_bin_sync[12]\, \wptr_bin_sync2[13]_net_1\, 
        \wptr_bin_sync[13]\, \rptr_bin_sync2[9]_net_1\, 
        \rptr_bin_sync[9]\, \rptr_bin_sync2[10]_net_1\, 
        \rptr_bin_sync[10]\, \rptr_bin_sync2[11]_net_1\, 
        \rptr_bin_sync[11]\, \rptr_bin_sync2[12]_net_1\, 
        \rptr_bin_sync[12]\, \rptr_bin_sync2[13]_net_1\, 
        \rptr_bin_sync[13]\, \fifo_MEMWADDR[7]\, 
        \memwaddr_r_2[7]_net_1\, \fifo_MEMWE\, \fifo_MEMWADDR[8]\, 
        \memwaddr_r_2[8]_net_1\, \fifo_MEMWADDR[9]\, 
        \memwaddr_r_2[9]_net_1\, \fifo_MEMWADDR[10]\, 
        \memwaddr_r_2[10]_net_1\, \fifo_MEMWADDR[11]\, 
        \memwaddr_r_2[11]_net_1\, \fifo_MEMWADDR[12]\, 
        \memwaddr_r_2[12]_net_1\, \rptr_bin_sync2[0]_net_1\, 
        \rptr_bin_sync[0]\, \rptr_bin_sync2[1]_net_1\, 
        \rptr_bin_sync[1]\, \rptr_bin_sync2[2]_net_1\, 
        \rptr_bin_sync[2]\, \rptr_bin_sync2[3]_net_1\, 
        \rptr_bin_sync[3]\, \rptr_bin_sync2[4]_net_1\, bin_N_6_i, 
        \rptr_bin_sync2[5]_net_1\, \rptr_bin_sync[5]\, 
        \rptr_bin_sync2[6]_net_1\, bin_N_4_0_i, 
        \rptr_bin_sync2[7]_net_1\, \rptr_bin_sync[7]\, 
        \rptr_bin_sync2[8]_net_1\, \rptr_bin_sync[8]\, 
        \fifo_MEMRADDR[5]\, \memraddr_r_2[5]_net_1\, \fifo_MEMRE\, 
        \fifo_MEMRADDR[6]\, un1_memraddr_r_cry_6_S, 
        \fifo_MEMRADDR[7]\, \memraddr_r_2[7]_net_1\, 
        \fifo_MEMRADDR[8]\, \memraddr_r_2[8]_net_1\, 
        \fifo_MEMRADDR[9]\, \memraddr_r_2[9]_net_1\, 
        \fifo_MEMRADDR[10]\, \memraddr_r_2[10]_net_1\, 
        \fifo_MEMRADDR[11]\, \memraddr_r_2[11]_net_1\, 
        \fifo_MEMRADDR[12]\, \memraddr_r_2[12]_net_1\, 
        \fifo_MEMWADDR[1]\, un1_memwaddr_r_cry_1_S, 
        \fifo_MEMWADDR[2]\, un1_memwaddr_r_cry_2_S, 
        \fifo_MEMWADDR[3]\, un1_memwaddr_r_cry_3_S, 
        \fifo_MEMWADDR[4]\, un1_memwaddr_r_cry_4_S, 
        \fifo_MEMWADDR[5]\, \memwaddr_r_2[5]_net_1\, 
        \fifo_MEMWADDR[6]\, un1_memwaddr_r_cry_6_S, 
        \fifo_MEMRADDR[1]\, un1_memraddr_r_cry_1_S, 
        \fifo_MEMRADDR[2]\, un1_memraddr_r_cry_2_S, 
        \fifo_MEMRADDR[3]\, un1_memraddr_r_cry_3_S, 
        \fifo_MEMRADDR[4]\, un1_memraddr_r_cry_4_S, 
        \iRX_FIFO_Full_0\, fulli, N_6_i, N_5_i, 
        \iRX_FIFO_Empty_0\, empty_r_3, \wptr[1]_net_1\, 
        \wptr_s[1]\, \wptr[2]_net_1\, \wptr_s[2]\, 
        \wptr[3]_net_1\, \wptr_s[3]\, \wptr[4]_net_1\, 
        \wptr_s[4]\, \wptr[5]_net_1\, \wptr_s[5]\, 
        \wptr[6]_net_1\, \wptr_s[6]\, \wptr[7]_net_1\, 
        \wptr_s[7]\, \wptr[8]_net_1\, \wptr_s[8]\, 
        \wptr[9]_net_1\, \wptr_s[9]\, \wptr[10]_net_1\, 
        \wptr_s[10]\, \wptr[11]_net_1\, \wptr_s[11]\, 
        \wptr[12]_net_1\, \wptr_s[12]\, \wptr_s[13]_net_1\, 
        \rptr[1]_net_1\, \rptr_s[1]\, \rptr[2]_net_1\, 
        \rptr_s[2]\, \rptr[3]_net_1\, \rptr_s[3]\, 
        \rptr[4]_net_1\, \rptr_s[4]\, \rptr[5]_net_1\, 
        \rptr_s[5]\, \rptr[6]_net_1\, \rptr_s[6]\, 
        \rptr[7]_net_1\, \rptr_s[7]\, \rptr[8]_net_1\, 
        \rptr_s[8]\, \rptr[9]_net_1\, \rptr_s[9]\, 
        \rptr[10]_net_1\, \rptr_s[10]\, \rptr[11]_net_1\, 
        \rptr_s[11]\, \rptr[12]_net_1\, \rptr_s[12]\, 
        \rptr_s[13]_net_1\, \rdiff_bus_cry_0\, 
        rdiff_bus_cry_0_Y_0, \rdiff_bus_cry_1\, \rdiff_bus[1]\, 
        \rdiff_bus_cry_2\, \rdiff_bus[2]\, \rdiff_bus_cry_3\, 
        \rdiff_bus[3]\, \rdiff_bus_cry_4\, \rdiff_bus[4]\, 
        \rdiff_bus_cry_5\, \rdiff_bus[5]\, \rdiff_bus_cry_6\, 
        \rdiff_bus[6]\, \rdiff_bus_cry_7\, \rdiff_bus[7]\, 
        \rdiff_bus_cry_8\, \rdiff_bus[8]\, \rdiff_bus_cry_9\, 
        \rdiff_bus[9]\, \rdiff_bus_cry_10\, \rdiff_bus[10]\, 
        \rdiff_bus_cry_11\, \rdiff_bus[11]\, \rdiff_bus[13]\, 
        \rdiff_bus_cry_12\, \rdiff_bus[12]\, \wdiff_bus_cry_0\, 
        wdiff_bus_cry_0_Y_0, \wdiff_bus_cry_1\, \wdiff_bus[1]\, 
        \wdiff_bus_cry_2\, \wdiff_bus[2]\, \wdiff_bus_cry_3\, 
        \wdiff_bus[3]\, \wdiff_bus_cry_4\, \wdiff_bus[4]\, 
        \wdiff_bus_cry_5\, \wdiff_bus[5]\, \wdiff_bus_cry_6\, 
        \wdiff_bus[6]\, \wdiff_bus_cry_7\, \wdiff_bus[7]\, 
        \wdiff_bus_cry_8\, \wdiff_bus[8]\, \wdiff_bus_cry_9\, 
        \wdiff_bus[9]\, \wdiff_bus_cry_10\, \wdiff_bus[10]\, 
        \wdiff_bus_cry_11\, \wdiff_bus[11]\, \wdiff_bus[13]\, 
        \wdiff_bus_cry_12\, \wdiff_bus[12]\, rptr_s_908_FCO, 
        \rptr_cry[1]_net_1\, \rptr_cry[2]_net_1\, 
        \rptr_cry[3]_net_1\, \rptr_cry[4]_net_1\, 
        \rptr_cry[5]_net_1\, \rptr_cry[6]_net_1\, 
        \rptr_cry[7]_net_1\, \rptr_cry[8]_net_1\, 
        \rptr_cry[9]_net_1\, \rptr_cry[10]_net_1\, 
        \rptr_cry[11]_net_1\, \rptr_cry[12]_net_1\, 
        wptr_s_909_FCO, \wptr_cry[1]_net_1\, \wptr_cry[2]_net_1\, 
        \wptr_cry[3]_net_1\, \wptr_cry[4]_net_1\, 
        \wptr_cry[5]_net_1\, \wptr_cry[6]_net_1\, 
        \wptr_cry[7]_net_1\, \wptr_cry[8]_net_1\, 
        \wptr_cry[9]_net_1\, \wptr_cry[10]_net_1\, 
        \wptr_cry[11]_net_1\, \wptr_cry[12]_net_1\, 
        un1_memraddr_r_s_1_923_FCO, \un1_memraddr_r_cry_1\, 
        \un1_memraddr_r_cry_2\, \un1_memraddr_r_cry_3\, 
        \un1_memraddr_r_cry_4\, \un1_memraddr_r_cry_5\, 
        un1_memraddr_r_cry_5_S, \un1_memraddr_r_cry_6\, 
        \un1_memraddr_r_cry_7\, un1_memraddr_r_cry_7_S, 
        \un1_memraddr_r_cry_8\, un1_memraddr_r_cry_8_S, 
        \un1_memraddr_r_cry_9\, un1_memraddr_r_cry_9_S, 
        \un1_memraddr_r_cry_10\, un1_memraddr_r_cry_10_S, 
        un1_memraddr_r_s_12_S, \un1_memraddr_r_cry_11\, 
        un1_memraddr_r_cry_11_S, un1_memwaddr_r_s_1_924_FCO, 
        \un1_memwaddr_r_cry_1\, \un1_memwaddr_r_cry_2\, 
        \un1_memwaddr_r_cry_3\, \un1_memwaddr_r_cry_4\, 
        \un1_memwaddr_r_cry_5\, un1_memwaddr_r_cry_5_S, 
        \un1_memwaddr_r_cry_6\, \un1_memwaddr_r_cry_7\, 
        un1_memwaddr_r_cry_7_S, \un1_memwaddr_r_cry_8\, 
        un1_memwaddr_r_cry_8_S, \un1_memwaddr_r_cry_9\, 
        un1_memwaddr_r_cry_9_S, \un1_memwaddr_r_cry_10\, 
        un1_memwaddr_r_cry_10_S, un1_memwaddr_r_s_12_S, 
        \un1_memwaddr_r_cry_11\, un1_memwaddr_r_cry_11_S, 
        \fulli_0_1\, N_12, \fulli_0_a3_3\, empty_r_3_0_a2_3, 
        un4_re_i_0, un4_we_i_0, empty_r_3_0_a2_9, un4_re_i_8, 
        un4_re_i_7, un4_we_i_8, un4_we_i_7, empty_r_3_0_a2_11, 
        un4_re_i_9, un4_we_i_9, N_7, \fulli_0_a3_0_3\, 
        empty_r_3_0_a2_7, \wptr_gray_sync[0]\, 
        \wptr_gray_sync[1]\, \wptr_gray_sync[2]\, 
        \wptr_gray_sync[3]\, \wptr_gray_sync[4]\, 
        \wptr_gray_sync[5]\, \wptr_gray_sync[6]\, 
        \wptr_gray_sync[7]\, \wptr_gray_sync[8]\, 
        \wptr_gray_sync[9]\, \wptr_gray_sync[10]\, 
        \wptr_gray_sync[11]\, \wptr_gray_sync[12]\, 
        \rptr_gray_sync[0]\, \rptr_gray_sync[1]\, 
        \rptr_gray_sync[2]\, \rptr_gray_sync[3]\, 
        \rptr_gray_sync[4]\, \rptr_gray_sync[5]\, 
        \rptr_gray_sync[6]\, \rptr_gray_sync[7]\, 
        \rptr_gray_sync[8]\, \rptr_gray_sync[9]\, 
        \rptr_gray_sync[10]\, \rptr_gray_sync[11]\, 
        \rptr_gray_sync[12]\ : std_logic;
    signal nc2, nc1 : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_0
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_0(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3
	Use entity work.
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3(DEF_ARCH);
begin 

    fifo_MEMRADDR(12) <= \fifo_MEMRADDR[12]\;
    fifo_MEMRADDR(11) <= \fifo_MEMRADDR[11]\;
    fifo_MEMRADDR(10) <= \fifo_MEMRADDR[10]\;
    fifo_MEMRADDR(9) <= \fifo_MEMRADDR[9]\;
    fifo_MEMRADDR(8) <= \fifo_MEMRADDR[8]\;
    fifo_MEMRADDR(7) <= \fifo_MEMRADDR[7]\;
    fifo_MEMRADDR(6) <= \fifo_MEMRADDR[6]\;
    fifo_MEMRADDR(5) <= \fifo_MEMRADDR[5]\;
    fifo_MEMRADDR(4) <= \fifo_MEMRADDR[4]\;
    fifo_MEMRADDR(3) <= \fifo_MEMRADDR[3]\;
    fifo_MEMRADDR(2) <= \fifo_MEMRADDR[2]\;
    fifo_MEMRADDR(1) <= \fifo_MEMRADDR[1]\;
    fifo_MEMRADDR(0) <= \fifo_MEMRADDR[0]\;
    fifo_MEMWADDR(12) <= \fifo_MEMWADDR[12]\;
    fifo_MEMWADDR(11) <= \fifo_MEMWADDR[11]\;
    fifo_MEMWADDR(10) <= \fifo_MEMWADDR[10]\;
    fifo_MEMWADDR(9) <= \fifo_MEMWADDR[9]\;
    fifo_MEMWADDR(8) <= \fifo_MEMWADDR[8]\;
    fifo_MEMWADDR(7) <= \fifo_MEMWADDR[7]\;
    fifo_MEMWADDR(6) <= \fifo_MEMWADDR[6]\;
    fifo_MEMWADDR(5) <= \fifo_MEMWADDR[5]\;
    fifo_MEMWADDR(4) <= \fifo_MEMWADDR[4]\;
    fifo_MEMWADDR(3) <= \fifo_MEMWADDR[3]\;
    fifo_MEMWADDR(2) <= \fifo_MEMWADDR[2]\;
    fifo_MEMWADDR(1) <= \fifo_MEMWADDR[1]\;
    fifo_MEMWADDR(0) <= \fifo_MEMWADDR[0]\;
    iRX_FIFO_Empty_0 <= \iRX_FIFO_Empty_0\;
    iRX_FIFO_Full_0 <= \iRX_FIFO_Full_0\;
    fifo_MEMRE <= \fifo_MEMRE\;
    fifo_MEMWE <= \fifo_MEMWE\;

    \rptr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[4]_net_1\, S
         => \rptr_s[5]\, Y => OPEN, FCO => \rptr_cry[5]_net_1\);
    
    \memwaddr_r_2[9]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_9_S, D => un4_we_i_9, Y => 
        \memwaddr_r_2[9]_net_1\);
    
    wdiff_bus_cry_8 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[8]_net_1\, B => 
        \rptr_bin_sync2[8]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_7\, S => \wdiff_bus[8]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_8\);
    
    \wptr_bin_sync2[12]\ : SLE
      port map(D => \wptr_bin_sync[12]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[12]_net_1\);
    
    \L1.empty_r_3_0_a2_11\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \rdiff_bus[4]\, B => \rdiff_bus[5]\, C => 
        empty_r_3_0_a2_3, D => empty_r_3_0_a2_9, Y => 
        empty_r_3_0_a2_11);
    
    wdiff_bus_cry_11 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[11]_net_1\, B => 
        \rptr_bin_sync2[11]_net_1\, C => GND_net_1, D => 
        GND_net_1, FCI => \wdiff_bus_cry_10\, S => 
        \wdiff_bus[11]\, Y => OPEN, FCO => \wdiff_bus_cry_11\);
    
    \wptr_gray[4]\ : SLE
      port map(D => \wptr_gray_1[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[4]_net_1\);
    
    \rptr_gray_1[3]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[3]_net_1\, B => \rptr[4]_net_1\, Y => 
        \rptr_gray_1[3]_net_1\);
    
    \rptr_bin_sync2[6]\ : SLE
      port map(D => bin_N_4_0_i, CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \rptr_bin_sync2[6]_net_1\);
    
    \rptr[1]\ : SLE
      port map(D => \rptr_s[1]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[1]_net_1\);
    
    fulli_0_a3_0_3 : CFG4
      generic map(INIT => x"8000")

      port map(A => \wdiff_bus[2]\, B => 
        RX_FIFO_TxColDetDis_wr_en, C => iRX_FIFO_wr_en_0_0, D => 
        \wdiff_bus[3]\, Y => \fulli_0_a3_0_3\);
    
    \wptr_gray_1[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[9]_net_1\, B => \wptr[10]_net_1\, Y => 
        \wptr_gray_1[9]_net_1\);
    
    \rptr_gray_1[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[5]_net_1\, B => \rptr[6]_net_1\, Y => 
        \rptr_gray_1[5]_net_1\);
    
    \rptr_gray[9]\ : SLE
      port map(D => \rptr_gray_1[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[9]_net_1\);
    
    un1_memwaddr_r_cry_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_6\, 
        S => un1_memwaddr_r_cry_7_S, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_7\);
    
    un1_memraddr_r_s_1_923 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[0]\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => un1_memraddr_r_s_1_923_FCO);
    
    \rptr_gray[8]\ : SLE
      port map(D => \rptr_gray_1[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[8]_net_1\);
    
    un1_memraddr_r_cry_11 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[11]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_10\, 
        S => un1_memraddr_r_cry_11_S, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_11\);
    
    \rptr_gray_1[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[2]_net_1\, B => \rptr[3]_net_1\, Y => 
        \rptr_gray_1[2]_net_1\);
    
    \rptr_bin_sync2[7]\ : SLE
      port map(D => \rptr_bin_sync[7]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[7]_net_1\);
    
    \memwaddr_r[1]\ : SLE
      port map(D => un1_memwaddr_r_cry_1_S, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[1]\);
    
    \wptr_gray_1[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[7]_net_1\, B => \wptr[8]_net_1\, Y => 
        \wptr_gray_1[7]_net_1\);
    
    \rptr_gray[13]\ : SLE
      port map(D => \rptr[13]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[13]_net_1\);
    
    \memraddr_r[0]\ : SLE
      port map(D => \fifo_MEMRADDR_i[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[0]\);
    
    \memraddr_r_2[9]\ : CFG4
      generic map(INIT => x"7F00")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => un4_re_i_9, 
        D => un1_memraddr_r_cry_9_S, Y => \memraddr_r_2[9]_net_1\);
    
    un1_memwaddr_r_s_1_924 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[0]\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => un1_memwaddr_r_s_1_924_FCO);
    
    \wptr[0]\ : SLE
      port map(D => \wptr_s[0]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[0]_net_1\);
    
    \rptr_bin_sync2[8]\ : SLE
      port map(D => \rptr_bin_sync[8]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[8]_net_1\);
    
    \rptr_gray_1[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[1]_net_1\, B => \rptr[2]_net_1\, Y => 
        \rptr_gray_1[1]_net_1\);
    
    \rptr_gray[10]\ : SLE
      port map(D => \rptr_gray_1[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[10]_net_1\);
    
    \wptr_gray_1[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[0]_net_1\, B => \wptr[1]_net_1\, Y => 
        \wptr_gray_1[0]_net_1\);
    
    wdiff_bus_cry_9 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[9]_net_1\, B => 
        \rptr_bin_sync2[9]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_8\, S => \wdiff_bus[9]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_9\);
    
    \rptr[5]\ : SLE
      port map(D => \rptr_s[5]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[5]_net_1\);
    
    \rptr_gray[3]\ : SLE
      port map(D => \rptr_gray_1[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[3]_net_1\);
    
    \rptr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[5]_net_1\, S
         => \rptr_s[6]\, Y => OPEN, FCO => \rptr_cry[6]_net_1\);
    
    \wptr_gray[3]\ : SLE
      port map(D => \wptr_gray_1[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[3]_net_1\);
    
    \rptr_gray_1[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[10]_net_1\, B => \rptr[11]_net_1\, Y
         => \rptr_gray_1[10]_net_1\);
    
    un1_memraddr_r_cry_10 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_9\, 
        S => un1_memraddr_r_cry_10_S, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_10\);
    
    \rptr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[7]_net_1\, S
         => \rptr_s[8]\, Y => OPEN, FCO => \rptr_cry[8]_net_1\);
    
    \rptr[7]\ : SLE
      port map(D => \rptr_s[7]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[7]_net_1\);
    
    rdiff_bus_cry_4 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[4]_net_1\, B => 
        \rptr[4]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_3\, S => \rdiff_bus[4]\, Y => OPEN, FCO
         => \rdiff_bus_cry_4\);
    
    \rptr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[9]_net_1\, S
         => \rptr_s[10]\, Y => OPEN, FCO => \rptr_cry[10]_net_1\);
    
    \rptr_bin_sync2[12]\ : SLE
      port map(D => \rptr_bin_sync[12]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[12]_net_1\);
    
    memwe_0_a3 : CFG3
      generic map(INIT => x"20")

      port map(A => RX_FIFO_TxColDetDis_wr_en, B => 
        \iRX_FIFO_Full_0\, C => iRX_FIFO_wr_en_0_0, Y => 
        \fifo_MEMWE\);
    
    \rptr_bin_sync2[0]\ : SLE
      port map(D => \rptr_bin_sync[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[0]_net_1\);
    
    \L1.empty_r_3_0_a2_7\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \rdiff_bus[3]\, B => \rdiff_bus[2]\, C => 
        \rdiff_bus[1]\, D => N_7, Y => empty_r_3_0_a2_7);
    
    \wptr[11]\ : SLE
      port map(D => \wptr_s[11]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[11]_net_1\);
    
    rdiff_bus_cry_1 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[1]_net_1\, B => 
        \rptr[1]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_0\, S => \rdiff_bus[1]\, Y => OPEN, FCO
         => \rdiff_bus_cry_1\);
    
    \memraddr_r[1]\ : SLE
      port map(D => un1_memraddr_r_cry_1_S, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[1]\);
    
    \L1.empty_r_3_0_a2_9\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \rdiff_bus[8]\, B => \rdiff_bus[9]\, C => 
        \rdiff_bus[10]\, D => \rdiff_bus[11]\, Y => 
        empty_r_3_0_a2_9);
    
    \rptr_bin_sync2[2]\ : SLE
      port map(D => \rptr_bin_sync[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[2]_net_1\);
    
    \memraddr_r_2[7]\ : CFG4
      generic map(INIT => x"7F00")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => un4_re_i_9, 
        D => un1_memraddr_r_cry_7_S, Y => \memraddr_r_2[7]_net_1\);
    
    un1_memwaddr_r_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_5\, 
        S => un1_memwaddr_r_cry_6_S, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_6\);
    
    rdiff_bus_cry_6 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[6]_net_1\, B => 
        \rptr[6]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_5\, S => \rdiff_bus[6]\, Y => OPEN, FCO
         => \rdiff_bus_cry_6\);
    
    \memwaddr_r_2[10]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_10_S, D => un4_we_i_9, Y => 
        \memwaddr_r_2[10]_net_1\);
    
    \memraddr_r_2[5]\ : CFG4
      generic map(INIT => x"7F00")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => un4_re_i_9, 
        D => un1_memraddr_r_cry_5_S, Y => \memraddr_r_2[5]_net_1\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    un1_memwaddr_r_cry_9 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[9]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_8\, 
        S => un1_memwaddr_r_cry_9_S, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_9\);
    
    \rptr_gray[1]\ : SLE
      port map(D => \rptr_gray_1[1]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[1]_net_1\);
    
    \memwaddr_r[7]\ : SLE
      port map(D => \memwaddr_r_2[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[7]\);
    
    \wptr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[3]_net_1\, S
         => \wptr_s[4]\, Y => OPEN, FCO => \wptr_cry[4]_net_1\);
    
    \wptr_gray_1[12]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[13]_net_1\, B => \wptr[12]_net_1\, Y
         => \wptr_gray_1[12]_net_1\);
    
    \wptr[12]\ : SLE
      port map(D => \wptr_s[12]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[12]_net_1\);
    
    \L1.empty_r_3_0_o2\ : CFG2
      generic map(INIT => x"E")

      port map(A => rdiff_bus_cry_0_Y_0, B => iRX_FIFO_rd_en_0, Y
         => N_7);
    
    \wptr_cry[10]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[10]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[9]_net_1\, S
         => \wptr_s[10]\, Y => OPEN, FCO => \wptr_cry[10]_net_1\);
    
    wdiff_bus_cry_5 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[5]_net_1\, B => 
        \rptr_bin_sync2[5]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_4\, S => \wdiff_bus[5]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_5\);
    
    \rptr_gray[12]\ : SLE
      port map(D => \rptr_gray_1[12]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[12]_net_1\);
    
    \memwaddr_r[4]\ : SLE
      port map(D => un1_memwaddr_r_cry_4_S, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[4]\);
    
    \wptr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[1]_net_1\, S
         => \wptr_s[2]\, Y => OPEN, FCO => \wptr_cry[2]_net_1\);
    
    \memraddr_r_2[10]\ : CFG4
      generic map(INIT => x"7F00")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => un4_re_i_9, 
        D => un1_memraddr_r_cry_10_S, Y => 
        \memraddr_r_2[10]_net_1\);
    
    rdiff_bus_cry_11 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[11]_net_1\, B => 
        \rptr[11]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_10\, S => \rdiff_bus[11]\, Y => OPEN, FCO
         => \rdiff_bus_cry_11\);
    
    wdiff_bus_cry_0 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[0]_net_1\, B => 
        \rptr_bin_sync2[0]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => VCC_net_1, S => OPEN, Y => wdiff_bus_cry_0_Y_0, 
        FCO => \wdiff_bus_cry_0\);
    
    \wptr[1]\ : SLE
      port map(D => \wptr_s[1]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[1]_net_1\);
    
    \rptr_bin_sync2[4]\ : SLE
      port map(D => bin_N_6_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[4]_net_1\);
    
    \wptr_bin_sync2[6]\ : SLE
      port map(D => \wptr_bin_sync[6]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[6]_net_1\);
    
    \rptr[3]\ : SLE
      port map(D => \rptr_s[3]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[3]_net_1\);
    
    \wptr_gray[13]\ : SLE
      port map(D => \wptr[13]_net_1\, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr_gray[13]_net_1\);
    
    \wptr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[2]_net_1\, S
         => \wptr_s[3]\, Y => OPEN, FCO => \wptr_cry[3]_net_1\);
    
    \rptr[6]\ : SLE
      port map(D => \rptr_s[6]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[6]_net_1\);
    
    rdiff_bus_cry_8 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[8]_net_1\, B => 
        \rptr[8]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_7\, S => \rdiff_bus[8]\, Y => OPEN, FCO
         => \rdiff_bus_cry_8\);
    
    \wptr_gray[10]\ : SLE
      port map(D => \wptr_gray_1[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[10]_net_1\);
    
    rdiff_bus_cry_7 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[7]_net_1\, B => 
        \rptr[7]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_6\, S => \rdiff_bus[7]\, Y => OPEN, FCO
         => \rdiff_bus_cry_7\);
    
    \wptr_bin_sync2[7]\ : SLE
      port map(D => \wptr_bin_sync[7]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[7]_net_1\);
    
    \rptr_gray_1[11]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[11]_net_1\, B => \rptr[12]_net_1\, Y
         => \rptr_gray_1[11]_net_1\);
    
    \rptr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[8]_net_1\, S
         => \rptr_s[9]\, Y => OPEN, FCO => \rptr_cry[9]_net_1\);
    
    un1_memwaddr_r_cry_1 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[1]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        un1_memwaddr_r_s_1_924_FCO, S => un1_memwaddr_r_cry_1_S, 
        Y => OPEN, FCO => \un1_memwaddr_r_cry_1\);
    
    \rptr_gray[5]\ : SLE
      port map(D => \rptr_gray_1[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[5]_net_1\);
    
    un1_memwaddr_r_s_12 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[12]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_11\, 
        S => un1_memwaddr_r_s_12_S, Y => OPEN, FCO => OPEN);
    
    \wptr_gray_1[2]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[2]_net_1\, B => \wptr[3]_net_1\, Y => 
        \wptr_gray_1[2]_net_1\);
    
    rptr_s_908 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => rptr_s_908_FCO);
    
    \wptr[5]\ : SLE
      port map(D => \wptr_s[5]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[5]_net_1\);
    
    rdiff_bus_cry_5 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[5]_net_1\, B => 
        \rptr[5]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_4\, S => \rdiff_bus[5]\, Y => OPEN, FCO
         => \rdiff_bus_cry_5\);
    
    \wptr_bin_sync2[8]\ : SLE
      port map(D => \wptr_bin_sync[8]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[8]_net_1\);
    
    fulli_0_a3_3 : CFG4
      generic map(INIT => x"8000")

      port map(A => \wdiff_bus[7]\, B => \wdiff_bus[8]\, C => 
        \wdiff_bus[9]\, D => \wdiff_bus[10]\, Y => \fulli_0_a3_3\);
    
    \wptr[7]\ : SLE
      port map(D => \wptr_s[7]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[7]_net_1\);
    
    un1_memwaddr_r_cry_2 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[2]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_1\, 
        S => un1_memwaddr_r_cry_2_S, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_2\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \wptr_gray[1]\ : SLE
      port map(D => \wptr_gray_1[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[1]_net_1\);
    
    \rptr_gray_1[9]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[9]_net_1\, B => \rptr[10]_net_1\, Y => 
        \rptr_gray_1[9]_net_1\);
    
    \rptr_bin_sync2[5]\ : SLE
      port map(D => \rptr_bin_sync[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[5]_net_1\);
    
    \rptr_bin_sync2[1]\ : SLE
      port map(D => \rptr_bin_sync[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[1]_net_1\);
    
    \memwaddr_r[10]\ : SLE
      port map(D => \memwaddr_r_2[10]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[10]\);
    
    wdiff_bus_cry_7 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[7]_net_1\, B => 
        \rptr_bin_sync2[7]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_6\, S => \wdiff_bus[7]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_7\);
    
    \wptr_bin_sync2[0]\ : SLE
      port map(D => \wptr_bin_sync[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => rdiff_bus);
    
    un1_memwaddr_r_cry_8 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[8]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_7\, 
        S => un1_memwaddr_r_cry_8_S, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_8\);
    
    \wptr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => wptr_s_909_FCO, S => 
        \wptr_s[1]\, Y => OPEN, FCO => \wptr_cry[1]_net_1\);
    
    un1_memwaddr_r_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_3\, 
        S => un1_memwaddr_r_cry_4_S, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_4\);
    
    un1_memwaddr_r_cry_3 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[3]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_2\, 
        S => un1_memwaddr_r_cry_3_S, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_3\);
    
    \memraddr_r[8]\ : SLE
      port map(D => \memraddr_r_2[8]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[8]\);
    
    \rptr[9]\ : SLE
      port map(D => \rptr_s[9]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[9]_net_1\);
    
    \wptr_gray_1[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[6]_net_1\, B => \wptr[7]_net_1\, Y => 
        \wptr_gray_1[6]_net_1\);
    
    \wptr_gray[12]\ : SLE
      port map(D => \wptr_gray_1[12]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[12]_net_1\);
    
    \wptr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[6]_net_1\, S
         => \wptr_s[7]\, Y => OPEN, FCO => \wptr_cry[7]_net_1\);
    
    \wptr_bin_sync2[2]\ : SLE
      port map(D => \wptr_bin_sync[2]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[2]_net_1\);
    
    fulli_0_1 : CFG4
      generic map(INIT => x"01FF")

      port map(A => \wdiff_bus[6]\, B => \wdiff_bus[5]\, C => 
        N_12, D => \fulli_0_a3_3\, Y => \fulli_0_1\);
    
    \L1.un4_re_i_9\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \fifo_MEMRADDR[11]\, B => \fifo_MEMRADDR[10]\, 
        C => \fifo_MEMRADDR[0]\, D => un4_re_i_0, Y => un4_re_i_9);
    
    un1_memraddr_r_cry_3 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[3]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_2\, 
        S => un1_memraddr_r_cry_3_S, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_3\);
    
    \rptr_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \rptr[0]_net_1\, Y => \rptr_s[0]\);
    
    un1_memraddr_r_cry_1 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[1]\, C => 
        GND_net_1, D => GND_net_1, FCI => 
        un1_memraddr_r_s_1_923_FCO, S => un1_memraddr_r_cry_1_S, 
        Y => OPEN, FCO => \un1_memraddr_r_cry_1\);
    
    \rptr[4]\ : SLE
      port map(D => \rptr_s[4]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[4]_net_1\);
    
    \memwaddr_r_2[5]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_5_S, D => un4_we_i_9, Y => 
        \memwaddr_r_2[5]_net_1\);
    
    \wptr_gray[6]\ : SLE
      port map(D => \wptr_gray_1[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[6]_net_1\);
    
    \wptr_gray_1[3]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[3]_net_1\, B => \wptr[4]_net_1\, Y => 
        \wptr_gray_1[3]_net_1\);
    
    \wptr_cry[5]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[5]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[4]_net_1\, S
         => \wptr_s[5]\, Y => OPEN, FCO => \wptr_cry[5]_net_1\);
    
    un1_memraddr_r_cry_9 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[9]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_8\, 
        S => un1_memraddr_r_cry_9_S, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_9\);
    
    fulli_0_a3_0 : CFG4
      generic map(INIT => x"4000")

      port map(A => wdiff_bus_cry_0_Y_0, B => \wdiff_bus[1]\, C
         => \wdiff_bus[4]\, D => \fulli_0_a3_0_3\, Y => N_12);
    
    \rptr_gray[4]\ : SLE
      port map(D => \rptr_gray_1[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[4]_net_1\);
    
    un1_memraddr_r_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_4\, 
        S => un1_memraddr_r_cry_5_S, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_5\);
    
    \wptr_bin_sync2[4]\ : SLE
      port map(D => \wptr_bin_sync[4]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[4]_net_1\);
    
    \wptr[3]\ : SLE
      port map(D => \wptr_s[3]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[3]_net_1\);
    
    \L1.un4_we_i_9\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \fifo_MEMWADDR[4]\, B => \fifo_MEMWADDR[3]\, 
        C => \fifo_MEMWADDR[0]\, D => un4_we_i_0, Y => un4_we_i_9);
    
    \memwaddr_r[6]\ : SLE
      port map(D => un1_memwaddr_r_cry_6_S, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[6]\);
    
    \wptr[6]\ : SLE
      port map(D => \wptr_s[6]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[6]_net_1\);
    
    \memwaddr_r[9]\ : SLE
      port map(D => \memwaddr_r_2[9]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[9]\);
    
    \memraddr_r[10]\ : SLE
      port map(D => \memraddr_r_2[10]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[10]\);
    
    \L1.un4_re_i_8\ : CFG4
      generic map(INIT => x"0080")

      port map(A => \fifo_MEMRADDR[9]\, B => \fifo_MEMRADDR[8]\, 
        C => \fifo_MEMRADDR[7]\, D => \fifo_MEMRADDR[6]\, Y => 
        un4_re_i_8);
    
    \memwaddr_r[3]\ : SLE
      port map(D => un1_memwaddr_r_cry_3_S, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[3]\);
    
    \rptr_gray_1[12]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[13]_net_1\, B => \rptr[12]_net_1\, Y
         => \rptr_gray_1[12]_net_1\);
    
    full_r : SLE
      port map(D => fulli, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \iRX_FIFO_Full_0\);
    
    \rptr_bin_sync2[3]\ : SLE
      port map(D => \rptr_bin_sync[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[3]_net_1\);
    
    \wptr_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \wptr[0]_net_1\, Y => \wptr_s[0]\);
    
    \rptr[2]\ : SLE
      port map(D => \rptr_s[2]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[2]_net_1\);
    
    \memraddr_r[3]\ : SLE
      port map(D => un1_memraddr_r_cry_3_S, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[3]\);
    
    \wptr[13]\ : SLE
      port map(D => \wptr_s[13]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \wptr[13]_net_1\);
    
    \rptr_bin_sync2[9]\ : SLE
      port map(D => \rptr_bin_sync[9]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[9]_net_1\);
    
    \wptr_bin_sync2[13]\ : SLE
      port map(D => \wptr_bin_sync[13]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[13]_net_1\);
    
    \rptr[11]\ : SLE
      port map(D => \rptr_s[11]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rptr[11]_net_1\);
    
    \wptr_cry[6]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[6]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[5]_net_1\, S
         => \wptr_s[6]\, Y => OPEN, FCO => \wptr_cry[6]_net_1\);
    
    \rptr_bin_sync2[11]\ : SLE
      port map(D => \rptr_bin_sync[11]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[11]_net_1\);
    
    \wptr_bin_sync2[5]\ : SLE
      port map(D => \wptr_bin_sync[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[5]_net_1\);
    
    \L1.un4_we_i_8\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \fifo_MEMWADDR[10]\, B => \fifo_MEMWADDR[9]\, 
        C => \fifo_MEMWADDR[8]\, D => \fifo_MEMWADDR[7]\, Y => 
        un4_we_i_8);
    
    \wptr_cry[8]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[8]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[7]_net_1\, S
         => \wptr_s[8]\, Y => OPEN, FCO => \wptr_cry[8]_net_1\);
    
    \wptr_bin_sync2[1]\ : SLE
      port map(D => \wptr_bin_sync[1]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[1]_net_1\);
    
    Wr_corefifo_grayToBinConv : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3_0
      port map(wptr_bin_sync(13) => \wptr_bin_sync[13]\, 
        wptr_bin_sync(12) => \wptr_bin_sync[12]\, 
        wptr_bin_sync(11) => \wptr_bin_sync[11]\, 
        wptr_bin_sync(10) => \wptr_bin_sync[10]\, 
        wptr_bin_sync(9) => \wptr_bin_sync[9]\, wptr_bin_sync(8)
         => \wptr_bin_sync[8]\, wptr_bin_sync(7) => 
        \wptr_bin_sync[7]\, wptr_bin_sync(6) => 
        \wptr_bin_sync[6]\, wptr_bin_sync(5) => 
        \wptr_bin_sync[5]\, wptr_bin_sync(4) => 
        \wptr_bin_sync[4]\, wptr_bin_sync(3) => 
        \wptr_bin_sync[3]\, wptr_bin_sync(2) => 
        \wptr_bin_sync[2]\, wptr_bin_sync(1) => 
        \wptr_bin_sync[1]\, wptr_bin_sync(0) => 
        \wptr_bin_sync[0]\, wptr_gray_sync(12) => 
        \wptr_gray_sync[12]\, wptr_gray_sync(11) => 
        \wptr_gray_sync[11]\, wptr_gray_sync(10) => 
        \wptr_gray_sync[10]\, wptr_gray_sync(9) => 
        \wptr_gray_sync[9]\, wptr_gray_sync(8) => 
        \wptr_gray_sync[8]\, wptr_gray_sync(7) => 
        \wptr_gray_sync[7]\, wptr_gray_sync(6) => 
        \wptr_gray_sync[6]\, wptr_gray_sync(5) => 
        \wptr_gray_sync[5]\, wptr_gray_sync(4) => 
        \wptr_gray_sync[4]\, wptr_gray_sync(3) => 
        \wptr_gray_sync[3]\, wptr_gray_sync(2) => 
        \wptr_gray_sync[2]\, wptr_gray_sync(1) => 
        \wptr_gray_sync[1]\, wptr_gray_sync(0) => 
        \wptr_gray_sync[0]\);
    
    \wptr_gray_1[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[4]_net_1\, B => \wptr[5]_net_1\, Y => 
        \wptr_gray_1[4]_net_1\);
    
    \rptr_bin_sync2[13]\ : SLE
      port map(D => \rptr_bin_sync[13]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[13]_net_1\);
    
    \L1.un4_re_i_7\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \fifo_MEMRADDR[4]\, B => \fifo_MEMRADDR[3]\, 
        C => \fifo_MEMRADDR[2]\, D => \fifo_MEMRADDR[1]\, Y => 
        un4_re_i_7);
    
    overflow_r : SLE
      port map(D => N_6_i, CLK => CommsFPGA_CCC_0_GL0, EN => 
        VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        iRX_FIFO_OVERFLOW_0);
    
    fulli_0 : CFG4
      generic map(INIT => x"BAAA")

      port map(A => \wdiff_bus[13]\, B => \fulli_0_1\, C => 
        \wdiff_bus[11]\, D => \wdiff_bus[12]\, Y => fulli);
    
    \memraddr_r_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \fifo_MEMRADDR[0]\, Y => \fifo_MEMRADDR_i[0]\);
    
    \memraddr_r_2[8]\ : CFG4
      generic map(INIT => x"7F00")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => un4_re_i_9, 
        D => un1_memraddr_r_cry_8_S, Y => \memraddr_r_2[8]_net_1\);
    
    \rptr_gray[11]\ : SLE
      port map(D => \rptr_gray_1[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[11]_net_1\);
    
    \wptr_bin_sync2[10]\ : SLE
      port map(D => \wptr_bin_sync[10]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[10]_net_1\);
    
    \rptr[10]\ : SLE
      port map(D => \rptr_s[10]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rptr[10]_net_1\);
    
    \wptr[9]\ : SLE
      port map(D => \wptr_s[9]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[9]_net_1\);
    
    Wr_corefifo_doubleSync : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync
      port map(wptr_gray(13) => \wptr_gray[13]_net_1\, 
        wptr_gray(12) => \wptr_gray[12]_net_1\, wptr_gray(11) => 
        \wptr_gray[11]_net_1\, wptr_gray(10) => 
        \wptr_gray[10]_net_1\, wptr_gray(9) => 
        \wptr_gray[9]_net_1\, wptr_gray(8) => 
        \wptr_gray[8]_net_1\, wptr_gray(7) => 
        \wptr_gray[7]_net_1\, wptr_gray(6) => 
        \wptr_gray[6]_net_1\, wptr_gray(5) => 
        \wptr_gray[5]_net_1\, wptr_gray(4) => 
        \wptr_gray[4]_net_1\, wptr_gray(3) => 
        \wptr_gray[3]_net_1\, wptr_gray(2) => 
        \wptr_gray[2]_net_1\, wptr_gray(1) => 
        \wptr_gray[1]_net_1\, wptr_gray(0) => 
        \wptr_gray[0]_net_1\, wptr_gray_sync(12) => 
        \wptr_gray_sync[12]\, wptr_gray_sync(11) => 
        \wptr_gray_sync[11]\, wptr_gray_sync(10) => 
        \wptr_gray_sync[10]\, wptr_gray_sync(9) => 
        \wptr_gray_sync[9]\, wptr_gray_sync(8) => 
        \wptr_gray_sync[8]\, wptr_gray_sync(7) => 
        \wptr_gray_sync[7]\, wptr_gray_sync(6) => 
        \wptr_gray_sync[6]\, wptr_gray_sync(5) => 
        \wptr_gray_sync[5]\, wptr_gray_sync(4) => 
        \wptr_gray_sync[4]\, wptr_gray_sync(3) => 
        \wptr_gray_sync[3]\, wptr_gray_sync(2) => 
        \wptr_gray_sync[2]\, wptr_gray_sync(1) => 
        \wptr_gray_sync[1]\, wptr_gray_sync(0) => 
        \wptr_gray_sync[0]\, wptr_bin_sync_0 => 
        \wptr_bin_sync[13]\, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, irx_fifo_rst_i => 
        irx_fifo_rst_i);
    
    un1_memwaddr_r_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[5]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_4\, 
        S => un1_memwaddr_r_cry_5_S, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_5\);
    
    \rptr_gray[0]\ : SLE
      port map(D => \rptr_gray_1[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[0]_net_1\);
    
    empty_r : SLE
      port map(D => empty_r_3, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \iRX_FIFO_Empty_0\);
    
    \memwaddr_r_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \fifo_MEMWADDR[0]\, Y => \fifo_MEMWADDR_i[0]\);
    
    \L1.empty_r_3_0_a2_3\ : CFG2
      generic map(INIT => x"1")

      port map(A => \rdiff_bus[7]\, B => \rdiff_bus[6]\, Y => 
        empty_r_3_0_a2_3);
    
    \memwaddr_r_2[12]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_s_12_S, D => un4_we_i_9, Y => 
        \memwaddr_r_2[12]_net_1\);
    
    \rptr_gray_1[7]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[7]_net_1\, B => \rptr[8]_net_1\, Y => 
        \rptr_gray_1[7]_net_1\);
    
    un1_memraddr_r_cry_2 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[2]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_1\, 
        S => un1_memraddr_r_cry_2_S, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_2\);
    
    wdiff_bus_cry_12 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[12]_net_1\, B => 
        \rptr_bin_sync2[12]_net_1\, C => GND_net_1, D => 
        GND_net_1, FCI => \wdiff_bus_cry_11\, S => 
        \wdiff_bus[12]\, Y => OPEN, FCO => \wdiff_bus_cry_12\);
    
    \wptr[4]\ : SLE
      port map(D => \wptr_s[4]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[4]_net_1\);
    
    un1_memraddr_r_cry_8 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[8]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_7\, 
        S => un1_memraddr_r_cry_8_S, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_8\);
    
    \rptr_s[13]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[13]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[12]_net_1\, S
         => \rptr_s[13]_net_1\, Y => OPEN, FCO => OPEN);
    
    \memwaddr_r[8]\ : SLE
      port map(D => \memwaddr_r_2[8]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[8]\);
    
    \memwaddr_r[2]\ : SLE
      port map(D => un1_memwaddr_r_cry_2_S, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[2]\);
    
    \wptr_bin_sync2[11]\ : SLE
      port map(D => \wptr_bin_sync[11]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[11]_net_1\);
    
    \L1.un4_we_i_7\ : CFG4
      generic map(INIT => x"0008")

      port map(A => \fifo_MEMWADDR[12]\, B => \fifo_MEMWADDR[11]\, 
        C => \fifo_MEMWADDR[6]\, D => \fifo_MEMWADDR[5]\, Y => 
        un4_we_i_7);
    
    \wptr_gray_1[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[1]_net_1\, B => \wptr[2]_net_1\, Y => 
        \wptr_gray_1[1]_net_1\);
    
    underflow_r : SLE
      port map(D => N_5_i, CLK => m2s010_som_sb_0_CCC_71MHz, EN
         => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => iRX_FIFO_UNDERRUN_0);
    
    \memwaddr_r_2[11]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_11_S, D => un4_we_i_9, Y => 
        \memwaddr_r_2[11]_net_1\);
    
    \memraddr_r_2[12]\ : CFG4
      generic map(INIT => x"7F00")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => un4_re_i_9, 
        D => un1_memraddr_r_s_12_S, Y => \memraddr_r_2[12]_net_1\);
    
    \wptr_gray[5]\ : SLE
      port map(D => \wptr_gray_1[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[5]_net_1\);
    
    overflow_r_RNO : CFG3
      generic map(INIT => x"80")

      port map(A => RX_FIFO_TxColDetDis_wr_en, B => 
        \iRX_FIFO_Full_0\, C => iRX_FIFO_wr_en_0_0, Y => N_6_i);
    
    \memraddr_r[7]\ : SLE
      port map(D => \memraddr_r_2[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[7]\);
    
    un1_memraddr_r_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[6]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_5\, 
        S => un1_memraddr_r_cry_6_S, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_6\);
    
    \rptr_bin_sync2[10]\ : SLE
      port map(D => \rptr_bin_sync[10]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_bin_sync2[10]_net_1\);
    
    wdiff_bus_s_13 : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \rptr_bin_sync2[13]_net_1\, C
         => \wptr[13]_net_1\, D => GND_net_1, FCI => 
        \wdiff_bus_cry_12\, S => \wdiff_bus[13]\, Y => OPEN, FCO
         => OPEN);
    
    wdiff_bus_cry_10 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[10]_net_1\, B => 
        \rptr_bin_sync2[10]_net_1\, C => GND_net_1, D => 
        GND_net_1, FCI => \wdiff_bus_cry_9\, S => \wdiff_bus[10]\, 
        Y => OPEN, FCO => \wdiff_bus_cry_10\);
    
    \memwaddr_r[11]\ : SLE
      port map(D => \memwaddr_r_2[11]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[11]\);
    
    \wptr_gray[8]\ : SLE
      port map(D => \wptr_gray_1[8]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[8]_net_1\);
    
    \memraddr_r_2[11]\ : CFG4
      generic map(INIT => x"7F00")

      port map(A => un4_re_i_8, B => un4_re_i_7, C => un4_re_i_9, 
        D => un1_memraddr_r_cry_11_S, Y => 
        \memraddr_r_2[11]_net_1\);
    
    un1_memraddr_r_s_12 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[12]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_11\, 
        S => un1_memraddr_r_s_12_S, Y => OPEN, FCO => OPEN);
    
    \wptr_gray[7]\ : SLE
      port map(D => \wptr_gray_1[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[7]_net_1\);
    
    \wptr_gray_1[5]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[5]_net_1\, B => \wptr[6]_net_1\, Y => 
        \wptr_gray_1[5]_net_1\);
    
    \memwaddr_r[5]\ : SLE
      port map(D => \memwaddr_r_2[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[5]\);
    
    \L1.empty_r_3_0_a2\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \rdiff_bus[12]\, B => \rdiff_bus[13]\, C => 
        empty_r_3_0_a2_7, D => empty_r_3_0_a2_11, Y => empty_r_3);
    
    un1_memraddr_r_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[4]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_3\, 
        S => un1_memraddr_r_cry_4_S, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_4\);
    
    \rptr[8]\ : SLE
      port map(D => \rptr_s[8]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[8]_net_1\);
    
    Rd_corefifo_doubleSync : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_doubleSync_0
      port map(rptr_gray(13) => \rptr_gray[13]_net_1\, 
        rptr_gray(12) => \rptr_gray[12]_net_1\, rptr_gray(11) => 
        \rptr_gray[11]_net_1\, rptr_gray(10) => 
        \rptr_gray[10]_net_1\, rptr_gray(9) => 
        \rptr_gray[9]_net_1\, rptr_gray(8) => 
        \rptr_gray[8]_net_1\, rptr_gray(7) => 
        \rptr_gray[7]_net_1\, rptr_gray(6) => 
        \rptr_gray[6]_net_1\, rptr_gray(5) => 
        \rptr_gray[5]_net_1\, rptr_gray(4) => 
        \rptr_gray[4]_net_1\, rptr_gray(3) => 
        \rptr_gray[3]_net_1\, rptr_gray(2) => 
        \rptr_gray[2]_net_1\, rptr_gray(1) => 
        \rptr_gray[1]_net_1\, rptr_gray(0) => 
        \rptr_gray[0]_net_1\, rptr_gray_sync(12) => 
        \rptr_gray_sync[12]\, rptr_gray_sync(11) => 
        \rptr_gray_sync[11]\, rptr_gray_sync(10) => 
        \rptr_gray_sync[10]\, rptr_gray_sync(9) => 
        \rptr_gray_sync[9]\, rptr_gray_sync(8) => 
        \rptr_gray_sync[8]\, rptr_gray_sync(7) => 
        \rptr_gray_sync[7]\, rptr_gray_sync(6) => 
        \rptr_gray_sync[6]\, rptr_gray_sync(5) => 
        \rptr_gray_sync[5]\, rptr_gray_sync(4) => 
        \rptr_gray_sync[4]\, rptr_gray_sync(3) => 
        \rptr_gray_sync[3]\, rptr_gray_sync(2) => 
        \rptr_gray_sync[2]\, rptr_gray_sync(1) => 
        \rptr_gray_sync[1]\, rptr_gray_sync(0) => 
        \rptr_gray_sync[0]\, rptr_bin_sync_0 => 
        \rptr_bin_sync[13]\, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, irx_fifo_rst_i => irx_fifo_rst_i);
    
    underflow_r_RNO : CFG2
      generic map(INIT => x"8")

      port map(A => iRX_FIFO_rd_en_0, B => \iRX_FIFO_Empty_0\, Y
         => N_5_i);
    
    \rptr_cry[4]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[4]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[3]_net_1\, S
         => \rptr_s[4]\, Y => OPEN, FCO => \rptr_cry[4]_net_1\);
    
    wptr_s_909 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => wptr_s_909_FCO);
    
    wdiff_bus_cry_2 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[2]_net_1\, B => 
        \rptr_bin_sync2[2]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_1\, S => \wdiff_bus[2]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_2\);
    
    \rptr_gray[2]\ : SLE
      port map(D => \rptr_gray_1[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[2]_net_1\);
    
    \wptr_cry[9]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[9]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[8]_net_1\, S
         => \wptr_s[9]\, Y => OPEN, FCO => \wptr_cry[9]_net_1\);
    
    \wptr_bin_sync2[3]\ : SLE
      port map(D => \wptr_bin_sync[3]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[3]_net_1\);
    
    \rptr[12]\ : SLE
      port map(D => \rptr_s[12]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rptr[12]_net_1\);
    
    \wptr[2]\ : SLE
      port map(D => \wptr_s[2]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[2]_net_1\);
    
    \rptr_cry[2]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[2]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[1]_net_1\, S
         => \rptr_s[2]\, Y => OPEN, FCO => \rptr_cry[2]_net_1\);
    
    rdiff_bus_cry_9 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[9]_net_1\, B => 
        \rptr[9]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_8\, S => \rdiff_bus[9]\, Y => OPEN, FCO
         => \rdiff_bus_cry_9\);
    
    \memwaddr_r[0]\ : SLE
      port map(D => \fifo_MEMWADDR_i[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[0]\);
    
    \wptr_gray[2]\ : SLE
      port map(D => \wptr_gray_1[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[2]_net_1\);
    
    \wptr_cry[12]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[12]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[11]_net_1\, S
         => \wptr_s[12]\, Y => OPEN, FCO => \wptr_cry[12]_net_1\);
    
    \memwaddr_r_2[7]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_7_S, D => un4_we_i_9, Y => 
        \memwaddr_r_2[7]_net_1\);
    
    wdiff_bus_cry_4 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[4]_net_1\, B => 
        \rptr_bin_sync2[4]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_3\, S => \wdiff_bus[4]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_4\);
    
    un1_memraddr_r_cry_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMRADDR[7]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memraddr_r_cry_6\, 
        S => un1_memraddr_r_cry_7_S, Y => OPEN, FCO => 
        \un1_memraddr_r_cry_7\);
    
    \wptr_s[13]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[13]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[12]_net_1\, S
         => \wptr_s[13]_net_1\, Y => OPEN, FCO => OPEN);
    
    \wptr_gray[11]\ : SLE
      port map(D => \wptr_gray_1[11]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[11]_net_1\);
    
    \wptr_bin_sync2[9]\ : SLE
      port map(D => \wptr_bin_sync[9]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_bin_sync2[9]_net_1\);
    
    \rptr_gray_1[6]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[6]_net_1\, B => \rptr[7]_net_1\, Y => 
        \rptr_gray_1[6]_net_1\);
    
    \wptr_gray_1[10]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[10]_net_1\, B => \wptr[11]_net_1\, Y
         => \wptr_gray_1[10]_net_1\);
    
    wdiff_bus_cry_6 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[6]_net_1\, B => 
        \rptr_bin_sync2[6]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_5\, S => \wdiff_bus[6]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_6\);
    
    \rptr_cry[3]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[3]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[2]_net_1\, S
         => \rptr_s[3]\, Y => OPEN, FCO => \rptr_cry[3]_net_1\);
    
    \memraddr_r[4]\ : SLE
      port map(D => un1_memraddr_r_cry_4_S, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[4]\);
    
    \rptr[13]\ : SLE
      port map(D => \rptr_s[13]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \rptr[13]_net_1\);
    
    \wptr_cry[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \wptr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \wptr_cry[10]_net_1\, S
         => \wptr_s[11]\, Y => OPEN, FCO => \wptr_cry[11]_net_1\);
    
    \memwaddr_r_2[8]\ : CFG4
      generic map(INIT => x"70F0")

      port map(A => un4_we_i_8, B => un4_we_i_7, C => 
        un1_memwaddr_r_cry_8_S, D => un4_we_i_9, Y => 
        \memwaddr_r_2[8]_net_1\);
    
    \memwaddr_r[12]\ : SLE
      port map(D => \memwaddr_r_2[12]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => \fifo_MEMWE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMWADDR[12]\);
    
    \L1.un4_re_i_0\ : CFG2
      generic map(INIT => x"4")

      port map(A => \fifo_MEMRADDR[5]\, B => \fifo_MEMRADDR[12]\, 
        Y => un4_re_i_0);
    
    \rptr_cry[12]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[12]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[11]_net_1\, S
         => \rptr_s[12]\, Y => OPEN, FCO => \rptr_cry[12]_net_1\);
    
    memre_0_a2 : CFG2
      generic map(INIT => x"2")

      port map(A => iRX_FIFO_rd_en_0, B => \iRX_FIFO_Empty_0\, Y
         => \fifo_MEMRE\);
    
    \memraddr_r[11]\ : SLE
      port map(D => \memraddr_r_2[11]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[11]\);
    
    rdiff_bus_cry_12 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[12]_net_1\, B => 
        \rptr[12]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_11\, S => \rdiff_bus[12]\, Y => OPEN, FCO
         => \rdiff_bus_cry_12\);
    
    \memraddr_r[5]\ : SLE
      port map(D => \memraddr_r_2[5]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[5]\);
    
    \rptr_gray[6]\ : SLE
      port map(D => \rptr_gray_1[6]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[6]_net_1\);
    
    \memraddr_r[9]\ : SLE
      port map(D => \memraddr_r_2[9]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[9]\);
    
    \rptr[0]\ : SLE
      port map(D => \rptr_s[0]\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \fifo_MEMRE\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rptr[0]_net_1\);
    
    \wptr[10]\ : SLE
      port map(D => \wptr_s[10]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[10]_net_1\);
    
    \L1.un4_we_i_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => \fifo_MEMWADDR[1]\, B => \fifo_MEMWADDR[2]\, 
        Y => un4_we_i_0);
    
    wdiff_bus_cry_1 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[1]_net_1\, B => 
        \rptr_bin_sync2[1]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_0\, S => \wdiff_bus[1]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_1\);
    
    rdiff_bus_cry_2 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[2]_net_1\, B => 
        \rptr[2]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_1\, S => \rdiff_bus[2]\, Y => OPEN, FCO
         => \rdiff_bus_cry_2\);
    
    \wptr_gray[9]\ : SLE
      port map(D => \wptr_gray_1[9]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[9]_net_1\);
    
    \rptr_gray_1[4]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[4]_net_1\, B => \rptr[5]_net_1\, Y => 
        \rptr_gray_1[4]_net_1\);
    
    \wptr_gray_1[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[8]_net_1\, B => \wptr[9]_net_1\, Y => 
        \wptr_gray_1[8]_net_1\);
    
    Rd_corefifo_grayToBinConv : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_grayToBinConv_1_3
      port map(rptr_bin_sync(13) => \rptr_bin_sync[13]\, 
        rptr_bin_sync(12) => \rptr_bin_sync[12]\, 
        rptr_bin_sync(11) => \rptr_bin_sync[11]\, 
        rptr_bin_sync(10) => \rptr_bin_sync[10]\, 
        rptr_bin_sync(9) => \rptr_bin_sync[9]\, rptr_bin_sync(8)
         => \rptr_bin_sync[8]\, rptr_bin_sync(7) => 
        \rptr_bin_sync[7]\, rptr_bin_sync(6) => nc2, 
        rptr_bin_sync(5) => \rptr_bin_sync[5]\, rptr_bin_sync(4)
         => nc1, rptr_bin_sync(3) => \rptr_bin_sync[3]\, 
        rptr_bin_sync(2) => \rptr_bin_sync[2]\, rptr_bin_sync(1)
         => \rptr_bin_sync[1]\, rptr_bin_sync(0) => 
        \rptr_bin_sync[0]\, rptr_gray_sync(12) => 
        \rptr_gray_sync[12]\, rptr_gray_sync(11) => 
        \rptr_gray_sync[11]\, rptr_gray_sync(10) => 
        \rptr_gray_sync[10]\, rptr_gray_sync(9) => 
        \rptr_gray_sync[9]\, rptr_gray_sync(8) => 
        \rptr_gray_sync[8]\, rptr_gray_sync(7) => 
        \rptr_gray_sync[7]\, rptr_gray_sync(6) => 
        \rptr_gray_sync[6]\, rptr_gray_sync(5) => 
        \rptr_gray_sync[5]\, rptr_gray_sync(4) => 
        \rptr_gray_sync[4]\, rptr_gray_sync(3) => 
        \rptr_gray_sync[3]\, rptr_gray_sync(2) => 
        \rptr_gray_sync[2]\, rptr_gray_sync(1) => 
        \rptr_gray_sync[1]\, rptr_gray_sync(0) => 
        \rptr_gray_sync[0]\, bin_N_6_i => bin_N_6_i, bin_N_4_0_i
         => bin_N_4_0_i);
    
    \rptr_cry[1]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[1]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => rptr_s_908_FCO, S => 
        \rptr_s[1]\, Y => OPEN, FCO => \rptr_cry[1]_net_1\);
    
    \rptr_cry[11]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[11]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[10]_net_1\, S
         => \rptr_s[11]\, Y => OPEN, FCO => \rptr_cry[11]_net_1\);
    
    rdiff_bus_cry_3 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[3]_net_1\, B => 
        \rptr[3]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_2\, S => \rdiff_bus[3]\, Y => OPEN, FCO
         => \rdiff_bus_cry_3\);
    
    rdiff_bus_cry_10 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr_bin_sync2[10]_net_1\, B => 
        \rptr[10]_net_1\, C => GND_net_1, D => GND_net_1, FCI => 
        \rdiff_bus_cry_9\, S => \rdiff_bus[10]\, Y => OPEN, FCO
         => \rdiff_bus_cry_10\);
    
    un1_memwaddr_r_cry_11 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[11]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_10\, 
        S => un1_memwaddr_r_cry_11_S, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_11\);
    
    \memraddr_r[6]\ : SLE
      port map(D => un1_memraddr_r_cry_6_S, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[6]\);
    
    \rptr_cry[7]\ : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \rptr[7]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => \rptr_cry[6]_net_1\, S
         => \rptr_s[7]\, Y => OPEN, FCO => \rptr_cry[7]_net_1\);
    
    rdiff_bus_cry_0 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => rdiff_bus, B => \rptr[0]_net_1\, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => rdiff_bus_cry_0_Y_0, FCO => \rdiff_bus_cry_0\);
    
    \memraddr_r[2]\ : SLE
      port map(D => un1_memraddr_r_cry_2_S, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[2]\);
    
    \wptr[8]\ : SLE
      port map(D => \wptr_s[8]\, CLK => CommsFPGA_CCC_0_GL0, EN
         => \fifo_MEMWE\, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \wptr[8]_net_1\);
    
    wdiff_bus_cry_3 : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \wptr[3]_net_1\, B => 
        \rptr_bin_sync2[3]_net_1\, C => GND_net_1, D => GND_net_1, 
        FCI => \wdiff_bus_cry_2\, S => \wdiff_bus[3]\, Y => OPEN, 
        FCO => \wdiff_bus_cry_3\);
    
    rdiff_bus_s_13 : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \rptr[13]_net_1\, C => 
        \wptr_bin_sync2[13]_net_1\, D => GND_net_1, FCI => 
        \rdiff_bus_cry_12\, S => \rdiff_bus[13]\, Y => OPEN, FCO
         => OPEN);
    
    \memraddr_r[12]\ : SLE
      port map(D => \memraddr_r_2[12]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \fifo_MEMRE\, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \fifo_MEMRADDR[12]\);
    
    \wptr_gray_1[11]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \wptr[11]_net_1\, B => \wptr[12]_net_1\, Y
         => \wptr_gray_1[11]_net_1\);
    
    \rptr_gray[7]\ : SLE
      port map(D => \rptr_gray_1[7]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rptr_gray[7]_net_1\);
    
    \wptr_gray[0]\ : SLE
      port map(D => \wptr_gray_1[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \wptr_gray[0]_net_1\);
    
    \rptr_gray_1[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[0]_net_1\, B => \rptr[1]_net_1\, Y => 
        \rptr_gray_1[0]_net_1\);
    
    un1_memwaddr_r_cry_10 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \fifo_MEMWADDR[10]\, C => 
        GND_net_1, D => GND_net_1, FCI => \un1_memwaddr_r_cry_9\, 
        S => un1_memwaddr_r_cry_10_S, Y => OPEN, FCO => 
        \un1_memwaddr_r_cry_10\);
    
    \rptr_gray_1[8]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \rptr[8]_net_1\, B => \rptr[9]_net_1\, Y => 
        \rptr_gray_1[8]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO is

    port( RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          RX_FIFO_DOUT_0            : out   std_logic_vector(8 downto 0);
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_wr_en_0_0        : in    std_logic;
          iRX_FIFO_rd_en_0          : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic;
          RX_FIFO_TxColDetDis_wr_en : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          irx_fifo_rst_i            : in    std_logic
        );

end FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO;

architecture DEF_ARCH of FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO is 

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper
    port( fifo_MEMRADDR             : in    std_logic_vector(12 downto 0) := (others => 'U');
          fifo_MEMWADDR             : in    std_logic_vector(12 downto 0) := (others => 'U');
          RDATA_int                 : out   std_logic_vector(8 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          fifo_MEMRE                : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          fifo_MEMWE                : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3
    port( fifo_MEMRADDR             : out   std_logic_vector(12 downto 0);
          fifo_MEMWADDR             : out   std_logic_vector(12 downto 0);
          iRX_FIFO_wr_en_0_0        : in    std_logic := 'U';
          iRX_FIFO_rd_en_0          : in    std_logic := 'U';
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          RX_FIFO_TxColDetDis_wr_en : in    std_logic := 'U';
          fifo_MEMRE                : out   std_logic;
          fifo_MEMWE                : out   std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          irx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \RDATA_r[0]_net_1\, VCC_net_1, \RDATA_int[0]\, 
        \un6_fifo_memre\, GND_net_1, \RDATA_r[1]_net_1\, 
        \RDATA_int[1]\, \RDATA_r[2]_net_1\, \RDATA_int[2]\, 
        \RDATA_r[3]_net_1\, \RDATA_int[3]\, \RDATA_r[4]_net_1\, 
        \RDATA_int[4]\, \RDATA_r[5]_net_1\, \RDATA_int[5]\, 
        \RDATA_r[6]_net_1\, \RDATA_int[6]\, \RDATA_r[7]_net_1\, 
        \RDATA_int[7]\, \RDATA_r[8]_net_1\, \RDATA_int[8]\, 
        \re_set\, \REN_d1\, \un9_fifo_memre\, fifo_MEMRE, \RE_d1\, 
        \re_pulse_d1\, \re_pulse\, \fifo_MEMRADDR[0]\, 
        \fifo_MEMRADDR[1]\, \fifo_MEMRADDR[2]\, 
        \fifo_MEMRADDR[3]\, \fifo_MEMRADDR[4]\, 
        \fifo_MEMRADDR[5]\, \fifo_MEMRADDR[6]\, 
        \fifo_MEMRADDR[7]\, \fifo_MEMRADDR[8]\, 
        \fifo_MEMRADDR[9]\, \fifo_MEMRADDR[10]\, 
        \fifo_MEMRADDR[11]\, \fifo_MEMRADDR[12]\, 
        \fifo_MEMWADDR[0]\, \fifo_MEMWADDR[1]\, 
        \fifo_MEMWADDR[2]\, \fifo_MEMWADDR[3]\, 
        \fifo_MEMWADDR[4]\, \fifo_MEMWADDR[5]\, 
        \fifo_MEMWADDR[6]\, \fifo_MEMWADDR[7]\, 
        \fifo_MEMWADDR[8]\, \fifo_MEMWADDR[9]\, 
        \fifo_MEMWADDR[10]\, \fifo_MEMWADDR[11]\, 
        \fifo_MEMWADDR[12]\, fifo_MEMWE : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper(DEF_ARCH);
    for all : FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3(DEF_ARCH);
begin 


    re_pulse : CFG3
      generic map(INIT => x"DC")

      port map(A => fifo_MEMRE, B => \re_set\, C => \REN_d1\, Y
         => \re_pulse\);
    
    \RDATA_r[3]\ : SLE
      port map(D => \RDATA_int[3]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \un6_fifo_memre\, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[3]_net_1\);
    
    \Q[6]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[6]_net_1\, C => 
        \RDATA_int[6]\, D => \RE_d1\, Y => RX_FIFO_DOUT_0(6));
    
    re_pulse_d1 : SLE
      port map(D => \re_pulse\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \re_pulse_d1\);
    
    \RDATA_r[5]\ : SLE
      port map(D => \RDATA_int[5]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \un6_fifo_memre\, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[5]_net_1\);
    
    un9_fifo_memre : CFG2
      generic map(INIT => x"6")

      port map(A => fifo_MEMRE, B => \REN_d1\, Y => 
        \un9_fifo_memre\);
    
    \RDATA_r[8]\ : SLE
      port map(D => \RDATA_int[8]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \un6_fifo_memre\, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[8]_net_1\);
    
    \Q[2]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[2]_net_1\, C => 
        \RDATA_int[2]\, D => \RE_d1\, Y => RX_FIFO_DOUT_0(2));
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \RW1.UI_ram_wrapper_1\ : FIFO_8Kx9_FIFO_8Kx9_0_ram_wrapper
      port map(fifo_MEMRADDR(12) => \fifo_MEMRADDR[12]\, 
        fifo_MEMRADDR(11) => \fifo_MEMRADDR[11]\, 
        fifo_MEMRADDR(10) => \fifo_MEMRADDR[10]\, 
        fifo_MEMRADDR(9) => \fifo_MEMRADDR[9]\, fifo_MEMRADDR(8)
         => \fifo_MEMRADDR[8]\, fifo_MEMRADDR(7) => 
        \fifo_MEMRADDR[7]\, fifo_MEMRADDR(6) => 
        \fifo_MEMRADDR[6]\, fifo_MEMRADDR(5) => 
        \fifo_MEMRADDR[5]\, fifo_MEMRADDR(4) => 
        \fifo_MEMRADDR[4]\, fifo_MEMRADDR(3) => 
        \fifo_MEMRADDR[3]\, fifo_MEMRADDR(2) => 
        \fifo_MEMRADDR[2]\, fifo_MEMRADDR(1) => 
        \fifo_MEMRADDR[1]\, fifo_MEMRADDR(0) => 
        \fifo_MEMRADDR[0]\, fifo_MEMWADDR(12) => 
        \fifo_MEMWADDR[12]\, fifo_MEMWADDR(11) => 
        \fifo_MEMWADDR[11]\, fifo_MEMWADDR(10) => 
        \fifo_MEMWADDR[10]\, fifo_MEMWADDR(9) => 
        \fifo_MEMWADDR[9]\, fifo_MEMWADDR(8) => 
        \fifo_MEMWADDR[8]\, fifo_MEMWADDR(7) => 
        \fifo_MEMWADDR[7]\, fifo_MEMWADDR(6) => 
        \fifo_MEMWADDR[6]\, fifo_MEMWADDR(5) => 
        \fifo_MEMWADDR[5]\, fifo_MEMWADDR(4) => 
        \fifo_MEMWADDR[4]\, fifo_MEMWADDR(3) => 
        \fifo_MEMWADDR[3]\, fifo_MEMWADDR(2) => 
        \fifo_MEMWADDR[2]\, fifo_MEMWADDR(1) => 
        \fifo_MEMWADDR[1]\, fifo_MEMWADDR(0) => 
        \fifo_MEMWADDR[0]\, RDATA_int(8) => \RDATA_int[8]\, 
        RDATA_int(7) => \RDATA_int[7]\, RDATA_int(6) => 
        \RDATA_int[6]\, RDATA_int(5) => \RDATA_int[5]\, 
        RDATA_int(4) => \RDATA_int[4]\, RDATA_int(3) => 
        \RDATA_int[3]\, RDATA_int(2) => \RDATA_int[2]\, 
        RDATA_int(1) => \RDATA_int[1]\, RDATA_int(0) => 
        \RDATA_int[0]\, RX_FIFO_DIN_pipe(8) => 
        RX_FIFO_DIN_pipe(8), RX_FIFO_DIN_pipe(7) => 
        RX_FIFO_DIN_pipe(7), RX_FIFO_DIN_pipe(6) => 
        RX_FIFO_DIN_pipe(6), RX_FIFO_DIN_pipe(5) => 
        RX_FIFO_DIN_pipe(5), RX_FIFO_DIN_pipe(4) => 
        RX_FIFO_DIN_pipe(4), RX_FIFO_DIN_pipe(3) => 
        RX_FIFO_DIN_pipe(3), RX_FIFO_DIN_pipe(2) => 
        RX_FIFO_DIN_pipe(2), RX_FIFO_DIN_pipe(1) => 
        RX_FIFO_DIN_pipe(1), RX_FIFO_DIN_pipe(0) => 
        RX_FIFO_DIN_pipe(0), m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, fifo_MEMRE => fifo_MEMRE, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, fifo_MEMWE
         => fifo_MEMWE);
    
    \RDATA_r[0]\ : SLE
      port map(D => \RDATA_int[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \un6_fifo_memre\, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[0]_net_1\);
    
    \Q[4]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[4]_net_1\, C => 
        \RDATA_int[4]\, D => \RE_d1\, Y => RX_FIFO_DOUT_0(4));
    
    \RDATA_r[2]\ : SLE
      port map(D => \RDATA_int[2]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \un6_fifo_memre\, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[2]_net_1\);
    
    \RDATA_r[6]\ : SLE
      port map(D => \RDATA_int[6]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \un6_fifo_memre\, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[6]_net_1\);
    
    \L31.U_corefifo_async\ : 
        FIFO_8Kx9_FIFO_8Kx9_0_corefifo_async_3
      port map(fifo_MEMRADDR(12) => \fifo_MEMRADDR[12]\, 
        fifo_MEMRADDR(11) => \fifo_MEMRADDR[11]\, 
        fifo_MEMRADDR(10) => \fifo_MEMRADDR[10]\, 
        fifo_MEMRADDR(9) => \fifo_MEMRADDR[9]\, fifo_MEMRADDR(8)
         => \fifo_MEMRADDR[8]\, fifo_MEMRADDR(7) => 
        \fifo_MEMRADDR[7]\, fifo_MEMRADDR(6) => 
        \fifo_MEMRADDR[6]\, fifo_MEMRADDR(5) => 
        \fifo_MEMRADDR[5]\, fifo_MEMRADDR(4) => 
        \fifo_MEMRADDR[4]\, fifo_MEMRADDR(3) => 
        \fifo_MEMRADDR[3]\, fifo_MEMRADDR(2) => 
        \fifo_MEMRADDR[2]\, fifo_MEMRADDR(1) => 
        \fifo_MEMRADDR[1]\, fifo_MEMRADDR(0) => 
        \fifo_MEMRADDR[0]\, fifo_MEMWADDR(12) => 
        \fifo_MEMWADDR[12]\, fifo_MEMWADDR(11) => 
        \fifo_MEMWADDR[11]\, fifo_MEMWADDR(10) => 
        \fifo_MEMWADDR[10]\, fifo_MEMWADDR(9) => 
        \fifo_MEMWADDR[9]\, fifo_MEMWADDR(8) => 
        \fifo_MEMWADDR[8]\, fifo_MEMWADDR(7) => 
        \fifo_MEMWADDR[7]\, fifo_MEMWADDR(6) => 
        \fifo_MEMWADDR[6]\, fifo_MEMWADDR(5) => 
        \fifo_MEMWADDR[5]\, fifo_MEMWADDR(4) => 
        \fifo_MEMWADDR[4]\, fifo_MEMWADDR(3) => 
        \fifo_MEMWADDR[3]\, fifo_MEMWADDR(2) => 
        \fifo_MEMWADDR[2]\, fifo_MEMWADDR(1) => 
        \fifo_MEMWADDR[1]\, fifo_MEMWADDR(0) => 
        \fifo_MEMWADDR[0]\, iRX_FIFO_wr_en_0_0 => 
        iRX_FIFO_wr_en_0_0, iRX_FIFO_rd_en_0 => iRX_FIFO_rd_en_0, 
        iRX_FIFO_Empty_0 => iRX_FIFO_Empty_0, iRX_FIFO_UNDERRUN_0
         => iRX_FIFO_UNDERRUN_0, iRX_FIFO_OVERFLOW_0 => 
        iRX_FIFO_OVERFLOW_0, iRX_FIFO_Full_0 => iRX_FIFO_Full_0, 
        RX_FIFO_TxColDetDis_wr_en => RX_FIFO_TxColDetDis_wr_en, 
        fifo_MEMRE => fifo_MEMRE, fifo_MEMWE => fifo_MEMWE, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz, 
        irx_fifo_rst_i => irx_fifo_rst_i);
    
    re_set : SLE
      port map(D => \REN_d1\, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \un9_fifo_memre\, ALn => irx_fifo_rst_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \re_set\);
    
    \Q[3]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[3]_net_1\, C => 
        \RDATA_int[3]\, D => \RE_d1\, Y => RX_FIFO_DOUT_0(3));
    
    \Q[7]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[7]_net_1\, C => 
        \RDATA_int[7]\, D => \RE_d1\, Y => RX_FIFO_DOUT_0(7));
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \Q[8]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[8]_net_1\, C => 
        \RDATA_int[8]\, D => \RE_d1\, Y => RX_FIFO_DOUT_0(8));
    
    RE_d1 : SLE
      port map(D => iRX_FIFO_rd_en_0, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => \RE_d1\);
    
    \RDATA_r[7]\ : SLE
      port map(D => \RDATA_int[7]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \un6_fifo_memre\, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[7]_net_1\);
    
    \RDATA_r[4]\ : SLE
      port map(D => \RDATA_int[4]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \un6_fifo_memre\, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[4]_net_1\);
    
    \Q[1]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[1]_net_1\, C => 
        \RDATA_int[1]\, D => \RE_d1\, Y => RX_FIFO_DOUT_0(1));
    
    \Q[0]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[0]_net_1\, C => 
        \RDATA_int[0]\, D => \RE_d1\, Y => RX_FIFO_DOUT_0(0));
    
    REN_d1 : SLE
      port map(D => fifo_MEMRE, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => irx_fifo_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \REN_d1\);
    
    \Q[5]\ : CFG4
      generic map(INIT => x"F0D8")

      port map(A => \re_pulse_d1\, B => \RDATA_r[5]_net_1\, C => 
        \RDATA_int[5]\, D => \RE_d1\, Y => RX_FIFO_DOUT_0(5));
    
    un6_fifo_memre : CFG2
      generic map(INIT => x"4")

      port map(A => fifo_MEMRE, B => \REN_d1\, Y => 
        \un6_fifo_memre\);
    
    \RDATA_r[1]\ : SLE
      port map(D => \RDATA_int[1]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \un6_fifo_memre\, ALn
         => irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \RDATA_r[1]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFO_8Kx9 is

    port( RX_FIFO_DOUT_0            : out   std_logic_vector(8 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0);
          iRX_FIFO_rd_en_0          : in    std_logic;
          iRX_FIFO_wr_en_0_0        : in    std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          irx_fifo_rst_i            : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz : in    std_logic;
          RX_FIFO_TxColDetDis_wr_en : in    std_logic;
          CommsFPGA_CCC_0_GL0       : in    std_logic
        );

end FIFO_8Kx9;

architecture DEF_ARCH of FIFO_8Kx9 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO
    port( RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          RX_FIFO_DOUT_0            : out   std_logic_vector(8 downto 0);
          iRX_FIFO_Full_0           : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_wr_en_0_0        : in    std_logic := 'U';
          iRX_FIFO_rd_en_0          : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U';
          RX_FIFO_TxColDetDis_wr_en : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          irx_fifo_rst_i            : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal GND_net_1, VCC_net_1 : std_logic;

    for all : FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO
	Use entity work.FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO(DEF_ARCH);
begin 


    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    FIFO_8Kx9_0 : FIFO_8Kx9_FIFO_8Kx9_0_COREFIFO
      port map(RX_FIFO_DIN_pipe(8) => RX_FIFO_DIN_pipe(8), 
        RX_FIFO_DIN_pipe(7) => RX_FIFO_DIN_pipe(7), 
        RX_FIFO_DIN_pipe(6) => RX_FIFO_DIN_pipe(6), 
        RX_FIFO_DIN_pipe(5) => RX_FIFO_DIN_pipe(5), 
        RX_FIFO_DIN_pipe(4) => RX_FIFO_DIN_pipe(4), 
        RX_FIFO_DIN_pipe(3) => RX_FIFO_DIN_pipe(3), 
        RX_FIFO_DIN_pipe(2) => RX_FIFO_DIN_pipe(2), 
        RX_FIFO_DIN_pipe(1) => RX_FIFO_DIN_pipe(1), 
        RX_FIFO_DIN_pipe(0) => RX_FIFO_DIN_pipe(0), 
        RX_FIFO_DOUT_0(8) => RX_FIFO_DOUT_0(8), RX_FIFO_DOUT_0(7)
         => RX_FIFO_DOUT_0(7), RX_FIFO_DOUT_0(6) => 
        RX_FIFO_DOUT_0(6), RX_FIFO_DOUT_0(5) => RX_FIFO_DOUT_0(5), 
        RX_FIFO_DOUT_0(4) => RX_FIFO_DOUT_0(4), RX_FIFO_DOUT_0(3)
         => RX_FIFO_DOUT_0(3), RX_FIFO_DOUT_0(2) => 
        RX_FIFO_DOUT_0(2), RX_FIFO_DOUT_0(1) => RX_FIFO_DOUT_0(1), 
        RX_FIFO_DOUT_0(0) => RX_FIFO_DOUT_0(0), iRX_FIFO_Full_0
         => iRX_FIFO_Full_0, iRX_FIFO_OVERFLOW_0 => 
        iRX_FIFO_OVERFLOW_0, iRX_FIFO_UNDERRUN_0 => 
        iRX_FIFO_UNDERRUN_0, iRX_FIFO_Empty_0 => iRX_FIFO_Empty_0, 
        iRX_FIFO_wr_en_0_0 => iRX_FIFO_wr_en_0_0, 
        iRX_FIFO_rd_en_0 => iRX_FIFO_rd_en_0, CommsFPGA_CCC_0_GL0
         => CommsFPGA_CCC_0_GL0, RX_FIFO_TxColDetDis_wr_en => 
        RX_FIFO_TxColDetDis_wr_en, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, irx_fifo_rst_i => 
        irx_fifo_rst_i);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity FIFOs is

    port( RX_FIFO_DIN_pipe             : in    std_logic_vector(8 downto 0);
          CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0);
          TX_FIFO_DOUT                 : out   std_logic_vector(7 downto 0);
          up_EOP_sync                  : in    std_logic_vector(2 downto 1);
          RX_FIFO_DOUT                 : out   std_logic_vector(8 downto 0);
          iRX_FIFO_Full                : out   std_logic_vector(3 downto 0);
          iRX_FIFO_UNDERRUN            : out   std_logic_vector(3 downto 0);
          iRX_FIFO_Empty               : out   std_logic_vector(3 downto 0);
          ReadFIFO_Write_Ptr           : out   std_logic_vector(1 downto 0);
          ReadFIFO_Read_Ptr            : out   std_logic_vector(1 downto 0);
          packet_available_clear_reg   : out   std_logic_vector(2 downto 0);
          RX_FIFO_TxColDetDis_wr_en    : in    std_logic;
          TX_FIFO_UNDERRUN             : out   std_logic;
          TX_FIFO_UNDERRUN_i           : out   std_logic;
          TX_FIFO_OVERFLOW             : out   std_logic;
          TX_FIFO_OVERFLOW_i           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic;
          TX_FIFO_Full                 : out   std_logic;
          TX_FIFO_wr_en                : in    std_logic;
          TX_FIFO_Empty                : out   std_logic;
          N_114                        : in    std_logic;
          BIT_CLK                      : in    std_logic;
          RX_FIFO_RST                  : in    std_logic;
          TX_FIFO_RST                  : in    std_logic;
          RESET                        : in    std_logic;
          RX_FIFO_rd_en                : in    std_logic;
          rx_packet_complt             : in    std_logic;
          RX_FIFO_Full                 : out   std_logic;
          RX_FIFO_Empty                : out   std_logic;
          rx_packet_avail_int          : in    std_logic;
          CommsFPGA_CCC_0_GL0          : in    std_logic;
          RX_FIFO_OVERFLOW_i           : out   std_logic;
          RX_FIFO_OVERFLOW             : out   std_logic;
          RX_FIFO_UNDERRUN_i           : out   std_logic;
          RX_FIFO_UNDERRUN             : out   std_logic
        );

end FIFOs;

architecture DEF_ARCH of FIFOs is 

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component FIFO_2Kx8
    port( TX_FIFO_DOUT                 : out   std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0) := (others => 'U');
          itx_fifo_rst_i               : in    std_logic := 'U';
          BIT_CLK                      : in    std_logic := 'U';
          N_114                        : in    std_logic := 'U';
          TX_FIFO_Empty                : out   std_logic;
          TX_FIFO_wr_en                : in    std_logic := 'U';
          TX_FIFO_Full                 : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic := 'U';
          TX_FIFO_OVERFLOW_i           : out   std_logic;
          TX_FIFO_OVERFLOW             : out   std_logic;
          TX_FIFO_UNDERRUN_i           : out   std_logic;
          TX_FIFO_UNDERRUN             : out   std_logic
        );
  end component;

  component FIFO_8Kx9_0
    port( RX_FIFO_DOUT_1            : out   std_logic_vector(8 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          iRX_FIFO_rd_en_0          : in    std_logic := 'U';
          iRX_FIFO_wr_en_0_0        : in    std_logic := 'U';
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          irx_fifo_rst_i            : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          RX_FIFO_TxColDetDis_wr_en : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9_1
    port( RX_FIFO_DOUT_2            : out   std_logic_vector(8 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          iRX_FIFO_rd_en_0          : in    std_logic := 'U';
          iRX_FIFO_wr_en_0_0        : in    std_logic := 'U';
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          irx_fifo_rst_i            : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          RX_FIFO_TxColDetDis_wr_en : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component FIFO_8Kx9_2
    port( RX_FIFO_DOUT_3            : out   std_logic_vector(8 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          iRX_FIFO_rd_en_0          : in    std_logic := 'U';
          iRX_FIFO_wr_en_0_0        : in    std_logic := 'U';
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          irx_fifo_rst_i            : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          RX_FIFO_TxColDetDis_wr_en : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U'
        );
  end component;

  component FIFO_8Kx9
    port( RX_FIFO_DOUT_0            : out   std_logic_vector(8 downto 0);
          RX_FIFO_DIN_pipe          : in    std_logic_vector(8 downto 0) := (others => 'U');
          iRX_FIFO_rd_en_0          : in    std_logic := 'U';
          iRX_FIFO_wr_en_0_0        : in    std_logic := 'U';
          iRX_FIFO_Empty_0          : out   std_logic;
          iRX_FIFO_UNDERRUN_0       : out   std_logic;
          iRX_FIFO_OVERFLOW_0       : out   std_logic;
          iRX_FIFO_Full_0           : out   std_logic;
          irx_fifo_rst_i            : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz : in    std_logic := 'U';
          RX_FIFO_TxColDetDis_wr_en : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0       : in    std_logic := 'U'
        );
  end component;

    signal itx_fifo_rst_i, \itx_fifo_rst\, irx_fifo_rst_i, 
        \irx_fifo_rst\, \RX_FIFO_UNDERRUN\, \RX_FIFO_OVERFLOW\, 
        \packet_available_clear_reg[0]_net_1\, VCC_net_1, 
        GND_net_1, \packet_available_clear_reg[1]_net_1\, 
        \ReadFIFO_Read_Ptr[0]_net_1\, \ReadFIFO_Read_Ptr_2[0]\, 
        \ReadFIFO_Read_Ptr[1]_net_1\, \ReadFIFO_Read_Ptr_2[1]\, 
        \ReadFIFO_Write_Ptr[0]_net_1\, \ReadFIFO_Write_Ptr_3[0]\, 
        \ReadFIFO_Write_Ptr[1]_net_1\, \ReadFIFO_Write_Ptr_3[1]\, 
        \iRX_FIFO_Empty[2]\, \iRX_FIFO_Empty[3]\, 
        RX_FIFO_Empty_3_0_0_y0, RX_FIFO_Empty_3_0_0_co0, 
        \iRX_FIFO_Empty[0]\, \iRX_FIFO_Empty[1]\, 
        \iRX_FIFO_UNDERRUN[2]\, \iRX_FIFO_UNDERRUN[3]\, 
        RX_FIFO_UNDERRUN_3_0_0_y0, RX_FIFO_UNDERRUN_3_0_0_co0, 
        \iRX_FIFO_UNDERRUN[0]\, \iRX_FIFO_UNDERRUN[1]\, 
        \iRX_FIFO_OVERFLOW[2]\, \iRX_FIFO_OVERFLOW[3]\, 
        RX_FIFO_OVERFLOW_3_0_0_y0, RX_FIFO_OVERFLOW_3_0_0_co0, 
        \iRX_FIFO_OVERFLOW[0]\, \iRX_FIFO_OVERFLOW[1]\, 
        \iRX_FIFO_Full[2]\, \iRX_FIFO_Full[3]\, 
        RX_FIFO_Full_3_0_0_y0, RX_FIFO_Full_3_0_0_co0, 
        \iRX_FIFO_Full[0]\, \iRX_FIFO_Full[1]\, 
        \RX_FIFO_DOUT_2[2]\, \RX_FIFO_DOUT_3[2]\, 
        \RX_FIFO_DOUT_3_0_0_y0[2]\, \RX_FIFO_DOUT_3_0_0_co0[2]\, 
        \RX_FIFO_DOUT_0[2]\, \RX_FIFO_DOUT_1[2]\, 
        \RX_FIFO_DOUT_2[8]\, \RX_FIFO_DOUT_3[8]\, 
        \RX_FIFO_DOUT_3_0_0_y0[8]\, \RX_FIFO_DOUT_3_0_0_co0[8]\, 
        \RX_FIFO_DOUT_0[8]\, \RX_FIFO_DOUT_1[8]\, 
        \RX_FIFO_DOUT_2[6]\, \RX_FIFO_DOUT_3[6]\, 
        \RX_FIFO_DOUT_3_0_0_y0[6]\, \RX_FIFO_DOUT_3_0_0_co0[6]\, 
        \RX_FIFO_DOUT_0[6]\, \RX_FIFO_DOUT_1[6]\, 
        \RX_FIFO_DOUT_2[5]\, \RX_FIFO_DOUT_3[5]\, 
        \RX_FIFO_DOUT_3_0_0_y0[5]\, \RX_FIFO_DOUT_3_0_0_co0[5]\, 
        \RX_FIFO_DOUT_0[5]\, \RX_FIFO_DOUT_1[5]\, 
        \RX_FIFO_DOUT_2[4]\, \RX_FIFO_DOUT_3[4]\, 
        \RX_FIFO_DOUT_3_0_0_y0[4]\, \RX_FIFO_DOUT_3_0_0_co0[4]\, 
        \RX_FIFO_DOUT_0[4]\, \RX_FIFO_DOUT_1[4]\, 
        \RX_FIFO_DOUT_2[1]\, \RX_FIFO_DOUT_3[1]\, 
        \RX_FIFO_DOUT_3_0_0_y0[1]\, \RX_FIFO_DOUT_3_0_0_co0[1]\, 
        \RX_FIFO_DOUT_0[1]\, \RX_FIFO_DOUT_1[1]\, 
        \RX_FIFO_DOUT_2[0]\, \RX_FIFO_DOUT_3[0]\, 
        \RX_FIFO_DOUT_3_0_0_y0[0]\, \RX_FIFO_DOUT_3_0_0_co0[0]\, 
        \RX_FIFO_DOUT_0[0]\, \RX_FIFO_DOUT_1[0]\, 
        \RX_FIFO_DOUT_2[7]\, \RX_FIFO_DOUT_3[7]\, 
        \RX_FIFO_DOUT_3_0_0_y0[7]\, \RX_FIFO_DOUT_3_0_0_co0[7]\, 
        \RX_FIFO_DOUT_0[7]\, \RX_FIFO_DOUT_1[7]\, 
        \RX_FIFO_DOUT_2[3]\, \RX_FIFO_DOUT_3[3]\, 
        \RX_FIFO_DOUT_3_0_0_y0[3]\, \RX_FIFO_DOUT_3_0_0_co0[3]\, 
        \RX_FIFO_DOUT_0[3]\, \RX_FIFO_DOUT_1[3]\, 
        \iRX_FIFO_wr_en_0[1]\, \iRX_FIFO_wr_en_0[0]\, 
        \iRX_FIFO_wr_en_0[2]\, \iRX_FIFO_wr_en_0[3]\, 
        \iRX_FIFO_rd_en[2]\, \iRX_FIFO_rd_en[0]\, 
        \iRX_FIFO_rd_en[3]\, \iRX_FIFO_rd_en[1]\ : std_logic;

    for all : FIFO_2Kx8
	Use entity work.FIFO_2Kx8(DEF_ARCH);
    for all : FIFO_8Kx9_0
	Use entity work.FIFO_8Kx9_0(DEF_ARCH);
    for all : FIFO_8Kx9_1
	Use entity work.FIFO_8Kx9_1(DEF_ARCH);
    for all : FIFO_8Kx9_2
	Use entity work.FIFO_8Kx9_2(DEF_ARCH);
    for all : FIFO_8Kx9
	Use entity work.FIFO_8Kx9(DEF_ARCH);
begin 

    iRX_FIFO_Full(3) <= \iRX_FIFO_Full[3]\;
    iRX_FIFO_Full(2) <= \iRX_FIFO_Full[2]\;
    iRX_FIFO_Full(1) <= \iRX_FIFO_Full[1]\;
    iRX_FIFO_Full(0) <= \iRX_FIFO_Full[0]\;
    iRX_FIFO_UNDERRUN(3) <= \iRX_FIFO_UNDERRUN[3]\;
    iRX_FIFO_UNDERRUN(2) <= \iRX_FIFO_UNDERRUN[2]\;
    iRX_FIFO_UNDERRUN(1) <= \iRX_FIFO_UNDERRUN[1]\;
    iRX_FIFO_UNDERRUN(0) <= \iRX_FIFO_UNDERRUN[0]\;
    iRX_FIFO_Empty(3) <= \iRX_FIFO_Empty[3]\;
    iRX_FIFO_Empty(2) <= \iRX_FIFO_Empty[2]\;
    iRX_FIFO_Empty(1) <= \iRX_FIFO_Empty[1]\;
    iRX_FIFO_Empty(0) <= \iRX_FIFO_Empty[0]\;
    ReadFIFO_Write_Ptr(1) <= \ReadFIFO_Write_Ptr[1]_net_1\;
    ReadFIFO_Write_Ptr(0) <= \ReadFIFO_Write_Ptr[0]_net_1\;
    ReadFIFO_Read_Ptr(1) <= \ReadFIFO_Read_Ptr[1]_net_1\;
    ReadFIFO_Read_Ptr(0) <= \ReadFIFO_Read_Ptr[0]_net_1\;
    packet_available_clear_reg(1) <= 
        \packet_available_clear_reg[1]_net_1\;
    packet_available_clear_reg(0) <= 
        \packet_available_clear_reg[0]_net_1\;
    RX_FIFO_OVERFLOW <= \RX_FIFO_OVERFLOW\;
    RX_FIFO_UNDERRUN <= \RX_FIFO_UNDERRUN\;

    RX_FIFO_Full_3_0_0_wmux : ARI1
      generic map(INIT => x"0FA44")

      port map(A => \ReadFIFO_Read_Ptr[0]_net_1\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \iRX_FIFO_Full[0]\, D
         => \iRX_FIFO_Full[1]\, FCI => VCC_net_1, S => OPEN, Y
         => RX_FIFO_Full_3_0_0_y0, FCO => RX_FIFO_Full_3_0_0_co0);
    
    \RX_FIFO_DOUT_3_0_0_wmux_0[6]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \RX_FIFO_DOUT_3_0_0_y0[6]\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \RX_FIFO_DOUT_2[6]\, D
         => \RX_FIFO_DOUT_3[6]\, FCI => 
        \RX_FIFO_DOUT_3_0_0_co0[6]\, S => OPEN, Y => 
        RX_FIFO_DOUT(6), FCO => OPEN);
    
    irx_fifo_rst_RNIS228 : CLKINT
      port map(A => \irx_fifo_rst\, Y => irx_fifo_rst_i);
    
    \RX_FIFO_DOUT_3_0_0_wmux[6]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => \ReadFIFO_Read_Ptr[0]_net_1\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \RX_FIFO_DOUT_0[6]\, D
         => \RX_FIFO_DOUT_1[6]\, FCI => VCC_net_1, S => OPEN, Y
         => \RX_FIFO_DOUT_3_0_0_y0[6]\, FCO => 
        \RX_FIFO_DOUT_3_0_0_co0[6]\);
    
    \ReadFIFO_Read_Ptr_RNO[1]\ : CFG4
      generic map(INIT => x"B4F0")

      port map(A => up_EOP_sync(1), B => up_EOP_sync(2), C => 
        \ReadFIFO_Read_Ptr[1]_net_1\, D => 
        \ReadFIFO_Read_Ptr[0]_net_1\, Y => 
        \ReadFIFO_Read_Ptr_2[1]\);
    
    RX_FIFO_UNDERRUN_3_0_0_wmux : ARI1
      generic map(INIT => x"0FA44")

      port map(A => \ReadFIFO_Read_Ptr[0]_net_1\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \iRX_FIFO_UNDERRUN[0]\, 
        D => \iRX_FIFO_UNDERRUN[1]\, FCI => VCC_net_1, S => OPEN, 
        Y => RX_FIFO_UNDERRUN_3_0_0_y0, FCO => 
        RX_FIFO_UNDERRUN_3_0_0_co0);
    
    RX_FIFO_Empty_3_0_0_wmux : ARI1
      generic map(INIT => x"0FA44")

      port map(A => \ReadFIFO_Read_Ptr[0]_net_1\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \iRX_FIFO_Empty[0]\, D
         => \iRX_FIFO_Empty[1]\, FCI => VCC_net_1, S => OPEN, Y
         => RX_FIFO_Empty_3_0_0_y0, FCO => 
        RX_FIFO_Empty_3_0_0_co0);
    
    RX_FIFO_OVERFLOW_3_0_0_wmux : ARI1
      generic map(INIT => x"0FA44")

      port map(A => \ReadFIFO_Read_Ptr[0]_net_1\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \iRX_FIFO_OVERFLOW[0]\, 
        D => \iRX_FIFO_OVERFLOW[1]\, FCI => VCC_net_1, S => OPEN, 
        Y => RX_FIFO_OVERFLOW_3_0_0_y0, FCO => 
        RX_FIFO_OVERFLOW_3_0_0_co0);
    
    \RX_FIFO_DOUT_3_0_0_wmux[7]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => \ReadFIFO_Read_Ptr[0]_net_1\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \RX_FIFO_DOUT_0[7]\, D
         => \RX_FIFO_DOUT_1[7]\, FCI => VCC_net_1, S => OPEN, Y
         => \RX_FIFO_DOUT_3_0_0_y0[7]\, FCO => 
        \RX_FIFO_DOUT_3_0_0_co0[7]\);
    
    \ReadFIFO_Read_Ptr_RNO[0]\ : CFG3
      generic map(INIT => x"9C")

      port map(A => up_EOP_sync(1), B => 
        \ReadFIFO_Read_Ptr[0]_net_1\, C => up_EOP_sync(2), Y => 
        \ReadFIFO_Read_Ptr_2[0]\);
    
    TRANSMIT_FIFO : FIFO_2Kx8
      port map(TX_FIFO_DOUT(7) => TX_FIFO_DOUT(7), 
        TX_FIFO_DOUT(6) => TX_FIFO_DOUT(6), TX_FIFO_DOUT(5) => 
        TX_FIFO_DOUT(5), TX_FIFO_DOUT(4) => TX_FIFO_DOUT(4), 
        TX_FIFO_DOUT(3) => TX_FIFO_DOUT(3), TX_FIFO_DOUT(2) => 
        TX_FIFO_DOUT(2), TX_FIFO_DOUT(1) => TX_FIFO_DOUT(1), 
        TX_FIFO_DOUT(0) => TX_FIFO_DOUT(0), 
        CoreAPB3_0_APBmslave0_PWDATA(7) => 
        CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), itx_fifo_rst_i => 
        itx_fifo_rst_i, BIT_CLK => BIT_CLK, N_114 => N_114, 
        TX_FIFO_Empty => TX_FIFO_Empty, TX_FIFO_wr_en => 
        TX_FIFO_wr_en, TX_FIFO_Full => TX_FIFO_Full, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz, 
        TX_FIFO_OVERFLOW_i => TX_FIFO_OVERFLOW_i, 
        TX_FIFO_OVERFLOW => TX_FIFO_OVERFLOW, TX_FIFO_UNDERRUN_i
         => TX_FIFO_UNDERRUN_i, TX_FIFO_UNDERRUN => 
        TX_FIFO_UNDERRUN);
    
    \RX_FIFO_DOUT_3_0_0_wmux[0]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => \ReadFIFO_Read_Ptr[0]_net_1\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \RX_FIFO_DOUT_0[0]\, D
         => \RX_FIFO_DOUT_1[0]\, FCI => VCC_net_1, S => OPEN, Y
         => \RX_FIFO_DOUT_3_0_0_y0[0]\, FCO => 
        \RX_FIFO_DOUT_3_0_0_co0[0]\);
    
    RECEIVE_FIFO_1 : FIFO_8Kx9_0
      port map(RX_FIFO_DOUT_1(8) => \RX_FIFO_DOUT_1[8]\, 
        RX_FIFO_DOUT_1(7) => \RX_FIFO_DOUT_1[7]\, 
        RX_FIFO_DOUT_1(6) => \RX_FIFO_DOUT_1[6]\, 
        RX_FIFO_DOUT_1(5) => \RX_FIFO_DOUT_1[5]\, 
        RX_FIFO_DOUT_1(4) => \RX_FIFO_DOUT_1[4]\, 
        RX_FIFO_DOUT_1(3) => \RX_FIFO_DOUT_1[3]\, 
        RX_FIFO_DOUT_1(2) => \RX_FIFO_DOUT_1[2]\, 
        RX_FIFO_DOUT_1(1) => \RX_FIFO_DOUT_1[1]\, 
        RX_FIFO_DOUT_1(0) => \RX_FIFO_DOUT_1[0]\, 
        RX_FIFO_DIN_pipe(8) => RX_FIFO_DIN_pipe(8), 
        RX_FIFO_DIN_pipe(7) => RX_FIFO_DIN_pipe(7), 
        RX_FIFO_DIN_pipe(6) => RX_FIFO_DIN_pipe(6), 
        RX_FIFO_DIN_pipe(5) => RX_FIFO_DIN_pipe(5), 
        RX_FIFO_DIN_pipe(4) => RX_FIFO_DIN_pipe(4), 
        RX_FIFO_DIN_pipe(3) => RX_FIFO_DIN_pipe(3), 
        RX_FIFO_DIN_pipe(2) => RX_FIFO_DIN_pipe(2), 
        RX_FIFO_DIN_pipe(1) => RX_FIFO_DIN_pipe(1), 
        RX_FIFO_DIN_pipe(0) => RX_FIFO_DIN_pipe(0), 
        iRX_FIFO_rd_en_0 => \iRX_FIFO_rd_en[1]\, 
        iRX_FIFO_wr_en_0_0 => \iRX_FIFO_wr_en_0[1]\, 
        iRX_FIFO_Empty_0 => \iRX_FIFO_Empty[1]\, 
        iRX_FIFO_UNDERRUN_0 => \iRX_FIFO_UNDERRUN[1]\, 
        iRX_FIFO_OVERFLOW_0 => \iRX_FIFO_OVERFLOW[1]\, 
        iRX_FIFO_Full_0 => \iRX_FIFO_Full[1]\, irx_fifo_rst_i => 
        irx_fifo_rst_i, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, RX_FIFO_TxColDetDis_wr_en => 
        RX_FIFO_TxColDetDis_wr_en, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0);
    
    \ReadFIFO_Read_Ptr_RNIH36R_0[0]\ : CFG3
      generic map(INIT => x"40")

      port map(A => \ReadFIFO_Read_Ptr[1]_net_1\, B => 
        \ReadFIFO_Read_Ptr[0]_net_1\, C => RX_FIFO_rd_en, Y => 
        \iRX_FIFO_rd_en[1]\);
    
    \RX_FIFO_DOUT_3_0_0_wmux_0[4]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \RX_FIFO_DOUT_3_0_0_y0[4]\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \RX_FIFO_DOUT_2[4]\, D
         => \RX_FIFO_DOUT_3[4]\, FCI => 
        \RX_FIFO_DOUT_3_0_0_co0[4]\, S => OPEN, Y => 
        RX_FIFO_DOUT(4), FCO => OPEN);
    
    \RX_FIFO_DOUT_3_0_0_wmux_0[5]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \RX_FIFO_DOUT_3_0_0_y0[5]\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \RX_FIFO_DOUT_2[5]\, D
         => \RX_FIFO_DOUT_3[5]\, FCI => 
        \RX_FIFO_DOUT_3_0_0_co0[5]\, S => OPEN, Y => 
        RX_FIFO_DOUT(5), FCO => OPEN);
    
    RECEIVE_FIFO_2 : FIFO_8Kx9_1
      port map(RX_FIFO_DOUT_2(8) => \RX_FIFO_DOUT_2[8]\, 
        RX_FIFO_DOUT_2(7) => \RX_FIFO_DOUT_2[7]\, 
        RX_FIFO_DOUT_2(6) => \RX_FIFO_DOUT_2[6]\, 
        RX_FIFO_DOUT_2(5) => \RX_FIFO_DOUT_2[5]\, 
        RX_FIFO_DOUT_2(4) => \RX_FIFO_DOUT_2[4]\, 
        RX_FIFO_DOUT_2(3) => \RX_FIFO_DOUT_2[3]\, 
        RX_FIFO_DOUT_2(2) => \RX_FIFO_DOUT_2[2]\, 
        RX_FIFO_DOUT_2(1) => \RX_FIFO_DOUT_2[1]\, 
        RX_FIFO_DOUT_2(0) => \RX_FIFO_DOUT_2[0]\, 
        RX_FIFO_DIN_pipe(8) => RX_FIFO_DIN_pipe(8), 
        RX_FIFO_DIN_pipe(7) => RX_FIFO_DIN_pipe(7), 
        RX_FIFO_DIN_pipe(6) => RX_FIFO_DIN_pipe(6), 
        RX_FIFO_DIN_pipe(5) => RX_FIFO_DIN_pipe(5), 
        RX_FIFO_DIN_pipe(4) => RX_FIFO_DIN_pipe(4), 
        RX_FIFO_DIN_pipe(3) => RX_FIFO_DIN_pipe(3), 
        RX_FIFO_DIN_pipe(2) => RX_FIFO_DIN_pipe(2), 
        RX_FIFO_DIN_pipe(1) => RX_FIFO_DIN_pipe(1), 
        RX_FIFO_DIN_pipe(0) => RX_FIFO_DIN_pipe(0), 
        iRX_FIFO_rd_en_0 => \iRX_FIFO_rd_en[2]\, 
        iRX_FIFO_wr_en_0_0 => \iRX_FIFO_wr_en_0[2]\, 
        iRX_FIFO_Empty_0 => \iRX_FIFO_Empty[2]\, 
        iRX_FIFO_UNDERRUN_0 => \iRX_FIFO_UNDERRUN[2]\, 
        iRX_FIFO_OVERFLOW_0 => \iRX_FIFO_OVERFLOW[2]\, 
        iRX_FIFO_Full_0 => \iRX_FIFO_Full[2]\, irx_fifo_rst_i => 
        irx_fifo_rst_i, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, RX_FIFO_TxColDetDis_wr_en => 
        RX_FIFO_TxColDetDis_wr_en, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \ReadFIFO_Read_Ptr[0]\ : SLE
      port map(D => \ReadFIFO_Read_Ptr_2[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \ReadFIFO_Read_Ptr[0]_net_1\);
    
    \ReadFIFO_Read_Ptr_RNIH36R_2[0]\ : CFG3
      generic map(INIT => x"10")

      port map(A => \ReadFIFO_Read_Ptr[1]_net_1\, B => 
        \ReadFIFO_Read_Ptr[0]_net_1\, C => RX_FIFO_rd_en, Y => 
        \iRX_FIFO_rd_en[0]\);
    
    itx_fifo_rst_RNIUMSA : CLKINT
      port map(A => \itx_fifo_rst\, Y => itx_fifo_rst_i);
    
    RX_FIFO_UNDERRUN_3_0_0_wmux_0_RNIS837 : CFG1
      generic map(INIT => "01")

      port map(A => \RX_FIFO_UNDERRUN\, Y => RX_FIFO_UNDERRUN_i);
    
    irx_fifo_rst : CFG2
      generic map(INIT => x"1")

      port map(A => RX_FIFO_RST, B => RESET, Y => \irx_fifo_rst\);
    
    \packet_available_clear_reg[0]\ : SLE
      port map(D => rx_packet_avail_int, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \packet_available_clear_reg[0]_net_1\);
    
    \ReadFIFO_Write_Ptr_RNIBKOU[1]\ : CFG2
      generic map(INIT => x"8")

      port map(A => \ReadFIFO_Write_Ptr[0]_net_1\, B => 
        \ReadFIFO_Write_Ptr[1]_net_1\, Y => \iRX_FIFO_wr_en_0[3]\);
    
    \RX_FIFO_DOUT_3_0_0_wmux_0[7]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \RX_FIFO_DOUT_3_0_0_y0[7]\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \RX_FIFO_DOUT_2[7]\, D
         => \RX_FIFO_DOUT_3[7]\, FCI => 
        \RX_FIFO_DOUT_3_0_0_co0[7]\, S => OPEN, Y => 
        RX_FIFO_DOUT(7), FCO => OPEN);
    
    \RX_FIFO_DOUT_3_0_0_wmux_0[2]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \RX_FIFO_DOUT_3_0_0_y0[2]\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \RX_FIFO_DOUT_2[2]\, D
         => \RX_FIFO_DOUT_3[2]\, FCI => 
        \RX_FIFO_DOUT_3_0_0_co0[2]\, S => OPEN, Y => 
        RX_FIFO_DOUT(2), FCO => OPEN);
    
    \ReadFIFO_Write_Ptr_RNIBKOU_0[1]\ : CFG2
      generic map(INIT => x"4")

      port map(A => \ReadFIFO_Write_Ptr[0]_net_1\, B => 
        \ReadFIFO_Write_Ptr[1]_net_1\, Y => \iRX_FIFO_wr_en_0[2]\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \ReadFIFO_Write_Ptr_RNO[1]\ : CFG3
      generic map(INIT => x"78")

      port map(A => \ReadFIFO_Write_Ptr[0]_net_1\, B => 
        rx_packet_complt, C => \ReadFIFO_Write_Ptr[1]_net_1\, Y
         => \ReadFIFO_Write_Ptr_3[1]\);
    
    \RX_FIFO_DOUT_3_0_0_wmux[3]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => \ReadFIFO_Read_Ptr[0]_net_1\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \RX_FIFO_DOUT_0[3]\, D
         => \RX_FIFO_DOUT_1[3]\, FCI => VCC_net_1, S => OPEN, Y
         => \RX_FIFO_DOUT_3_0_0_y0[3]\, FCO => 
        \RX_FIFO_DOUT_3_0_0_co0[3]\);
    
    RX_FIFO_UNDERRUN_3_0_0_wmux_0 : ARI1
      generic map(INIT => x"0F588")

      port map(A => RX_FIFO_UNDERRUN_3_0_0_y0, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \iRX_FIFO_UNDERRUN[2]\, 
        D => \iRX_FIFO_UNDERRUN[3]\, FCI => 
        RX_FIFO_UNDERRUN_3_0_0_co0, S => OPEN, Y => 
        \RX_FIFO_UNDERRUN\, FCO => OPEN);
    
    RX_FIFO_Empty_3_0_0_wmux_0 : ARI1
      generic map(INIT => x"0F588")

      port map(A => RX_FIFO_Empty_3_0_0_y0, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \iRX_FIFO_Empty[2]\, D
         => \iRX_FIFO_Empty[3]\, FCI => RX_FIFO_Empty_3_0_0_co0, 
        S => OPEN, Y => RX_FIFO_Empty, FCO => OPEN);
    
    \ReadFIFO_Write_Ptr[0]\ : SLE
      port map(D => \ReadFIFO_Write_Ptr_3[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \ReadFIFO_Write_Ptr[0]_net_1\);
    
    \RX_FIFO_DOUT_3_0_0_wmux_0[0]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \RX_FIFO_DOUT_3_0_0_y0[0]\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \RX_FIFO_DOUT_2[0]\, D
         => \RX_FIFO_DOUT_3[0]\, FCI => 
        \RX_FIFO_DOUT_3_0_0_co0[0]\, S => OPEN, Y => 
        RX_FIFO_DOUT(0), FCO => OPEN);
    
    RECEIVE_FIFO_3 : FIFO_8Kx9_2
      port map(RX_FIFO_DOUT_3(8) => \RX_FIFO_DOUT_3[8]\, 
        RX_FIFO_DOUT_3(7) => \RX_FIFO_DOUT_3[7]\, 
        RX_FIFO_DOUT_3(6) => \RX_FIFO_DOUT_3[6]\, 
        RX_FIFO_DOUT_3(5) => \RX_FIFO_DOUT_3[5]\, 
        RX_FIFO_DOUT_3(4) => \RX_FIFO_DOUT_3[4]\, 
        RX_FIFO_DOUT_3(3) => \RX_FIFO_DOUT_3[3]\, 
        RX_FIFO_DOUT_3(2) => \RX_FIFO_DOUT_3[2]\, 
        RX_FIFO_DOUT_3(1) => \RX_FIFO_DOUT_3[1]\, 
        RX_FIFO_DOUT_3(0) => \RX_FIFO_DOUT_3[0]\, 
        RX_FIFO_DIN_pipe(8) => RX_FIFO_DIN_pipe(8), 
        RX_FIFO_DIN_pipe(7) => RX_FIFO_DIN_pipe(7), 
        RX_FIFO_DIN_pipe(6) => RX_FIFO_DIN_pipe(6), 
        RX_FIFO_DIN_pipe(5) => RX_FIFO_DIN_pipe(5), 
        RX_FIFO_DIN_pipe(4) => RX_FIFO_DIN_pipe(4), 
        RX_FIFO_DIN_pipe(3) => RX_FIFO_DIN_pipe(3), 
        RX_FIFO_DIN_pipe(2) => RX_FIFO_DIN_pipe(2), 
        RX_FIFO_DIN_pipe(1) => RX_FIFO_DIN_pipe(1), 
        RX_FIFO_DIN_pipe(0) => RX_FIFO_DIN_pipe(0), 
        iRX_FIFO_rd_en_0 => \iRX_FIFO_rd_en[3]\, 
        iRX_FIFO_wr_en_0_0 => \iRX_FIFO_wr_en_0[3]\, 
        iRX_FIFO_Empty_0 => \iRX_FIFO_Empty[3]\, 
        iRX_FIFO_UNDERRUN_0 => \iRX_FIFO_UNDERRUN[3]\, 
        iRX_FIFO_OVERFLOW_0 => \iRX_FIFO_OVERFLOW[3]\, 
        iRX_FIFO_Full_0 => \iRX_FIFO_Full[3]\, irx_fifo_rst_i => 
        irx_fifo_rst_i, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, RX_FIFO_TxColDetDis_wr_en => 
        RX_FIFO_TxColDetDis_wr_en, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0);
    
    \RX_FIFO_DOUT_3_0_0_wmux_0[8]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \RX_FIFO_DOUT_3_0_0_y0[8]\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \RX_FIFO_DOUT_2[8]\, D
         => \RX_FIFO_DOUT_3[8]\, FCI => 
        \RX_FIFO_DOUT_3_0_0_co0[8]\, S => OPEN, Y => 
        RX_FIFO_DOUT(8), FCO => OPEN);
    
    \ReadFIFO_Read_Ptr_RNIH36R[0]\ : CFG3
      generic map(INIT => x"80")

      port map(A => \ReadFIFO_Read_Ptr[1]_net_1\, B => 
        \ReadFIFO_Read_Ptr[0]_net_1\, C => RX_FIFO_rd_en, Y => 
        \iRX_FIFO_rd_en[3]\);
    
    \ReadFIFO_Write_Ptr_RNIBKOU_1[1]\ : CFG2
      generic map(INIT => x"2")

      port map(A => \ReadFIFO_Write_Ptr[0]_net_1\, B => 
        \ReadFIFO_Write_Ptr[1]_net_1\, Y => \iRX_FIFO_wr_en_0[1]\);
    
    \ReadFIFO_Write_Ptr_RNO[0]\ : CFG2
      generic map(INIT => x"6")

      port map(A => rx_packet_complt, B => 
        \ReadFIFO_Write_Ptr[0]_net_1\, Y => 
        \ReadFIFO_Write_Ptr_3[0]\);
    
    itx_fifo_rst : CFG2
      generic map(INIT => x"1")

      port map(A => RESET, B => TX_FIFO_RST, Y => \itx_fifo_rst\);
    
    \RX_FIFO_DOUT_3_0_0_wmux[8]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => \ReadFIFO_Read_Ptr[0]_net_1\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \RX_FIFO_DOUT_0[8]\, D
         => \RX_FIFO_DOUT_1[8]\, FCI => VCC_net_1, S => OPEN, Y
         => \RX_FIFO_DOUT_3_0_0_y0[8]\, FCO => 
        \RX_FIFO_DOUT_3_0_0_co0[8]\);
    
    RECEIVE_FIFO_0 : FIFO_8Kx9
      port map(RX_FIFO_DOUT_0(8) => \RX_FIFO_DOUT_0[8]\, 
        RX_FIFO_DOUT_0(7) => \RX_FIFO_DOUT_0[7]\, 
        RX_FIFO_DOUT_0(6) => \RX_FIFO_DOUT_0[6]\, 
        RX_FIFO_DOUT_0(5) => \RX_FIFO_DOUT_0[5]\, 
        RX_FIFO_DOUT_0(4) => \RX_FIFO_DOUT_0[4]\, 
        RX_FIFO_DOUT_0(3) => \RX_FIFO_DOUT_0[3]\, 
        RX_FIFO_DOUT_0(2) => \RX_FIFO_DOUT_0[2]\, 
        RX_FIFO_DOUT_0(1) => \RX_FIFO_DOUT_0[1]\, 
        RX_FIFO_DOUT_0(0) => \RX_FIFO_DOUT_0[0]\, 
        RX_FIFO_DIN_pipe(8) => RX_FIFO_DIN_pipe(8), 
        RX_FIFO_DIN_pipe(7) => RX_FIFO_DIN_pipe(7), 
        RX_FIFO_DIN_pipe(6) => RX_FIFO_DIN_pipe(6), 
        RX_FIFO_DIN_pipe(5) => RX_FIFO_DIN_pipe(5), 
        RX_FIFO_DIN_pipe(4) => RX_FIFO_DIN_pipe(4), 
        RX_FIFO_DIN_pipe(3) => RX_FIFO_DIN_pipe(3), 
        RX_FIFO_DIN_pipe(2) => RX_FIFO_DIN_pipe(2), 
        RX_FIFO_DIN_pipe(1) => RX_FIFO_DIN_pipe(1), 
        RX_FIFO_DIN_pipe(0) => RX_FIFO_DIN_pipe(0), 
        iRX_FIFO_rd_en_0 => \iRX_FIFO_rd_en[0]\, 
        iRX_FIFO_wr_en_0_0 => \iRX_FIFO_wr_en_0[0]\, 
        iRX_FIFO_Empty_0 => \iRX_FIFO_Empty[0]\, 
        iRX_FIFO_UNDERRUN_0 => \iRX_FIFO_UNDERRUN[0]\, 
        iRX_FIFO_OVERFLOW_0 => \iRX_FIFO_OVERFLOW[0]\, 
        iRX_FIFO_Full_0 => \iRX_FIFO_Full[0]\, irx_fifo_rst_i => 
        irx_fifo_rst_i, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, RX_FIFO_TxColDetDis_wr_en => 
        RX_FIFO_TxColDetDis_wr_en, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0);
    
    \ReadFIFO_Read_Ptr[1]\ : SLE
      port map(D => \ReadFIFO_Read_Ptr_2[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \ReadFIFO_Read_Ptr[1]_net_1\);
    
    \RX_FIFO_DOUT_3_0_0_wmux_0[3]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \RX_FIFO_DOUT_3_0_0_y0[3]\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \RX_FIFO_DOUT_2[3]\, D
         => \RX_FIFO_DOUT_3[3]\, FCI => 
        \RX_FIFO_DOUT_3_0_0_co0[3]\, S => OPEN, Y => 
        RX_FIFO_DOUT(3), FCO => OPEN);
    
    \RX_FIFO_DOUT_3_0_0_wmux[1]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => \ReadFIFO_Read_Ptr[0]_net_1\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \RX_FIFO_DOUT_0[1]\, D
         => \RX_FIFO_DOUT_1[1]\, FCI => VCC_net_1, S => OPEN, Y
         => \RX_FIFO_DOUT_3_0_0_y0[1]\, FCO => 
        \RX_FIFO_DOUT_3_0_0_co0[1]\);
    
    \packet_available_clear_reg[1]\ : SLE
      port map(D => \packet_available_clear_reg[0]_net_1\, CLK
         => CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \packet_available_clear_reg[1]_net_1\);
    
    RX_FIFO_Full_3_0_0_wmux_0 : ARI1
      generic map(INIT => x"0F588")

      port map(A => RX_FIFO_Full_3_0_0_y0, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \iRX_FIFO_Full[2]\, D
         => \iRX_FIFO_Full[3]\, FCI => RX_FIFO_Full_3_0_0_co0, S
         => OPEN, Y => RX_FIFO_Full, FCO => OPEN);
    
    \ReadFIFO_Read_Ptr_RNIH36R_1[0]\ : CFG3
      generic map(INIT => x"20")

      port map(A => \ReadFIFO_Read_Ptr[1]_net_1\, B => 
        \ReadFIFO_Read_Ptr[0]_net_1\, C => RX_FIFO_rd_en, Y => 
        \iRX_FIFO_rd_en[2]\);
    
    \RX_FIFO_DOUT_3_0_0_wmux[2]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => \ReadFIFO_Read_Ptr[0]_net_1\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \RX_FIFO_DOUT_0[2]\, D
         => \RX_FIFO_DOUT_1[2]\, FCI => VCC_net_1, S => OPEN, Y
         => \RX_FIFO_DOUT_3_0_0_y0[2]\, FCO => 
        \RX_FIFO_DOUT_3_0_0_co0[2]\);
    
    RX_FIFO_OVERFLOW_3_0_0_wmux_0 : ARI1
      generic map(INIT => x"0F588")

      port map(A => RX_FIFO_OVERFLOW_3_0_0_y0, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \iRX_FIFO_OVERFLOW[2]\, 
        D => \iRX_FIFO_OVERFLOW[3]\, FCI => 
        RX_FIFO_OVERFLOW_3_0_0_co0, S => OPEN, Y => 
        \RX_FIFO_OVERFLOW\, FCO => OPEN);
    
    RX_FIFO_OVERFLOW_3_0_0_wmux_0_RNITUE2 : CFG1
      generic map(INIT => "01")

      port map(A => \RX_FIFO_OVERFLOW\, Y => RX_FIFO_OVERFLOW_i);
    
    \RX_FIFO_DOUT_3_0_0_wmux[5]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => \ReadFIFO_Read_Ptr[0]_net_1\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \RX_FIFO_DOUT_0[5]\, D
         => \RX_FIFO_DOUT_1[5]\, FCI => VCC_net_1, S => OPEN, Y
         => \RX_FIFO_DOUT_3_0_0_y0[5]\, FCO => 
        \RX_FIFO_DOUT_3_0_0_co0[5]\);
    
    \ReadFIFO_Write_Ptr[1]\ : SLE
      port map(D => \ReadFIFO_Write_Ptr_3[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \ReadFIFO_Write_Ptr[1]_net_1\);
    
    \ReadFIFO_Write_Ptr_RNIBKOU_2[1]\ : CFG2
      generic map(INIT => x"1")

      port map(A => \ReadFIFO_Write_Ptr[0]_net_1\, B => 
        \ReadFIFO_Write_Ptr[1]_net_1\, Y => \iRX_FIFO_wr_en_0[0]\);
    
    \packet_available_clear_reg[2]\ : SLE
      port map(D => \packet_available_clear_reg[1]_net_1\, CLK
         => CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => 
        irx_fifo_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        packet_available_clear_reg(2));
    
    \RX_FIFO_DOUT_3_0_0_wmux_0[1]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \RX_FIFO_DOUT_3_0_0_y0[1]\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \RX_FIFO_DOUT_2[1]\, D
         => \RX_FIFO_DOUT_3[1]\, FCI => 
        \RX_FIFO_DOUT_3_0_0_co0[1]\, S => OPEN, Y => 
        RX_FIFO_DOUT(1), FCO => OPEN);
    
    \RX_FIFO_DOUT_3_0_0_wmux[4]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => \ReadFIFO_Read_Ptr[0]_net_1\, B => 
        \ReadFIFO_Read_Ptr[1]_net_1\, C => \RX_FIFO_DOUT_0[4]\, D
         => \RX_FIFO_DOUT_1[4]\, FCI => VCC_net_1, S => OPEN, Y
         => \RX_FIFO_DOUT_3_0_0_y0[4]\, FCO => 
        \RX_FIFO_DOUT_3_0_0_co0[4]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity Interrupts is

    port( CoreAPB3_0_APBmslave0_PADDR  : in    std_logic_vector(3 downto 2);
          CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 1);
          int_reg                      : out   std_logic_vector(7 downto 1);
          i_int_mask_reg               : in    std_logic_vector(7 downto 1);
          up_EOP_del                   : out   std_logic_vector(5 downto 0);
          N_218                        : in    std_logic;
          write_reg_en                 : in    std_logic;
          CommsFPGA_top_0_INT          : out   std_logic;
          RESET                        : in    std_logic;
          int_reg_clr                  : out   std_logic;
          long_reset                   : in    std_logic;
          RX_packet_depth_status       : in    std_logic;
          tx_packet_complt_int         : out   std_logic;
          TX_FIFO_UNDERRUN             : in    std_logic;
          un15_int_reg_clr             : out   std_logic;
          TX_FIFO_UNDERRUN_set         : in    std_logic;
          TX_FIFO_OVERFLOW             : in    std_logic;
          un19_int_reg_clr             : out   std_logic;
          TX_FIFO_OVERFLOW_set         : in    std_logic;
          RX_FIFO_UNDERRUN             : in    std_logic;
          un23_int_reg_clr             : out   std_logic;
          rx_FIFO_UNDERRUN_int         : out   std_logic;
          RX_FIFO_UNDERRUN_set         : in    std_logic;
          RX_FIFO_OVERFLOW             : in    std_logic;
          un27_int_reg_clr             : out   std_logic;
          rx_FIFO_OVERFLOW_int         : out   std_logic;
          RX_FIFO_OVERFLOW_set         : in    std_logic;
          rx_CRC_error                 : in    std_logic;
          un31_int_reg_clr             : out   std_logic;
          rx_CRC_error_int             : out   std_logic;
          rx_CRC_error_set             : in    std_logic;
          rx_packet_avail_int          : out   std_logic;
          tx_packet_complt             : in    std_logic;
          iup_EOP                      : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic;
          CommsFPGA_CCC_0_GL0          : in    std_logic;
          RESET_i                      : in    std_logic;
          block_int_until_rd           : out   std_logic
        );

end Interrupts;

architecture DEF_ARCH of Interrupts is 

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal un2_apb3_reset, un2_apb3_reset_0, 
        block_int_until_rd_net_1, block_int_until_rd_i, 
        \tx_packet_complt_toClk16x\, tx_packet_complt_toClk16x_i, 
        un2_apb3_reset_i, \tx_packet_complt_d[6]_net_1\, 
        VCC_net_1, \tx_packet_complt_d[5]_net_1\, GND_net_1, 
        \tx_packet_complt_d[7]_net_1\, \up_EOP_del[0]_net_1\, 
        \up_EOP_del[1]_net_1\, \up_EOP_del[2]_net_1\, 
        \up_EOP_del[3]_net_1\, \up_EOP_del[4]_net_1\, 
        \up_EOP_del[5]_net_1\, \tx_packet_complt_d[0]_net_1\, 
        \tx_packet_complt_d[1]_net_1\, 
        \tx_packet_complt_d[2]_net_1\, 
        \tx_packet_complt_d[3]_net_1\, 
        \tx_packet_complt_d[4]_net_1\, \rx_packet_avail_int\, 
        un15_apb3_reset_i, un1_N_5_mux_0_i, 
        \block_int_until_rd_RNO\, un2_apb3_reset_rs_3, 
        rx_CRC_error_intrs, rx_CRC_error_int_net_1, 
        \un31_int_reg_clr\, un2_apb3_reset_rs_2, 
        rx_FIFO_OVERFLOW_intrs, rx_FIFO_OVERFLOW_int_net_1, 
        \un27_int_reg_clr\, un2_apb3_reset_rs_1, 
        rx_FIFO_UNDERRUN_intrs, rx_FIFO_UNDERRUN_int_net_1, 
        \un23_int_reg_clr\, tx_FIFO_OVERFLOW_intrs, 
        un2_apb3_reset_rs_0, \tx_FIFO_OVERFLOW_int\, 
        \un19_int_reg_clr\, tx_FIFO_UNDERRUN_intrs, 
        un2_apb3_reset_rs, \tx_FIFO_UNDERRUN_int\, 
        \un15_int_reg_clr\, \tx_packet_complt_toClk16x_set\, 
        tx_packet_complt_intrs, un6_apb3_reset_rs, 
        tx_packet_complt_int_net_1, un6_apb3_reset_i, 
        un5_int_reg_clr, un1_N_5_mux_0_i_1, N_385, \int_reg[1]\, 
        \int_reg[2]\, \int_reg[3]\, \int_reg[4]\, \int_reg[5]\, 
        \int_reg[6]\, \int_reg[7]\, \INT_4\ : std_logic;

begin 

    int_reg(7) <= \int_reg[7]\;
    int_reg(6) <= \int_reg[6]\;
    int_reg(5) <= \int_reg[5]\;
    int_reg(4) <= \int_reg[4]\;
    int_reg(3) <= \int_reg[3]\;
    int_reg(2) <= \int_reg[2]\;
    int_reg(1) <= \int_reg[1]\;
    up_EOP_del(5) <= \up_EOP_del[5]_net_1\;
    up_EOP_del(4) <= \up_EOP_del[4]_net_1\;
    up_EOP_del(3) <= \up_EOP_del[3]_net_1\;
    up_EOP_del(2) <= \up_EOP_del[2]_net_1\;
    up_EOP_del(1) <= \up_EOP_del[1]_net_1\;
    up_EOP_del(0) <= \up_EOP_del[0]_net_1\;
    tx_packet_complt_int <= tx_packet_complt_int_net_1;
    un15_int_reg_clr <= \un15_int_reg_clr\;
    un19_int_reg_clr <= \un19_int_reg_clr\;
    un23_int_reg_clr <= \un23_int_reg_clr\;
    rx_FIFO_UNDERRUN_int <= rx_FIFO_UNDERRUN_int_net_1;
    un27_int_reg_clr <= \un27_int_reg_clr\;
    rx_FIFO_OVERFLOW_int <= rx_FIFO_OVERFLOW_int_net_1;
    un31_int_reg_clr <= \un31_int_reg_clr\;
    rx_CRC_error_int <= rx_CRC_error_int_net_1;
    rx_packet_avail_int <= \rx_packet_avail_int\;
    block_int_until_rd <= block_int_until_rd_net_1;

    irx_packet_avail_int_RNIF9DL : CFG2
      generic map(INIT => x"2")

      port map(A => \rx_packet_avail_int\, B => i_int_mask_reg(6), 
        Y => \int_reg[6]\);
    
    \TX_PACKET_COMPLETE_INTR.un2_apb3_reset_rs_3\ : SLE
      port map(D => VCC_net_1, CLK => rx_CRC_error, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        un2_apb3_reset_rs_3);
    
    \up_EOP_del[1]\ : SLE
      port map(D => \up_EOP_del[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \up_EOP_del[1]_net_1\);
    
    \TX_PACKET_COMPLETE_INTR.un2_apb3_reset_rs_1_RNIVKP21\ : CFG2
      generic map(INIT => x"2")

      port map(A => rx_FIFO_UNDERRUN_int_net_1, B => 
        i_int_mask_reg(3), Y => \int_reg[3]\);
    
    tx_packet_complt_toClk16x_set_RNO : CFG1
      generic map(INIT => "01")

      port map(A => \tx_packet_complt_toClk16x\, Y => 
        tx_packet_complt_toClk16x_i);
    
    \REGISTER_CLEAR_INST.un1_write_reg_en\ : CFG4
      generic map(INIT => x"0800")

      port map(A => write_reg_en, B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => N_218, Y => N_385);
    
    \RX_PACKET_AVAILABLE_INTR.un15_apb3_reset\ : CFG4
      generic map(INIT => x"0001")

      port map(A => rx_FIFO_UNDERRUN_int_net_1, B => 
        rx_FIFO_OVERFLOW_int_net_1, C => rx_CRC_error_int_net_1, 
        D => un2_apb3_reset, Y => un15_apb3_reset_i);
    
    tx_FIFO_UNDERRUN_int_RNI6GG01 : CFG3
      generic map(INIT => x"EC")

      port map(A => TX_FIFO_UNDERRUN_set, B => 
        tx_FIFO_UNDERRUN_intrs, C => un2_apb3_reset_rs, Y => 
        \tx_FIFO_UNDERRUN_int\);
    
    \TX_FIFO_UNDERRUN_INTR.un15_int_reg_clr_0_a2\ : CFG3
      generic map(INIT => x"20")

      port map(A => N_385, B => long_reset, C => 
        CoreAPB3_0_APBmslave0_PWDATA(5), Y => \un15_int_reg_clr\);
    
    \RX_FIFO_OVERFLOW_INTR.un27_int_reg_clr\ : CFG3
      generic map(INIT => x"20")

      port map(A => N_385, B => long_reset, C => 
        CoreAPB3_0_APBmslave0_PWDATA(2), Y => \un27_int_reg_clr\);
    
    \up_EOP_del[0]\ : SLE
      port map(D => iup_EOP, CLK => m2s010_som_sb_0_CCC_71MHz, EN
         => VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \up_EOP_del[0]_net_1\);
    
    \TX_PACKET_COMPLETE_INTR.un2_apb3_reset_rs_3_RNIL7BV\ : CFG2
      generic map(INIT => x"2")

      port map(A => rx_CRC_error_int_net_1, B => 
        i_int_mask_reg(1), Y => \int_reg[1]\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \up_EOP_del[5]\ : SLE
      port map(D => \up_EOP_del[4]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \up_EOP_del[5]_net_1\);
    
    irx_packet_avail_int : SLE
      port map(D => block_int_until_rd_i, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un1_N_5_mux_0_i, ALn => 
        un15_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \rx_packet_avail_int\);
    
    \TX_FIFO_OVERFLOW_INTR.un19_int_reg_clr\ : CFG3
      generic map(INIT => x"20")

      port map(A => N_385, B => long_reset, C => 
        CoreAPB3_0_APBmslave0_PWDATA(4), Y => \un19_int_reg_clr\);
    
    \tx_packet_complt_d[0]\ : SLE
      port map(D => tx_packet_complt, CLK => CommsFPGA_CCC_0_GL0, 
        EN => VCC_net_1, ALn => RESET_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \tx_packet_complt_d[0]_net_1\);
    
    \RX_CRC_ERROR_INTR.un31_int_reg_clr\ : CFG3
      generic map(INIT => x"20")

      port map(A => N_385, B => long_reset, C => 
        CoreAPB3_0_APBmslave0_PWDATA(1), Y => \un31_int_reg_clr\);
    
    int_reg_clr_0_a2_0_a2 : CFG2
      generic map(INIT => x"4")

      port map(A => long_reset, B => N_385, Y => int_reg_clr);
    
    \TX_PACKET_COMPLETE_INTR.un5_int_reg_clr\ : CFG3
      generic map(INIT => x"20")

      port map(A => N_385, B => long_reset, C => 
        CoreAPB3_0_APBmslave0_PWDATA(7), Y => un5_int_reg_clr);
    
    \TX_PACKET_COMPLETE_INTR.un2_apb3_reset_rs_2_RNIL9OK\ : CFG3
      generic map(INIT => x"F8")

      port map(A => RX_FIFO_OVERFLOW_set, B => 
        un2_apb3_reset_rs_2, C => rx_FIFO_OVERFLOW_intrs, Y => 
        rx_FIFO_OVERFLOW_int_net_1);
    
    \TX_PACKET_COMPLETE_INTR.un2_apb3_reset_rs_0_RNI5SCL\ : CFG2
      generic map(INIT => x"2")

      port map(A => \tx_FIFO_OVERFLOW_int\, B => 
        i_int_mask_reg(4), Y => \int_reg[4]\);
    
    \tx_packet_complt_d[7]\ : SLE
      port map(D => \tx_packet_complt_d[6]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_packet_complt_d[7]_net_1\);
    
    \TX_PACKET_COMPLETE_INTR.un2_apb3_reset_rs_2\ : SLE
      port map(D => VCC_net_1, CLK => RX_FIFO_OVERFLOW, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        un2_apb3_reset_rs_2);
    
    tx_FIFO_OVERFLOW_int : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \un19_int_reg_clr\, ALn => un2_apb3_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => tx_FIFO_OVERFLOW_intrs);
    
    \rx_CRC_error_int\ : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \un31_int_reg_clr\, ALn => un2_apb3_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => rx_CRC_error_intrs);
    
    \TX_PACKET_COMPLETE_INTR.un2_apb3_reset_rs\ : SLE
      port map(D => VCC_net_1, CLK => TX_FIFO_UNDERRUN, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        un2_apb3_reset_rs);
    
    tx_FIFO_UNDERRUN_int : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \un15_int_reg_clr\, ALn => un2_apb3_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => tx_FIFO_UNDERRUN_intrs);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    tx_FIFO_UNDERRUN_int_RNILNM71 : CFG2
      generic map(INIT => x"2")

      port map(A => \tx_FIFO_UNDERRUN_int\, B => 
        i_int_mask_reg(5), Y => \int_reg[5]\);
    
    \tx_packet_complt_d[5]\ : SLE
      port map(D => \tx_packet_complt_d[4]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_packet_complt_d[5]_net_1\);
    
    \tx_packet_complt_d[4]\ : SLE
      port map(D => \tx_packet_complt_d[3]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_packet_complt_d[4]_net_1\);
    
    \TX_PACKET_COMPLETE_INTR.un2_apb3_reset_rs_1_RNIIFJR\ : CFG3
      generic map(INIT => x"F8")

      port map(A => RX_FIFO_UNDERRUN_set, B => 
        un2_apb3_reset_rs_1, C => rx_FIFO_UNDERRUN_intrs, Y => 
        rx_FIFO_UNDERRUN_int_net_1);
    
    \tx_packet_complt_d[3]\ : SLE
      port map(D => \tx_packet_complt_d[2]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_packet_complt_d[3]_net_1\);
    
    \TX_PACKET_COMPLETE_INTR.un2_apb3_reset_rs_3_RNIA45O\ : CFG3
      generic map(INIT => x"F8")

      port map(A => rx_CRC_error_set, B => un2_apb3_reset_rs_3, C
         => rx_CRC_error_intrs, Y => rx_CRC_error_int_net_1);
    
    \tx_packet_complt_int\ : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => un5_int_reg_clr, ALn => un6_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => tx_packet_complt_intrs);
    
    irx_packet_avail_int_RNO : CFG1
      generic map(INIT => "01")

      port map(A => block_int_until_rd_net_1, Y => 
        block_int_until_rd_i);
    
    \tx_packet_complt_d[6]\ : SLE
      port map(D => \tx_packet_complt_d[5]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_packet_complt_d[6]_net_1\);
    
    \TX_PACKET_COMPLETE_INTR.un2_apb3_reset\ : CFG2
      generic map(INIT => x"E")

      port map(A => long_reset, B => RESET, Y => un2_apb3_reset_0);
    
    INT_4 : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \int_reg[5]\, B => \int_reg[3]\, C => 
        \int_reg[2]\, D => \int_reg[1]\, Y => \INT_4\);
    
    \block_int_until_rd\ : SLE
      port map(D => \block_int_until_rd_RNO\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un1_N_5_mux_0_i, ALn => 
        un15_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        block_int_until_rd_net_1);
    
    \TX_PACKET_COMPLETE_INTR.un2_apb3_reset_rs_0\ : SLE
      port map(D => VCC_net_1, CLK => TX_FIFO_OVERFLOW, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        un2_apb3_reset_rs_0);
    
    block_int_until_rd_RNIRNGP1 : CFG4
      generic map(INIT => x"1D0C")

      port map(A => \rx_packet_avail_int\, B => 
        block_int_until_rd_net_1, C => un1_N_5_mux_0_i_1, D => 
        RX_packet_depth_status, Y => un1_N_5_mux_0_i);
    
    tx_packet_complt_toClk16x : CFG2
      generic map(INIT => x"2")

      port map(A => \tx_packet_complt_d[6]_net_1\, B => 
        \tx_packet_complt_d[7]_net_1\, Y => 
        \tx_packet_complt_toClk16x\);
    
    \TX_PACKET_COMPLETE_INTR.un2_apb3_reset_RNI0RDF_0\ : CFG1
      generic map(INIT => "01")

      port map(A => un2_apb3_reset, Y => un2_apb3_reset_i);
    
    \RX_FIFO_UNDERRUN_INTR.un23_int_reg_clr\ : CFG3
      generic map(INIT => x"20")

      port map(A => N_385, B => long_reset, C => 
        CoreAPB3_0_APBmslave0_PWDATA(3), Y => \un23_int_reg_clr\);
    
    \rx_FIFO_OVERFLOW_int\ : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \un27_int_reg_clr\, ALn => un2_apb3_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => rx_FIFO_OVERFLOW_intrs);
    
    \up_EOP_del_RNI9V2U[5]\ : CFG4
      generic map(INIT => x"00F7")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(6), B => N_385, 
        C => long_reset, D => \up_EOP_del[5]_net_1\, Y => 
        un1_N_5_mux_0_i_1);
    
    \TX_PACKET_COMPLETE_INTR.un2_apb3_reset_rs_2_RNI1EUR\ : CFG2
      generic map(INIT => x"2")

      port map(A => rx_FIFO_OVERFLOW_int_net_1, B => 
        i_int_mask_reg(2), Y => \int_reg[2]\);
    
    \up_EOP_del[4]\ : SLE
      port map(D => \up_EOP_del[3]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \up_EOP_del[4]_net_1\);
    
    \tx_packet_complt_d[1]\ : SLE
      port map(D => \tx_packet_complt_d[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_packet_complt_d[1]_net_1\);
    
    \tx_packet_complt_d[2]\ : SLE
      port map(D => \tx_packet_complt_d[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => RESET_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \tx_packet_complt_d[2]_net_1\);
    
    block_int_until_rd_RNO : CFG4
      generic map(INIT => x"08FF")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(6), B => N_385, 
        C => long_reset, D => block_int_until_rd_net_1, Y => 
        \block_int_until_rd_RNO\);
    
    tx_packet_complt_toClk16x_set_RNI9HQV : CFG2
      generic map(INIT => x"2")

      port map(A => tx_packet_complt_int_net_1, B => 
        i_int_mask_reg(7), Y => \int_reg[7]\);
    
    \TX_PACKET_COMPLETE_INTR.un6_apb3_reset\ : CFG2
      generic map(INIT => x"1")

      port map(A => un2_apb3_reset, B => \tx_FIFO_UNDERRUN_int\, 
        Y => un6_apb3_reset_i);
    
    \TX_PACKET_COMPLETE_INTR.un6_apb3_reset_rs\ : SLE
      port map(D => VCC_net_1, CLK => \tx_packet_complt_toClk16x\, 
        EN => VCC_net_1, ALn => un6_apb3_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        VCC_net_1, Q => un6_apb3_reset_rs);
    
    \TX_PACKET_COMPLETE_INTR.un2_apb3_reset_rs_1\ : SLE
      port map(D => VCC_net_1, CLK => RX_FIFO_UNDERRUN, EN => 
        VCC_net_1, ALn => un2_apb3_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => VCC_net_1, Q => 
        un2_apb3_reset_rs_1);
    
    \TX_PACKET_COMPLETE_INTR.un2_apb3_reset_rs_0_RNINL6E\ : CFG3
      generic map(INIT => x"EC")

      port map(A => TX_FIFO_OVERFLOW_set, B => 
        tx_FIFO_OVERFLOW_intrs, C => un2_apb3_reset_rs_0, Y => 
        \tx_FIFO_OVERFLOW_int\);
    
    INT : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \int_reg[7]\, B => \INT_4\, C => \int_reg[6]\, 
        D => \int_reg[4]\, Y => CommsFPGA_top_0_INT);
    
    \TX_PACKET_COMPLETE_INTR.un2_apb3_reset_RNI0RDF\ : CLKINT
      port map(A => un2_apb3_reset_0, Y => un2_apb3_reset);
    
    \up_EOP_del[3]\ : SLE
      port map(D => \up_EOP_del[2]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \up_EOP_del[3]_net_1\);
    
    \up_EOP_del[2]\ : SLE
      port map(D => \up_EOP_del[1]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        un2_apb3_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        \up_EOP_del[2]_net_1\);
    
    tx_packet_complt_toClk16x_set : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => un5_int_reg_clr, ALn => tx_packet_complt_toClk16x_i, 
        ADn => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \tx_packet_complt_toClk16x_set\);
    
    tx_packet_complt_toClk16x_set_RNIO7KO : CFG3
      generic map(INIT => x"EC")

      port map(A => \tx_packet_complt_toClk16x_set\, B => 
        tx_packet_complt_intrs, C => un6_apb3_reset_rs, Y => 
        tx_packet_complt_int_net_1);
    
    \rx_FIFO_UNDERRUN_int\ : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => \un23_int_reg_clr\, ALn => un2_apb3_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => rx_FIFO_UNDERRUN_intrs);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity uP_if is

    port( up_EOP_del                    : out   std_logic_vector(5 downto 0);
          int_reg                       : out   std_logic_vector(7 downto 1);
          RX_FIFO_DOUT                  : in    std_logic_vector(8 downto 0);
          CoreAPB3_0_APBmslave0_PADDR   : in    std_logic_vector(7 downto 0);
          RX_packet_depth               : out   std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PRDATA  : out   std_logic_vector(7 downto 0);
          consumer_type4_reg            : out   std_logic_vector(9 downto 0);
          consumer_type3_reg            : out   std_logic_vector(9 downto 0);
          consumer_type2_reg            : out   std_logic_vector(9 downto 0);
          consumer_type1_reg            : out   std_logic_vector(9 downto 0);
          CoreAPB3_0_APBmslave0_PWDATA  : in    std_logic_vector(7 downto 0);
          up_EOP_sync                   : out   std_logic_vector(2 downto 1);
          control_reg_0                 : out   std_logic;
          control_reg_2                 : out   std_logic;
          control_reg_3                 : out   std_logic;
          block_int_until_rd            : out   std_logic;
          RESET_i                       : in    std_logic;
          tx_packet_complt              : in    std_logic;
          rx_CRC_error_set              : in    std_logic;
          rx_CRC_error_int              : out   std_logic;
          un31_int_reg_clr              : out   std_logic;
          rx_CRC_error                  : in    std_logic;
          RX_FIFO_OVERFLOW_set          : in    std_logic;
          rx_FIFO_OVERFLOW_int          : out   std_logic;
          un27_int_reg_clr              : out   std_logic;
          RX_FIFO_OVERFLOW              : in    std_logic;
          RX_FIFO_UNDERRUN_set          : in    std_logic;
          rx_FIFO_UNDERRUN_int          : out   std_logic;
          un23_int_reg_clr              : out   std_logic;
          RX_FIFO_UNDERRUN              : in    std_logic;
          TX_FIFO_OVERFLOW_set          : in    std_logic;
          un19_int_reg_clr              : out   std_logic;
          TX_FIFO_OVERFLOW              : in    std_logic;
          TX_FIFO_UNDERRUN_set          : in    std_logic;
          un15_int_reg_clr              : out   std_logic;
          TX_FIFO_UNDERRUN              : in    std_logic;
          int_reg_clr                   : out   std_logic;
          RESET                         : in    std_logic;
          CommsFPGA_top_0_INT           : out   std_logic;
          TX_PreAmble                   : in    std_logic;
          N_480_i                       : out   std_logic;
          CoreAPB3_0_APBmslave0_PWRITE  : in    std_logic;
          RX_FIFO_Empty                 : in    std_logic;
          RX_FIFO_Full                  : in    std_logic;
          CoreAPB3_0_APBmslave0_PENABLE : in    std_logic;
          CoreAPB3_0_APBmslave0_PSELx   : in    std_logic;
          TX_FIFO_Empty                 : in    std_logic;
          TX_FIFO_Full                  : in    std_logic;
          rx_packet_avail_int           : out   std_logic;
          rx_packet_complt              : in    std_logic;
          RX_packet_depth_status        : out   std_logic;
          TX_FIFO_wr_en                 : out   std_logic;
          RX_FIFO_rd_en                 : out   std_logic;
          N_480_i_i                     : in    std_logic;
          TX_FIFO_RST                   : out   std_logic;
          rx_FIFO_rst_reg               : out   std_logic;
          start_tx_FIFO                 : out   std_logic;
          internal_loopback             : out   std_logic;
          external_loopback             : out   std_logic;
          long_reset                    : in    std_logic;
          CoreAPB3_0_APBmslave0_PREADY  : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz     : in    std_logic;
          long_reset_set                : in    std_logic;
          iup_EOP                       : out   std_logic;
          CommsFPGA_CCC_0_GL0           : in    std_logic;
          long_reset_i                  : in    std_logic
        );

end uP_if;

architecture DEF_ARCH of uP_if is 

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component Interrupts
    port( CoreAPB3_0_APBmslave0_PADDR  : in    std_logic_vector(3 downto 2) := (others => 'U');
          CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 1) := (others => 'U');
          int_reg                      : out   std_logic_vector(7 downto 1);
          i_int_mask_reg               : in    std_logic_vector(7 downto 1) := (others => 'U');
          up_EOP_del                   : out   std_logic_vector(5 downto 0);
          N_218                        : in    std_logic := 'U';
          write_reg_en                 : in    std_logic := 'U';
          CommsFPGA_top_0_INT          : out   std_logic;
          RESET                        : in    std_logic := 'U';
          int_reg_clr                  : out   std_logic;
          long_reset                   : in    std_logic := 'U';
          RX_packet_depth_status       : in    std_logic := 'U';
          tx_packet_complt_int         : out   std_logic;
          TX_FIFO_UNDERRUN             : in    std_logic := 'U';
          un15_int_reg_clr             : out   std_logic;
          TX_FIFO_UNDERRUN_set         : in    std_logic := 'U';
          TX_FIFO_OVERFLOW             : in    std_logic := 'U';
          un19_int_reg_clr             : out   std_logic;
          TX_FIFO_OVERFLOW_set         : in    std_logic := 'U';
          RX_FIFO_UNDERRUN             : in    std_logic := 'U';
          un23_int_reg_clr             : out   std_logic;
          rx_FIFO_UNDERRUN_int         : out   std_logic;
          RX_FIFO_UNDERRUN_set         : in    std_logic := 'U';
          RX_FIFO_OVERFLOW             : in    std_logic := 'U';
          un27_int_reg_clr             : out   std_logic;
          rx_FIFO_OVERFLOW_int         : out   std_logic;
          RX_FIFO_OVERFLOW_set         : in    std_logic := 'U';
          rx_CRC_error                 : in    std_logic := 'U';
          un31_int_reg_clr             : out   std_logic;
          rx_CRC_error_int             : out   std_logic;
          rx_CRC_error_set             : in    std_logic := 'U';
          rx_packet_avail_int          : out   std_logic;
          tx_packet_complt             : in    std_logic := 'U';
          iup_EOP                      : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0          : in    std_logic := 'U';
          RESET_i                      : in    std_logic := 'U';
          block_int_until_rd           : out   std_logic
        );
  end component;

    signal \iAPB3_READY[0]_net_1\, \iAPB3_READY_i[0]\, 
        \up_EOP_sync[0]_net_1\, VCC_net_1, iup_EOP_net_1, 
        GND_net_1, \up_EOP_sync[1]_net_1\, \up_EOP_sync[2]_net_1\, 
        \iAPB3_READYrs[0]\, un5_apb3_rst_rs, un5_apb3_rst_i, 
        CoreAPB3_0_APBmslave0_PREADYrs, 
        \CoreAPB3_0_APBmslave0_PREADY\, 
        \mac_3_byte_4_reg[7]_net_1\, un13_mac_3_byte_4_reg_en, 
        \mac_3_byte_3_reg[0]_net_1\, un13_mac_3_byte_3_reg_en, 
        \mac_3_byte_3_reg[1]_net_1\, \mac_3_byte_3_reg[2]_net_1\, 
        \mac_3_byte_3_reg[3]_net_1\, \mac_3_byte_3_reg[4]_net_1\, 
        \mac_3_byte_3_reg[5]_net_1\, \mac_3_byte_3_reg[6]_net_1\, 
        \mac_3_byte_3_reg[7]_net_1\, \mac_3_byte_5_reg[0]_net_1\, 
        un13_mac_3_byte_5_reg_en, \mac_3_byte_5_reg[1]_net_1\, 
        \mac_3_byte_5_reg[2]_net_1\, \mac_3_byte_5_reg[3]_net_1\, 
        \mac_3_byte_5_reg[4]_net_1\, \mac_3_byte_5_reg[5]_net_1\, 
        \mac_3_byte_5_reg[6]_net_1\, \mac_3_byte_5_reg[7]_net_1\, 
        \mac_3_byte_4_reg[0]_net_1\, \mac_3_byte_4_reg[1]_net_1\, 
        \mac_3_byte_4_reg[2]_net_1\, \mac_3_byte_4_reg[3]_net_1\, 
        \mac_3_byte_4_reg[4]_net_1\, \mac_3_byte_4_reg[5]_net_1\, 
        \mac_3_byte_4_reg[6]_net_1\, \mac_4_byte_1_reg[1]_net_1\, 
        un13_mac_4_byte_1_reg_en, \mac_4_byte_1_reg[2]_net_1\, 
        \mac_4_byte_1_reg[3]_net_1\, \mac_4_byte_1_reg[4]_net_1\, 
        \mac_4_byte_1_reg[5]_net_1\, \mac_4_byte_1_reg[6]_net_1\, 
        \mac_4_byte_1_reg[7]_net_1\, \mac_3_byte_6_reg[0]_net_1\, 
        un13_mac_3_byte_6_reg_en, \mac_3_byte_6_reg[1]_net_1\, 
        \mac_3_byte_6_reg[2]_net_1\, \mac_3_byte_6_reg[3]_net_1\, 
        \mac_3_byte_6_reg[4]_net_1\, \mac_3_byte_6_reg[5]_net_1\, 
        \mac_3_byte_6_reg[6]_net_1\, \mac_3_byte_6_reg[7]_net_1\, 
        \mac_4_byte_3_reg[2]_net_1\, un13_mac_4_byte_3_reg_en, 
        \mac_4_byte_3_reg[3]_net_1\, \mac_4_byte_3_reg[4]_net_1\, 
        \mac_4_byte_3_reg[5]_net_1\, \mac_4_byte_3_reg[6]_net_1\, 
        \mac_4_byte_3_reg[7]_net_1\, \mac_4_byte_2_reg[0]_net_1\, 
        un13_mac_4_byte_2_reg_en, \mac_4_byte_2_reg[1]_net_1\, 
        \mac_4_byte_2_reg[2]_net_1\, \mac_4_byte_2_reg[3]_net_1\, 
        \mac_4_byte_2_reg[4]_net_1\, \mac_4_byte_2_reg[5]_net_1\, 
        \mac_4_byte_2_reg[6]_net_1\, \mac_4_byte_2_reg[7]_net_1\, 
        \mac_4_byte_1_reg[0]_net_1\, \mac_4_byte_5_reg[3]_net_1\, 
        un13_mac_4_byte_5_reg_en, \mac_4_byte_5_reg[4]_net_1\, 
        \mac_4_byte_5_reg[5]_net_1\, \mac_4_byte_5_reg[6]_net_1\, 
        \mac_4_byte_5_reg[7]_net_1\, \mac_4_byte_4_reg[0]_net_1\, 
        un13_mac_4_byte_4_reg_en, \mac_4_byte_4_reg[1]_net_1\, 
        \mac_4_byte_4_reg[2]_net_1\, \mac_4_byte_4_reg[3]_net_1\, 
        \mac_4_byte_4_reg[4]_net_1\, \mac_4_byte_4_reg[5]_net_1\, 
        \mac_4_byte_4_reg[6]_net_1\, \mac_4_byte_4_reg[7]_net_1\, 
        \mac_4_byte_3_reg[0]_net_1\, \mac_4_byte_3_reg[1]_net_1\, 
        \mac_1_byte_1_reg[4]_net_1\, un13_mac_1_byte_1_reg_en, 
        \mac_1_byte_1_reg[5]_net_1\, \mac_1_byte_1_reg[6]_net_1\, 
        \mac_1_byte_1_reg[7]_net_1\, \scratch_pad_reg[0]_net_1\, 
        \write_scratch_reg_en\, \scratch_pad_reg[1]_net_1\, 
        \scratch_pad_reg[2]_net_1\, \scratch_pad_reg[3]_net_1\, 
        \scratch_pad_reg[4]_net_1\, \scratch_pad_reg[5]_net_1\, 
        \scratch_pad_reg[6]_net_1\, \scratch_pad_reg[7]_net_1\, 
        \mac_4_byte_5_reg[0]_net_1\, \mac_4_byte_5_reg[1]_net_1\, 
        \mac_4_byte_5_reg[2]_net_1\, \mac_1_byte_3_reg[5]_net_1\, 
        un13_mac_1_byte_3_reg_en, \mac_1_byte_3_reg[6]_net_1\, 
        \mac_1_byte_3_reg[7]_net_1\, \consumer_type1_reg[0]\, 
        un13_mac_1_byte_2_reg_en, \consumer_type1_reg[1]\, 
        \consumer_type1_reg[2]\, \consumer_type1_reg[3]\, 
        \consumer_type1_reg[4]\, \consumer_type1_reg[5]\, 
        \consumer_type1_reg[6]\, \consumer_type1_reg[7]\, 
        \consumer_type1_reg[8]\, \consumer_type1_reg[9]\, 
        \mac_1_byte_1_reg[2]_net_1\, \mac_1_byte_1_reg[3]_net_1\, 
        \mac_1_byte_5_reg[6]_net_1\, un13_mac_1_byte_5_reg_en, 
        \mac_1_byte_5_reg[7]_net_1\, \consumer_type2_reg[0]\, 
        un13_mac_1_byte_4_reg_en, \consumer_type2_reg[1]\, 
        \consumer_type2_reg[2]\, \consumer_type2_reg[3]\, 
        \consumer_type2_reg[4]\, \consumer_type2_reg[5]\, 
        \consumer_type2_reg[6]\, \consumer_type2_reg[7]\, 
        \consumer_type2_reg[8]\, \consumer_type2_reg[9]\, 
        \mac_1_byte_3_reg[2]_net_1\, \mac_1_byte_3_reg[3]_net_1\, 
        \mac_1_byte_3_reg[4]_net_1\, \mac_2_byte_1_reg[7]_net_1\, 
        un13_mac_2_byte_1_reg_en, \consumer_type3_reg[0]\, 
        un13_mac_1_byte_6_reg_en, \consumer_type3_reg[1]\, 
        \consumer_type3_reg[2]\, \consumer_type3_reg[3]\, 
        \consumer_type3_reg[4]\, \consumer_type3_reg[5]\, 
        \consumer_type3_reg[6]\, \consumer_type3_reg[7]\, 
        \consumer_type3_reg[8]\, \consumer_type3_reg[9]\, 
        \mac_1_byte_5_reg[2]_net_1\, \mac_1_byte_5_reg[3]_net_1\, 
        \mac_1_byte_5_reg[4]_net_1\, \mac_1_byte_5_reg[5]_net_1\, 
        \consumer_type4_reg[0]\, un13_mac_2_byte_2_reg_en, 
        \consumer_type4_reg[1]\, \consumer_type4_reg[2]\, 
        \consumer_type4_reg[3]\, \consumer_type4_reg[4]\, 
        \consumer_type4_reg[5]\, \consumer_type4_reg[6]\, 
        \consumer_type4_reg[7]\, \consumer_type4_reg[8]\, 
        \consumer_type4_reg[9]\, \mac_2_byte_1_reg[2]_net_1\, 
        \mac_2_byte_1_reg[3]_net_1\, \mac_2_byte_1_reg[4]_net_1\, 
        \mac_2_byte_1_reg[5]_net_1\, \mac_2_byte_1_reg[6]_net_1\, 
        \mac_2_byte_4_reg[1]_net_1\, un13_mac_2_byte_4_reg_en, 
        \mac_2_byte_4_reg[2]_net_1\, \mac_2_byte_4_reg[3]_net_1\, 
        \mac_2_byte_4_reg[4]_net_1\, \mac_2_byte_4_reg[5]_net_1\, 
        \mac_2_byte_4_reg[6]_net_1\, \mac_2_byte_4_reg[7]_net_1\, 
        \mac_2_byte_3_reg[0]_net_1\, un13_mac_2_byte_3_reg_en, 
        \mac_2_byte_3_reg[1]_net_1\, \mac_2_byte_3_reg[2]_net_1\, 
        \mac_2_byte_3_reg[3]_net_1\, \mac_2_byte_3_reg[4]_net_1\, 
        \mac_2_byte_3_reg[5]_net_1\, \mac_2_byte_3_reg[6]_net_1\, 
        \mac_2_byte_3_reg[7]_net_1\, \mac_2_byte_6_reg[2]_net_1\, 
        un13_mac_2_byte_6_reg_en, \mac_2_byte_6_reg[3]_net_1\, 
        \mac_2_byte_6_reg[4]_net_1\, \mac_2_byte_6_reg[5]_net_1\, 
        \mac_2_byte_6_reg[6]_net_1\, \mac_2_byte_6_reg[7]_net_1\, 
        \mac_2_byte_5_reg[0]_net_1\, un13_mac_2_byte_5_reg_en, 
        \mac_2_byte_5_reg[1]_net_1\, \mac_2_byte_5_reg[2]_net_1\, 
        \mac_2_byte_5_reg[3]_net_1\, \mac_2_byte_5_reg[4]_net_1\, 
        \mac_2_byte_5_reg[5]_net_1\, \mac_2_byte_5_reg[6]_net_1\, 
        \mac_2_byte_5_reg[7]_net_1\, \mac_2_byte_4_reg[0]_net_1\, 
        \mac_3_byte_2_reg[3]_net_1\, un13_mac_3_byte_2_reg_en, 
        \mac_3_byte_2_reg[4]_net_1\, \mac_3_byte_2_reg[5]_net_1\, 
        \mac_3_byte_2_reg[6]_net_1\, \mac_3_byte_2_reg[7]_net_1\, 
        \mac_3_byte_1_reg[0]_net_1\, un13_mac_3_byte_1_reg_en, 
        \mac_3_byte_1_reg[1]_net_1\, \mac_3_byte_1_reg[2]_net_1\, 
        \mac_3_byte_1_reg[3]_net_1\, \mac_3_byte_1_reg[4]_net_1\, 
        \mac_3_byte_1_reg[5]_net_1\, \mac_3_byte_1_reg[6]_net_1\, 
        \mac_3_byte_1_reg[7]_net_1\, \mac_2_byte_6_reg[0]_net_1\, 
        \mac_2_byte_6_reg[1]_net_1\, \i_int_mask_reg[4]_net_1\, 
        un13_int_mask_reg_en_i_i_a2, \i_int_mask_reg[5]_net_1\, 
        \i_int_mask_reg[6]_net_1\, \i_int_mask_reg[7]_net_1\, 
        \mac_4_byte_6_reg[0]_net_1\, un13_mac_4_byte_6_reg_en, 
        \mac_4_byte_6_reg[1]_net_1\, \mac_4_byte_6_reg[2]_net_1\, 
        \mac_4_byte_6_reg[3]_net_1\, \mac_4_byte_6_reg[4]_net_1\, 
        \mac_4_byte_6_reg[5]_net_1\, \mac_4_byte_6_reg[6]_net_1\, 
        \mac_4_byte_6_reg[7]_net_1\, \mac_3_byte_2_reg[0]_net_1\, 
        \mac_3_byte_2_reg[1]_net_1\, \mac_3_byte_2_reg[2]_net_1\, 
        \control_reg_0\, control_reg_22, \external_loopback\, 
        \control_reg_2\, \control_reg_3\, \internal_loopback\, 
        \start_tx_FIFO\, N_456_i, un1_control_reg_en_2_i_0, 
        \rx_FIFO_rst_reg\, \TX_FIFO_RST\, 
        \i_int_mask_reg[0]_net_1\, \i_int_mask_reg[1]_net_1\, 
        \i_int_mask_reg[2]_net_1\, \i_int_mask_reg[3]_net_1\, 
        \mac_4_byte_5_reg_en\, mac_4_byte_6_reg_en_1, N_363, 
        \mac_4_byte_4_reg_en\, N_362, \mac_4_byte_3_reg_en\, 
        N_361, N_479_i_i, N_336, un1_apb3_addr, 
        \mac_3_byte_2_reg_en\, N_354, \mac_3_byte_1_reg_en\, 
        N_353, \mac_2_byte_6_reg_en\, N_352, 
        \mac_2_byte_5_reg_en\, N_351, \mac_2_byte_4_reg_en\, 
        N_350, \mac_2_byte_3_reg_en\, N_349, 
        \mac_2_byte_2_reg_en\, N_348, \mac_3_byte_3_reg_en\, 
        N_355, \mac_3_byte_4_reg_en\, N_356, 
        \mac_3_byte_5_reg_en\, N_357, \mac_3_byte_6_reg_en\, 
        N_358, \mac_4_byte_1_reg_en\, N_359, 
        \mac_4_byte_2_reg_en\, N_360, \mac_4_byte_6_reg_en\, 
        N_364, N_813, N_804, N_812, N_803, \mac_1_byte_2_reg_en\, 
        N_342, \control_reg_en\, N_337, \mac_1_byte_4_reg_en\, 
        N_344, \mac_1_byte_6_reg_en\, N_346, \int_mask_reg_en\, 
        N_339, \mac_1_byte_5_reg_en\, N_345, 
        \mac_1_byte_1_reg_en\, N_341, N_335, 
        \mac_2_byte_1_reg_en\, N_347, \mac_1_byte_3_reg_en\, 
        N_343, \read_reg_en\, \write_reg_en\, un116_apb3_addr, 
        RX_packet_depth_status_net_1, rx_packet_depth_status2, 
        \APB3_RDATA_31_sqmuxa_i\, \APB3_RDATA_1[0]_net_1\, 
        \APB3_RDATA_1[1]\, \APB3_RDATA_1[2]\, 
        \APB3_RDATA_1[3]_net_1\, \APB3_RDATA_1[4]\, 
        \APB3_RDATA_1[5]\, \APB3_RDATA_1[6]_net_1\, 
        \APB3_RDATA_1[7]_net_1\, \RX_packet_depth[0]_net_1\, 
        \RX_packet_depth_s[0]\, N_1528_i, 
        \RX_packet_depth[1]_net_1\, \RX_packet_depth_s[1]\, 
        \RX_packet_depth[2]_net_1\, \RX_packet_depth_s[2]\, 
        \RX_packet_depth[3]_net_1\, \RX_packet_depth_s[3]\, 
        \RX_packet_depth[4]_net_1\, \RX_packet_depth_s[4]\, 
        \RX_packet_depth[5]_net_1\, \RX_packet_depth_s[5]\, 
        \RX_packet_depth[6]_net_1\, \RX_packet_depth_s[6]\, 
        \RX_packet_depth[7]_net_1\, \RX_packet_depth_s[7]_net_1\, 
        un12_mac_2_byte_1_reg_en_16_0_reto, 
        un12_mac_2_byte_1_reg_en_16_0, 
        un12_mac_2_byte_1_reg_en_16_1_reto, 
        un12_mac_2_byte_1_reg_en_16_1, 
        un12_mac_2_byte_1_reg_en_16_2_reto, 
        un12_mac_2_byte_1_reg_en_16_2, N_342_reto, 
        mac_4_byte_6_reg_en_1_reto, mac_1_byte_2_reg_en_reto, 
        N_341_reto, N_803_reto, mac_4_byte_6_reg_en_1_reto_0, 
        mac_1_byte_1_reg_en_reto, RX_packet_depth_s_914_FCO, 
        \RX_packet_depth_cry[0]_net_1\, 
        \RX_packet_depth_cry[1]_net_1\, 
        \RX_packet_depth_cry[2]_net_1\, 
        \RX_packet_depth_cry[3]_net_1\, 
        \RX_packet_depth_cry[4]_net_1\, 
        \RX_packet_depth_cry[5]_net_1\, 
        \RX_packet_depth_cry[6]_net_1\, APB3_RDATA_1_sn_i6_mux, 
        \APB3_RDATA_1_sn_m19_2\, APB3_RDATA_1_sn_N_18, 
        APB3_RDATA_1_sn_m19_4_1_0_y0, 
        APB3_RDATA_1_sn_m19_4_1_0_co0, \APB3_RDATA_1_sn_m19_0\, 
        \APB3_RDATA_1_25_0_wmux_0_Y[5]\, 
        \APB3_RDATA_1_25_0_0_y0[5]\, \APB3_RDATA_1_25_0_0_co0[5]\, 
        \APB3_RDATA_1_25_0_wmux_0_Y[4]\, 
        \APB3_RDATA_1_25_0_0_y0[4]\, \APB3_RDATA_1_25_0_0_co0[4]\, 
        \APB3_RDATA_1_25_0_wmux_0_Y[3]\, 
        \APB3_RDATA_1_25_0_0_y0[3]\, \APB3_RDATA_1_25_0_0_co0[3]\, 
        \APB3_RDATA_1_25_0_wmux_0_Y[2]\, 
        \APB3_RDATA_1_25_0_0_y0[2]\, \APB3_RDATA_1_25_0_0_co0[2]\, 
        \APB3_RDATA_1_25_0_wmux_0_Y[1]\, 
        \APB3_RDATA_1_25_0_0_y0[1]\, \APB3_RDATA_1_25_0_0_co0[1]\, 
        \APB3_RDATA_1_25_0_wmux_0_Y[0]\, 
        \APB3_RDATA_1_25_0_0_y0[0]\, \APB3_RDATA_1_25_0_0_co0[0]\, 
        \APB3_RDATA_1_25_0_wmux_0_Y[6]\, 
        \APB3_RDATA_1_25_0_0_y0[6]\, \APB3_RDATA_1_25_0_0_co0[6]\, 
        N_1687, \APB3_RDATA_1_17_0_0_y0[7]\, 
        \APB3_RDATA_1_17_0_0_co0[7]\, N_1718, 
        \APB3_RDATA_1_21_0_0_y0[6]\, \APB3_RDATA_1_21_0_0_co0[6]\, 
        N_120, \APB3_RDATA_1_18_0_0_y0[4]\, 
        \APB3_RDATA_1_18_0_0_co0[4]\, N_1714, 
        \APB3_RDATA_1_21_0_0_y0[2]\, \APB3_RDATA_1_21_0_0_co0[2]\, 
        N_1682, \APB3_RDATA_1_17_0_0_y0[2]\, 
        \APB3_RDATA_1_17_0_0_co0[2]\, N_1703, 
        \APB3_RDATA_1_19_0_0_y0[7]\, \APB3_RDATA_1_19_0_0_co0[7]\, 
        N_1698, \APB3_RDATA_1_19_0_0_y0[2]\, 
        \APB3_RDATA_1_19_0_0_co0[2]\, N_1719, 
        \APB3_RDATA_1_21_0_0_y0[7]\, \APB3_RDATA_1_21_0_0_co0[7]\, 
        N_1716, \APB3_RDATA_1_21_0_0_y0[4]\, 
        \APB3_RDATA_1_21_0_0_co0[4]\, N_1712, 
        \APB3_RDATA_1_21_0_0_y0[0]\, \APB3_RDATA_1_21_0_0_co0[0]\, 
        N_123, \APB3_RDATA_1_18_0_0_y0[7]\, 
        \APB3_RDATA_1_18_0_0_co0[7]\, N_121, 
        \APB3_RDATA_1_18_0_0_y0[5]\, \APB3_RDATA_1_18_0_0_co0[5]\, 
        N_118, \APB3_RDATA_1_18_0_0_y0[2]\, 
        \APB3_RDATA_1_18_0_0_co0[2]\, N_117, 
        \APB3_RDATA_1_18_0_0_y0[1]\, \APB3_RDATA_1_18_0_0_co0[1]\, 
        N_116, \APB3_RDATA_1_18_0_0_y0[0]\, 
        \APB3_RDATA_1_18_0_0_co0[0]\, N_1686, 
        \APB3_RDATA_1_17_0_0_y0[6]\, \APB3_RDATA_1_17_0_0_co0[6]\, 
        N_1685, \APB3_RDATA_1_17_0_0_y0[5]\, 
        \APB3_RDATA_1_17_0_0_co0[5]\, N_1684, 
        \APB3_RDATA_1_17_0_0_y0[4]\, \APB3_RDATA_1_17_0_0_co0[4]\, 
        N_1681, \APB3_RDATA_1_17_0_0_y0[1]\, 
        \APB3_RDATA_1_17_0_0_co0[1]\, N_1680, 
        \APB3_RDATA_1_17_0_0_y0[0]\, \APB3_RDATA_1_17_0_0_co0[0]\, 
        N_1717, \APB3_RDATA_1_21_0_0_y0[5]\, 
        \APB3_RDATA_1_21_0_0_co0[5]\, N_1715, 
        \APB3_RDATA_1_21_0_0_y0[3]\, \APB3_RDATA_1_21_0_0_co0[3]\, 
        N_1701, \APB3_RDATA_1_19_0_0_y0[5]\, 
        \APB3_RDATA_1_19_0_0_co0[5]\, N_1700, 
        \APB3_RDATA_1_19_0_0_y0[4]\, \APB3_RDATA_1_19_0_0_co0[4]\, 
        N_1699, \APB3_RDATA_1_19_0_0_y0[3]\, 
        \APB3_RDATA_1_19_0_0_co0[3]\, N_1696, 
        \APB3_RDATA_1_19_0_0_y0[0]\, \APB3_RDATA_1_19_0_0_co0[0]\, 
        N_1683, \APB3_RDATA_1_17_0_0_y0[3]\, 
        \APB3_RDATA_1_17_0_0_co0[3]\, N_1713, 
        \APB3_RDATA_1_21_0_0_y0[1]\, \APB3_RDATA_1_21_0_0_co0[1]\, 
        N_1702, \APB3_RDATA_1_19_0_0_y0[6]\, 
        \APB3_RDATA_1_19_0_0_co0[6]\, N_1697, 
        \APB3_RDATA_1_19_0_0_y0[1]\, \APB3_RDATA_1_19_0_0_co0[1]\, 
        N_119, \APB3_RDATA_1_18_0_0_y0[3]\, 
        \APB3_RDATA_1_18_0_0_co0[3]\, N_122, 
        \APB3_RDATA_1_18_0_0_y0[6]\, \APB3_RDATA_1_18_0_0_co0[6]\, 
        \APB3_RDATA_1_27_d_0_wmux_0_Y[3]\, 
        APB3_RDATA_1_sn_N_31_mux, N_1577, N_1659, 
        \APB3_RDATA_1_27_d_0_0_y0[3]\, 
        \APB3_RDATA_1_27_d_0_0_co0[3]\, \int_reg[3]\, N_1752, 
        \APB3_RDATA_1_25_4_0_y1[7]\, \APB3_RDATA_1_25_4_0_y3[7]\, 
        \APB3_RDATA_1_25_4_co1_0[7]\, N_57, N_1571, 
        \APB3_RDATA_1_25_4_y0_0[7]\, \APB3_RDATA_1_25_4_co0_0[7]\, 
        \APB3_RDATA_1_25_4_0_co1[7]\, \APB3_RDATA_1_25_4_0_y0[7]\, 
        \APB3_RDATA_1_25_4_0_co0[7]\, N_55, N_1569, 
        \APB3_RDATA_1_25_3[5]_net_1\, N_562, N_1568, 
        \APB3_RDATA_1_25_3[4]_net_1\, N_561, N_1567, 
        \APB3_RDATA_1_25_3[3]_net_1\, N_560, N_1566, 
        \APB3_RDATA_1_25_3[2]_net_1\, N_559, N_1565, 
        \APB3_RDATA_1_25_3[1]_net_1\, N_558, N_1564, 
        \APB3_RDATA_1_25_3[0]_net_1\, N_56, N_1570, 
        \APB3_RDATA_1_25_3[6]_net_1\, \N_455_i\, 
        APB3_RDATA_1_sn_N_10, N_3, \rx_packet_avail_int\, 
        \APB3_RDATA_1_27_d_0[6]_net_1\, tx_packet_complt_int, 
        N_1671, N_413, N_157, \APB3_RDATA_1_bm[1]_net_1\, 
        \APB3_RDATA_1_ns_1[1]_net_1\, N_1730, 
        APB3_RDATA_1_sn_N_33_mux, APB3_RDATA_1_sn_N_32_mux, 
        \APB3_RDATA_1_am_1[1]_net_1\, \APB3_RDATA_1_d_0[0]_net_1\, 
        \APB3_RDATA_1_1[0]_net_1\, \APB3_RDATA_1_1_0[0]_net_1\, 
        N_1753, N_1720, N_1738, APB3_RDATA_1_sn_N_14, N_1746, 
        \APB3_RDATA_1_4\, \APB3_RDATA_1_1[7]_net_1\, N_1760, 
        \APB3_RDATA_1_0_1[7]_net_1\, \APB3_RDATA_1_bm_1[2]_net_1\, 
        N_1731, \APB3_RDATA_1_bm[2]_net_1\, N_1576, N_1658, 
        APB3_RDATA_1_sn_m8_out, \APB3_RDATA_1_bm_1[5]_net_1\, 
        \APB3_RDATA_1_bm[5]_net_1\, \int_reg[5]\, 
        \APB3_RDATA_1_bm_1[4]_net_1\, N_1733, 
        \APB3_RDATA_1_bm[4]_net_1\, N_1578, N_1660, N_1805, 
        \APB3_RDATA_31_sqmuxa_i_1\, 
        \APB3_RDATA_31_sqmuxa_1_a3_0_2\, 
        \APB3_RDATA_1_29_d_am_1_0[5]_net_1\, 
        \APB3_RDATA_1_29_d_am[5]_net_1\, 
        \APB3_RDATA_1_29_d_1[6]_net_1\, 
        \APB3_RDATA_1_29_d[6]_net_1\, 
        \APB3_RDATA_1_22_1_0[7]_net_1\, N_1727, 
        \APB3_RDATA_1_27_d_3_1[6]_net_1\, 
        \APB3_RDATA_1_27_d_3[6]_net_1\, 
        \APB3_RDATA_1_29_d_ns[5]_net_1\, 
        \APB3_RDATA_1_ns_1[5]_net_1\, N_1777, 
        \APB3_RDATA_1_s[7]_net_1\, \APB3_RDATA_1_am[2]_net_1\, 
        \APB3_RDATA_1_am[4]_net_1\, \APB3_RDATA_1_d_bm[3]_net_1\, 
        \APB3_RDATA_1_d_am[3]_net_1\, 
        \APB3_RDATA_1_d_ns[3]_net_1\, 
        \APB3_RDATA_1_29_d_bm[5]_net_1\, 
        \APB3_RDATA_1_22_am[0]_net_1\, 
        \APB3_RDATA_1_22_bm[0]_net_1\, 
        \APB3_RDATA_1_22_am[1]_net_1\, 
        \APB3_RDATA_1_22_bm[1]_net_1\, N_1721, 
        \APB3_RDATA_1_27_d_1[6]_net_1\, 
        \APB3_RDATA_1_d_RNO[6]_net_1\, N_1750, N_1749, N_1748, 
        N_1747, N_1745, N_1751, \APB3_RDATA_1_29_s[6]_net_1\, 
        N_1744, N_802, un13_mac_4_byte_5_reg_en_0_a2_0_a2_0, 
        N_796, un1_control_reg_en_2_i_0_0_o2_0, N_201, N_202, 
        N_212, APB3_RDATA_1_sn_N_23, N_1757, N_1755, N_1754, 
        N_1743, N_1742, N_1741, N_1740, N_1739, N_1737, 
        un13_mac_4_byte_3_reg_en_0_a2_4_a2_2, 
        un13_mac_4_byte_4_reg_en_0_a2_0_a2_1, 
        un105_apb3_addr_0_a2_0_1, un1_RX_packet_depthlto7_5, 
        un1_RX_packet_depthlto7_4, N_407, 
        un13_mac_4_byte_2_reg_en_0_a2_3_o2_0, N_412, N_156, N_129, 
        \int_reg[4]\, N_1668, \int_reg[2]\, N_1666, \int_reg[1]\, 
        N_1665, N_199, N_200, N_1778, N_1776, N_1774, N_414, 
        N_213, N_218, APB3_RDATA_1_sn_N_25, N_131, 
        \APB3_RDATA_1_d_a0[0]_net_1\, 
        \APB3_RDATA_1_d_a1[0]_net_1\, N_420, 
        \APB3_RDATA_1_0_0[7]_net_1\, 
        un13_mac_4_byte_1_reg_en_0_a2_0_a2_1, N_1765, N_141, N_7, 
        N_10, N_11, N_146, \APB3_RDATA_1_d[6]_net_1\, N_160, 
        N_553, N_801 : std_logic;

    for all : Interrupts
	Use entity work.Interrupts(DEF_ARCH);
begin 

    int_reg(5) <= \int_reg[5]\;
    int_reg(4) <= \int_reg[4]\;
    int_reg(3) <= \int_reg[3]\;
    int_reg(2) <= \int_reg[2]\;
    int_reg(1) <= \int_reg[1]\;
    RX_packet_depth(7) <= \RX_packet_depth[7]_net_1\;
    RX_packet_depth(6) <= \RX_packet_depth[6]_net_1\;
    RX_packet_depth(5) <= \RX_packet_depth[5]_net_1\;
    RX_packet_depth(4) <= \RX_packet_depth[4]_net_1\;
    RX_packet_depth(3) <= \RX_packet_depth[3]_net_1\;
    RX_packet_depth(2) <= \RX_packet_depth[2]_net_1\;
    RX_packet_depth(1) <= \RX_packet_depth[1]_net_1\;
    RX_packet_depth(0) <= \RX_packet_depth[0]_net_1\;
    consumer_type4_reg(9) <= \consumer_type4_reg[9]\;
    consumer_type4_reg(8) <= \consumer_type4_reg[8]\;
    consumer_type4_reg(7) <= \consumer_type4_reg[7]\;
    consumer_type4_reg(6) <= \consumer_type4_reg[6]\;
    consumer_type4_reg(5) <= \consumer_type4_reg[5]\;
    consumer_type4_reg(4) <= \consumer_type4_reg[4]\;
    consumer_type4_reg(3) <= \consumer_type4_reg[3]\;
    consumer_type4_reg(2) <= \consumer_type4_reg[2]\;
    consumer_type4_reg(1) <= \consumer_type4_reg[1]\;
    consumer_type4_reg(0) <= \consumer_type4_reg[0]\;
    consumer_type3_reg(9) <= \consumer_type3_reg[9]\;
    consumer_type3_reg(8) <= \consumer_type3_reg[8]\;
    consumer_type3_reg(7) <= \consumer_type3_reg[7]\;
    consumer_type3_reg(6) <= \consumer_type3_reg[6]\;
    consumer_type3_reg(5) <= \consumer_type3_reg[5]\;
    consumer_type3_reg(4) <= \consumer_type3_reg[4]\;
    consumer_type3_reg(3) <= \consumer_type3_reg[3]\;
    consumer_type3_reg(2) <= \consumer_type3_reg[2]\;
    consumer_type3_reg(1) <= \consumer_type3_reg[1]\;
    consumer_type3_reg(0) <= \consumer_type3_reg[0]\;
    consumer_type2_reg(9) <= \consumer_type2_reg[9]\;
    consumer_type2_reg(8) <= \consumer_type2_reg[8]\;
    consumer_type2_reg(7) <= \consumer_type2_reg[7]\;
    consumer_type2_reg(6) <= \consumer_type2_reg[6]\;
    consumer_type2_reg(5) <= \consumer_type2_reg[5]\;
    consumer_type2_reg(4) <= \consumer_type2_reg[4]\;
    consumer_type2_reg(3) <= \consumer_type2_reg[3]\;
    consumer_type2_reg(2) <= \consumer_type2_reg[2]\;
    consumer_type2_reg(1) <= \consumer_type2_reg[1]\;
    consumer_type2_reg(0) <= \consumer_type2_reg[0]\;
    consumer_type1_reg(9) <= \consumer_type1_reg[9]\;
    consumer_type1_reg(8) <= \consumer_type1_reg[8]\;
    consumer_type1_reg(7) <= \consumer_type1_reg[7]\;
    consumer_type1_reg(6) <= \consumer_type1_reg[6]\;
    consumer_type1_reg(5) <= \consumer_type1_reg[5]\;
    consumer_type1_reg(4) <= \consumer_type1_reg[4]\;
    consumer_type1_reg(3) <= \consumer_type1_reg[3]\;
    consumer_type1_reg(2) <= \consumer_type1_reg[2]\;
    consumer_type1_reg(1) <= \consumer_type1_reg[1]\;
    consumer_type1_reg(0) <= \consumer_type1_reg[0]\;
    up_EOP_sync(2) <= \up_EOP_sync[2]_net_1\;
    up_EOP_sync(1) <= \up_EOP_sync[1]_net_1\;
    control_reg_0 <= \control_reg_0\;
    control_reg_2 <= \control_reg_2\;
    control_reg_3 <= \control_reg_3\;
    rx_packet_avail_int <= \rx_packet_avail_int\;
    RX_packet_depth_status <= RX_packet_depth_status_net_1;
    TX_FIFO_RST <= \TX_FIFO_RST\;
    rx_FIFO_rst_reg <= \rx_FIFO_rst_reg\;
    start_tx_FIFO <= \start_tx_FIFO\;
    internal_loopback <= \internal_loopback\;
    external_loopback <= \external_loopback\;
    CoreAPB3_0_APBmslave0_PREADY <= 
        \CoreAPB3_0_APBmslave0_PREADY\;
    iup_EOP <= iup_EOP_net_1;

    \mac_3_byte_1_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_1_reg[7]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un9_apb3_addr_0_a2_1\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_200, B => APB3_RDATA_1_sn_N_18, Y => N_218);
    
    \mac_2_byte_4_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_4_reg[3]_net_1\);
    
    \APB3_RDATA_1_19_0_wmux_0[7]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_19_0_0_y0[7]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \mac_2_byte_5_reg[7]_net_1\, D => 
        \mac_4_byte_1_reg[7]_net_1\, FCI => 
        \APB3_RDATA_1_19_0_0_co0[7]\, S => OPEN, Y => N_1703, FCO
         => OPEN);
    
    \APB3_RDATA_1_22_am[1]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \consumer_type3_reg[1]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \scratch_pad_reg[1]_net_1\, Y => 
        \APB3_RDATA_1_22_am[1]_net_1\);
    
    \mac_2_byte_3_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_3_reg[4]_net_1\);
    
    \mac_2_byte_2_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type4_reg[3]\);
    
    APB3_RDATA_31_sqmuxa_1_m3 : CFG4
      generic map(INIT => x"AAB8")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(7), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        CoreAPB3_0_APBmslave0_PADDR(5), D => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_1805);
    
    \APB3_RDATA_1_25_3[3]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_561, B => CoreAPB3_0_APBmslave0_PADDR(3), C
         => N_1567, Y => \APB3_RDATA_1_25_3[3]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_4_byte_5_reg_en_0_a2_0_a2\ : CFG4
      generic map(INIT => x"0008")

      port map(A => un13_mac_4_byte_5_reg_en_0_a2_0_a2_0, B => 
        N_553, C => \mac_1_byte_2_reg_en\, D => N_156, Y => 
        un13_mac_4_byte_5_reg_en);
    
    \i_int_mask_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_int_mask_reg_en_i_i_a2, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \i_int_mask_reg[3]_net_1\);
    
    \APB3_RDATA_1_ns_1[5]\ : CFG4
      generic map(INIT => x"5053")

      port map(A => N_1777, B => APB3_RDATA_1_sn_N_32_mux, C => 
        APB3_RDATA_1_sn_N_33_mux, D => APB3_RDATA_1_sn_N_31_mux, 
        Y => \APB3_RDATA_1_ns_1[5]_net_1\);
    
    \APB3_RDATA_1_21_0_0_wmux[2]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_2_byte_4_reg[2]_net_1\, D => 
        \mac_2_byte_6_reg[2]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_21_0_0_y0[2]\, FCO => 
        \APB3_RDATA_1_21_0_0_co0[2]\);
    
    \REG_WRITE_PROC.un13_mac_1_byte_3_reg_en_0_a2_0_a2_0\ : CFG3
      generic map(INIT => x"04")

      port map(A => \mac_1_byte_2_reg_en\, B => N_407, C => 
        \mac_1_byte_1_reg_en\, Y => N_414);
    
    iRX_FIFO_rd_en : SLE
      port map(D => \iAPB3_READY_i[0]\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_336, ALn => N_479_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => RX_FIFO_rd_en);
    
    \mac_3_byte_2_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_2_reg[0]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un97_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"0080")

      port map(A => N_201, B => un105_apb3_addr_0_a2_0_1, C => 
        CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => N_362);
    
    \APB3_RDATA_1_bm[2]\ : CFG3
      generic map(INIT => x"72")

      port map(A => APB3_RDATA_1_sn_N_31_mux, B => 
        \APB3_RDATA_1_bm_1[2]_net_1\, C => N_1731, Y => 
        \APB3_RDATA_1_bm[2]_net_1\);
    
    \i_int_mask_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_int_mask_reg_en_i_i_a2, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \i_int_mask_reg[4]_net_1\);
    
    \mac_2_byte_3_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_3_reg[3]_net_1\);
    
    \mac_2_byte_2_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type4_reg[4]\);
    
    \RX_packet_depth_cry[1]\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \RX_packet_depth[1]_net_1\, B => 
        rx_packet_complt, C => GND_net_1, D => GND_net_1, FCI => 
        \RX_packet_depth_cry[0]_net_1\, S => 
        \RX_packet_depth_s[1]\, Y => OPEN, FCO => 
        \RX_packet_depth_cry[1]_net_1\);
    
    \APB3_RDATA_1_17_0_0_wmux[1]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => \external_loopback\, 
        D => \mac_2_byte_3_reg[1]_net_1\, FCI => VCC_net_1, S => 
        OPEN, Y => \APB3_RDATA_1_17_0_0_y0[1]\, FCO => 
        \APB3_RDATA_1_17_0_0_co0[1]\);
    
    \RX_packet_depth_cry[5]\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \RX_packet_depth[5]_net_1\, B => 
        rx_packet_complt, C => GND_net_1, D => GND_net_1, FCI => 
        \RX_packet_depth_cry[4]_net_1\, S => 
        \RX_packet_depth_s[5]\, Y => OPEN, FCO => 
        \RX_packet_depth_cry[5]_net_1\);
    
    \APB3_RDATA_1_19_0_0_wmux[7]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \i_int_mask_reg[7]_net_1\, D => 
        \mac_1_byte_3_reg[7]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_19_0_0_y0[7]\, FCO => 
        \APB3_RDATA_1_19_0_0_co0[7]\);
    
    \mac_4_byte_5_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_5_reg[7]_net_1\);
    
    \mac_3_byte_3_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_3_reg[0]_net_1\);
    
    \up_EOP_sync[2]\ : SLE
      port map(D => \up_EOP_sync[1]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \up_EOP_sync[2]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_1_byte_5_reg_en_0_a2_1_a2\ : CFG4
      generic map(INIT => x"0200")

      port map(A => \mac_1_byte_5_reg_en\, B => 
        \mac_1_byte_4_reg_en\, C => \mac_1_byte_3_reg_en\, D => 
        N_414, Y => un13_mac_1_byte_5_reg_en);
    
    \WRITE_REGISTER_ENABLE_PROC.apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"4000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_200, D => N_201, Y
         => N_335);
    
    \APB3_RDATA_1_26[4]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_1716, B => N_120, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_1757);
    
    \mac_4_byte_5_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_5_reg[4]_net_1\);
    
    control_reg_en_0 : CFG4
      generic map(INIT => x"7430")

      port map(A => \CoreAPB3_0_APBmslave0_PREADY\, B => N_337, C
         => \control_reg_en\, D => \iAPB3_READY[0]_net_1\, Y => 
        N_3);
    
    \mac_2_byte_2_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type4_reg[2]\);
    
    \APB3_RDATA_1_19_0_0_wmux[4]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \i_int_mask_reg[4]_net_1\, D => 
        \mac_1_byte_3_reg[4]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_19_0_0_y0[4]\, FCO => 
        \APB3_RDATA_1_19_0_0_co0[4]\);
    
    \REG_WRITE_PROC.un13_mac_4_byte_6_reg_en_0_a2_4_o2\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => \mac_4_byte_5_reg_en\, B => 
        \mac_4_byte_4_reg_en\, C => \mac_4_byte_3_reg_en\, D => 
        \mac_4_byte_2_reg_en\, Y => N_157);
    
    \control_reg[5]\ : SLE
      port map(D => N_456_i, CLK => m2s010_som_sb_0_CCC_71MHz, EN
         => un1_control_reg_en_2_i_0, ALn => long_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \start_tx_FIFO\);
    
    \mac_2_byte_3_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_3_reg[2]_net_1\);
    
    \mac_3_byte_5_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_5_reg[3]_net_1\);
    
    mac_1_byte_3_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_343, ALn => N_480_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_1_byte_3_reg_en\);
    
    \APB3_RDATA_1_25_0_wmux_0[3]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_25_0_0_y0[3]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_1_reg[3]_net_1\, D => 
        \mac_3_byte_3_reg[3]_net_1\, FCI => 
        \APB3_RDATA_1_25_0_0_co0[3]\, S => OPEN, Y => 
        \APB3_RDATA_1_25_0_wmux_0_Y[3]\, FCO => OPEN);
    
    \mac_4_byte_6_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_6_reg[6]_net_1\);
    
    mac_4_byte_6_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_364, ALn => N_480_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_4_byte_6_reg_en\);
    
    \APB3_RDATA_1_28[4]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => N_1741, B => APB3_RDATA_1_sn_N_14, C => 
        N_1749, Y => N_1776);
    
    \APB3_RDATA_1_27_d_0[6]\ : CFG4
      generic map(INIT => x"F202")

      port map(A => \rx_packet_avail_int\, B => 
        \i_int_mask_reg[6]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => 
        CoreAPB3_0_APBmslave0_PADDR(6), Y => 
        \APB3_RDATA_1_27_d_0[6]_net_1\);
    
    \mac_3_byte_5_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_5_reg[6]_net_1\);
    
    \mac_1_byte_5_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type3_reg[8]\);
    
    \mac_2_byte_5_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_5_reg[2]_net_1\);
    
    \APB3_RDATA_1_3[6]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \consumer_type4_reg[6]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_4_reg[6]_net_1\, Y => N_1570);
    
    mac_1_byte_2_reg_en_ret_1 : SLE
      port map(D => N_342, CLK => m2s010_som_sb_0_CCC_71MHz, EN
         => VCC_net_1, ALn => N_480_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        N_342_reto);
    
    \APB3_RDATA_1_am[4]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => N_1776, B => APB3_RDATA_1_sn_N_33_mux, C => 
        N_1757, Y => \APB3_RDATA_1_am[4]_net_1\);
    
    \mac_4_byte_4_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_4_reg[2]_net_1\);
    
    \APB3_RDATA_1_19_0_wmux_0[5]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_19_0_0_y0[5]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \mac_2_byte_5_reg[5]_net_1\, D => 
        \mac_4_byte_1_reg[5]_net_1\, FCI => 
        \APB3_RDATA_1_19_0_0_co0[5]\, S => OPEN, Y => N_1701, FCO
         => OPEN);
    
    \APB3_RDATA[5]\ : SLE
      port map(D => \APB3_RDATA_1[5]\, CLK => 
        \APB3_RDATA_31_sqmuxa_i\, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => VCC_net_1, Q => 
        CoreAPB3_0_APBmslave0_PRDATA(5));
    
    \REG_WRITE_PROC.un13_mac_2_byte_2_reg_en_0_a2_0_a2\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_420, B => \mac_2_byte_2_reg_en\, Y => 
        un13_mac_2_byte_2_reg_en);
    
    \mac_4_byte_3_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_3_reg[5]_net_1\);
    
    \APB3_RDATA_1_ns[5]\ : CFG4
      generic map(INIT => x"22FC")

      port map(A => \APB3_RDATA_1_bm[5]_net_1\, B => 
        APB3_RDATA_1_sn_N_33_mux, C => 
        \APB3_RDATA_1_29_d_ns[5]_net_1\, D => 
        \APB3_RDATA_1_ns_1[5]_net_1\, Y => \APB3_RDATA_1[5]\);
    
    \APB3_RDATA_1_bm_1[4]\ : CFG3
      generic map(INIT => x"1B")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => N_1578, 
        C => N_1660, Y => \APB3_RDATA_1_bm_1[4]_net_1\);
    
    \APB3_RDATA_1_19_0_0_wmux[1]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \i_int_mask_reg[1]_net_1\, D => \consumer_type2_reg[9]\, 
        FCI => VCC_net_1, S => OPEN, Y => 
        \APB3_RDATA_1_19_0_0_y0[1]\, FCO => 
        \APB3_RDATA_1_19_0_0_co0[1]\);
    
    \APB3_RDATA_1_24[6]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_1686, B => CoreAPB3_0_APBmslave0_PADDR(3), 
        C => N_1702, Y => N_1743);
    
    \APB3_RDATA_1_22_ns[0]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        \APB3_RDATA_1_22_am[0]_net_1\, C => 
        \APB3_RDATA_1_22_bm[0]_net_1\, Y => N_1720);
    
    \WRITE_REGISTER_ENABLE_PROC.un57_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => APB3_RDATA_1_sn_N_18, B => N_199, C => 
        CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => N_352);
    
    \WRITE_REGISTER_ENABLE_PROC.un13_apb3_addr_0_a2_2\ : CFG4
      generic map(INIT => x"0001")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CoreAPB3_0_APBmslave0_PADDR(7), C => 
        CoreAPB3_0_APBmslave0_PADDR(1), D => 
        CoreAPB3_0_APBmslave0_PADDR(0), Y => N_200);
    
    \REG_WRITE_PROC.un13_mac_4_byte_1_reg_en_0_a2_0_a2\ : CFG4
      generic map(INIT => x"0010")

      port map(A => \mac_3_byte_3_reg_en\, B => 
        \mac_3_byte_4_reg_en\, C => 
        un13_mac_4_byte_1_reg_en_0_a2_0_a2_1, D => N_141, Y => 
        un13_mac_4_byte_1_reg_en);
    
    \mac_4_byte_5_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_5_reg[5]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_2_byte_4_reg_en_0_a2_1_a2\ : CFG4
      generic map(INIT => x"0200")

      port map(A => \mac_2_byte_4_reg_en\, B => 
        \mac_2_byte_3_reg_en\, C => \mac_2_byte_2_reg_en\, D => 
        N_420, Y => un13_mac_2_byte_4_reg_en);
    
    \APB3_RDATA_1_21_0_wmux_0[2]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_21_0_0_y0[2]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \consumer_type1_reg[2]\, D => \consumer_type2_reg[2]\, 
        FCI => \APB3_RDATA_1_21_0_0_co0[2]\, S => OPEN, Y => 
        N_1714, FCO => OPEN);
    
    \APB3_RDATA_1_19_0_wmux_0[3]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_19_0_0_y0[3]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \mac_2_byte_5_reg[3]_net_1\, D => 
        \mac_4_byte_1_reg[3]_net_1\, FCI => 
        \APB3_RDATA_1_19_0_0_co0[3]\, S => OPEN, Y => N_1699, FCO
         => OPEN);
    
    \APB3_RDATA_1_19_0_wmux_0[2]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_19_0_0_y0[2]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \mac_2_byte_5_reg[2]_net_1\, D => 
        \mac_4_byte_1_reg[2]_net_1\, FCI => 
        \APB3_RDATA_1_19_0_0_co0[2]\, S => OPEN, Y => N_1698, FCO
         => OPEN);
    
    \APB3_RDATA_1_19_0_wmux_0[4]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_19_0_0_y0[4]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \mac_2_byte_5_reg[4]_net_1\, D => 
        \mac_4_byte_1_reg[4]_net_1\, FCI => 
        \APB3_RDATA_1_19_0_0_co0[4]\, S => OPEN, Y => N_1700, FCO
         => OPEN);
    
    \scratch_pad_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \write_scratch_reg_en\, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \scratch_pad_reg[3]_net_1\);
    
    \APB3_RDATA_1[3]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => \APB3_RDATA_1_d_ns[3]_net_1\, B => N_1765, C
         => \APB3_RDATA_1_s[7]_net_1\, Y => 
        \APB3_RDATA_1[3]_net_1\);
    
    \APB3_RDATA_1_bm[4]\ : CFG3
      generic map(INIT => x"72")

      port map(A => APB3_RDATA_1_sn_N_31_mux, B => 
        \APB3_RDATA_1_bm_1[4]_net_1\, C => N_1733, Y => 
        \APB3_RDATA_1_bm[4]_net_1\);
    
    mac_1_byte_2_reg_en_ret_4 : SLE
      port map(D => \mac_1_byte_2_reg_en\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        N_480_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        mac_1_byte_2_reg_en_reto);
    
    APB3_RDATA_31_sqmuxa_i_1 : CFG4
      generic map(INIT => x"0007")

      port map(A => \APB3_RDATA_31_sqmuxa_1_a3_0_2\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        CoreAPB3_0_APBmslave0_PADDR(1), D => 
        CoreAPB3_0_APBmslave0_PADDR(0), Y => 
        \APB3_RDATA_31_sqmuxa_i_1\);
    
    \mac_1_byte_5_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_5_reg[7]_net_1\);
    
    \APB3_RDATA_1_19_0_wmux_0[6]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_19_0_0_y0[6]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \mac_2_byte_5_reg[6]_net_1\, D => 
        \mac_4_byte_1_reg[6]_net_1\, FCI => 
        \APB3_RDATA_1_19_0_0_co0[6]\, S => OPEN, Y => N_1702, FCO
         => OPEN);
    
    \WRITE_REGISTER_ENABLE_PROC.un53_apb3_addr_0_a2_1\ : CFG4
      generic map(INIT => x"0002")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CoreAPB3_0_APBmslave0_PADDR(7), C => 
        CoreAPB3_0_APBmslave0_PADDR(1), D => 
        CoreAPB3_0_APBmslave0_PADDR(0), Y => N_199);
    
    \mac_2_byte_1_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_1_reg[4]_net_1\);
    
    \mac_1_byte_5_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_5_reg[4]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_2_byte_5_reg_en_0_a2_1_o2\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \mac_2_byte_4_reg_en\, B => 
        \mac_2_byte_3_reg_en\, C => \mac_2_byte_2_reg_en\, Y => 
        N_129);
    
    \APB3_RDATA_1_17_0_0_wmux[6]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => \rx_FIFO_rst_reg\, D
         => \mac_2_byte_3_reg[6]_net_1\, FCI => VCC_net_1, S => 
        OPEN, Y => \APB3_RDATA_1_17_0_0_y0[6]\, FCO => 
        \APB3_RDATA_1_17_0_0_co0[6]\);
    
    \mac_3_byte_2_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_2_reg[7]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un105_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => N_201, B => un105_apb3_addr_0_a2_0_1, C => 
        CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => N_364);
    
    \REG_WRITE_PROC.un12_mac_2_byte_1_reg_en_16_1\ : CFG4
      generic map(INIT => x"FFCA")

      port map(A => \mac_1_byte_4_reg_en\, B => 
        mac_4_byte_6_reg_en_1, C => N_344, D => N_11, Y => 
        un12_mac_2_byte_1_reg_en_16_1);
    
    \APB3_RDATA_1_18_0_wmux_0[7]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_18_0_0_y0[7]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_5_reg[7]_net_1\, D => 
        \mac_4_byte_6_reg[7]_net_1\, FCI => 
        \APB3_RDATA_1_18_0_0_co0[7]\, S => OPEN, Y => N_123, FCO
         => OPEN);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \mac_4_byte_1_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_1_reg[1]_net_1\);
    
    \APB3_RDATA_1_17_0_wmux_0[0]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_17_0_0_y0[0]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \consumer_type1_reg[8]\, D => \mac_3_byte_5_reg[0]_net_1\, 
        FCI => \APB3_RDATA_1_17_0_0_co0[0]\, S => OPEN, Y => 
        N_1680, FCO => OPEN);
    
    mac_1_byte_6_reg_en_0 : CFG4
      generic map(INIT => x"ACCC")

      port map(A => mac_4_byte_6_reg_en_1, B => 
        \mac_1_byte_6_reg_en\, C => N_213, D => N_201, Y => N_10);
    
    control_reg_en_ret_0 : SLE
      port map(D => N_803, CLK => m2s010_som_sb_0_CCC_71MHz, EN
         => VCC_net_1, ALn => N_480_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        N_812);
    
    \control_reg_RNO_0[5]\ : CFG4
      generic map(INIT => x"0CAA")

      port map(A => TX_PreAmble, B => \control_reg_en\, C => 
        \write_scratch_reg_en\, D => N_160, Y => 
        un1_control_reg_en_2_i_0);
    
    \APB3_RDATA[7]\ : SLE
      port map(D => \APB3_RDATA_1[7]_net_1\, CLK => 
        \APB3_RDATA_31_sqmuxa_i\, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => VCC_net_1, Q => 
        CoreAPB3_0_APBmslave0_PRDATA(7));
    
    \mac_4_byte_5_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_5_reg[1]_net_1\);
    
    \APB3_RDATA_1_18_0_0_wmux[5]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_3_reg[5]_net_1\, D => 
        \mac_4_byte_4_reg[5]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_18_0_0_y0[5]\, FCO => 
        \APB3_RDATA_1_18_0_0_co0[5]\);
    
    \mac_2_byte_6_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_6_reg[1]_net_1\);
    
    \mac_2_byte_1_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type4_reg[8]\);
    
    \WRITE_REGISTER_ENABLE_PROC.un61_apb3_addr_0_a2_0\ : CFG2
      generic map(INIT => x"2")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_212);
    
    \mac_3_byte_3_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_3_reg[7]_net_1\);
    
    \mac_1_byte_6_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type3_reg[6]\);
    
    \APB3_RDATA_1_25_0_0_wmux[5]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_1_byte_5_reg[5]_net_1\, D => 
        \mac_2_byte_1_reg[5]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_25_0_0_y0[5]\, FCO => 
        \APB3_RDATA_1_25_0_0_co0[5]\);
    
    \APB3_RDATA_1_15[1]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \int_reg[1]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_2_reg[1]_net_1\, Y => N_1665);
    
    \mac_2_byte_6_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_6_reg[7]_net_1\);
    
    \mac_3_byte_3_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_3_reg[1]_net_1\);
    
    \REG_WRITE_PROC.un12_mac_1_byte_2_reg_en_20\ : CFG4
      generic map(INIT => x"FAFC")

      port map(A => mac_4_byte_6_reg_en_1_reto, B => 
        mac_1_byte_2_reg_en_reto, C => N_802, D => N_342_reto, Y
         => N_801);
    
    mac_3_byte_6_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_358, ALn => N_480_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_3_byte_6_reg_en\);
    
    \WRITE_REGISTER_ENABLE_PROC.un9_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"0800")

      port map(A => APB3_RDATA_1_sn_N_18, B => N_200, C => 
        CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => N_339);
    
    \APB3_RDATA_1_29_d_ns[5]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \APB3_RDATA_1_29_d_bm[5]_net_1\, B => 
        \APB3_RDATA_1_29_d_am[5]_net_1\, C => 
        APB3_RDATA_1_sn_N_32_mux, Y => 
        \APB3_RDATA_1_29_d_ns[5]_net_1\);
    
    \APB3_RDATA_1_d[6]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => APB3_RDATA_1_sn_N_33_mux, B => 
        \APB3_RDATA_1_d_RNO[6]_net_1\, C => N_1778, Y => 
        \APB3_RDATA_1_d[6]_net_1\);
    
    \mac_1_byte_4_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type2_reg[2]\);
    
    APB3_RDATA_1_sn_m19_4_1_wmux_0 : ARI1
      generic map(INIT => x"0F588")

      port map(A => APB3_RDATA_1_sn_m19_4_1_0_y0, B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \APB3_RDATA_1_sn_m19_2\, D => APB3_RDATA_1_sn_N_18, FCI
         => APB3_RDATA_1_sn_m19_4_1_0_co0, S => OPEN, Y => 
        APB3_RDATA_1_sn_i6_mux, FCO => OPEN);
    
    \mac_2_byte_2_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type4_reg[5]\);
    
    \APB3_RDATA_1_15[2]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \int_reg[2]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_2_reg[2]_net_1\, Y => N_1666);
    
    \mac_4_byte_4_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_4_reg[7]_net_1\);
    
    \mac_1_byte_3_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_3_reg[5]_net_1\);
    
    \mac_4_byte_4_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_4_reg[6]_net_1\);
    
    \mac_4_byte_3_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_3_reg[6]_net_1\);
    
    \APB3_RDATA_1_29_s[6]\ : CFG3
      generic map(INIT => x"10")

      port map(A => APB3_RDATA_1_sn_i6_mux, B => \N_455_i\, C => 
        APB3_RDATA_1_sn_m8_out, Y => \APB3_RDATA_1_29_s[6]_net_1\);
    
    \APB3_RDATA_1_22_bm[1]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => RX_FIFO_DOUT(1), B => RX_FIFO_Full, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => 
        \APB3_RDATA_1_22_bm[1]_net_1\);
    
    \mac_2_byte_1_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_1_reg[6]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_4_byte_1_reg_en_0_a2_0_o2\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \mac_3_byte_4_reg_en\, B => 
        \mac_3_byte_3_reg_en\, C => N_141, Y => N_146);
    
    \REG_WRITE_PROC.un12_mac_2_byte_1_reg_en_16_2\ : CFG4
      generic map(INIT => x"FFCA")

      port map(A => \mac_1_byte_5_reg_en\, B => 
        mac_4_byte_6_reg_en_1, C => N_345, D => N_10, Y => 
        un12_mac_2_byte_1_reg_en_16_2);
    
    \i_int_mask_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_int_mask_reg_en_i_i_a2, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \i_int_mask_reg[7]_net_1\);
    
    \APB3_RDATA_1_3[3]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \consumer_type4_reg[3]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_4_reg[3]_net_1\, Y => N_1567);
    
    \mac_1_byte_5_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_5_reg[5]_net_1\);
    
    \RX_packet_depth_cry[0]\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \RX_packet_depth[0]_net_1\, B => 
        rx_packet_complt, C => GND_net_1, D => GND_net_1, FCI => 
        RX_packet_depth_s_914_FCO, S => \RX_packet_depth_s[0]\, Y
         => OPEN, FCO => \RX_packet_depth_cry[0]_net_1\);
    
    \mac_4_byte_4_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_4_reg[3]_net_1\);
    
    \APB3_RDATA_1_18_0_0_wmux[2]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_3_reg[2]_net_1\, D => 
        \mac_4_byte_4_reg[2]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_18_0_0_y0[2]\, FCO => 
        \APB3_RDATA_1_18_0_0_co0[2]\);
    
    \mac_4_byte_3_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_3_reg[4]_net_1\);
    
    \mac_4_byte_2_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_2_reg[3]_net_1\);
    
    \APB3_RDATA_1_19_0_0_wmux[6]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \i_int_mask_reg[6]_net_1\, D => 
        \mac_1_byte_3_reg[6]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_19_0_0_y0[6]\, FCO => 
        \APB3_RDATA_1_19_0_0_co0[6]\);
    
    \APB3_RDATA_1_17_0_wmux_0[1]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_17_0_0_y0[1]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \consumer_type1_reg[9]\, D => \mac_3_byte_5_reg[1]_net_1\, 
        FCI => \APB3_RDATA_1_17_0_0_co0[1]\, S => OPEN, Y => 
        N_1681, FCO => OPEN);
    
    APB3_RDATA_1_sn_m13 : CFG2
      generic map(INIT => x"4")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => APB3_RDATA_1_sn_N_14);
    
    \mac_2_byte_6_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_6_reg[4]_net_1\);
    
    \APB3_RDATA_1_1_1[0]\ : CFG4
      generic map(INIT => x"535F")

      port map(A => N_1753, B => N_1720, C => 
        APB3_RDATA_1_sn_N_32_mux, D => APB3_RDATA_1_sn_N_31_mux, 
        Y => \APB3_RDATA_1_1_0[0]_net_1\);
    
    \APB3_RDATA_1_28[2]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => N_1739, B => APB3_RDATA_1_sn_N_14, C => 
        N_1747, Y => N_1774);
    
    \REG_WRITE_PROC.un13_mac_2_byte_3_reg_en_0_a2_0_a2\ : CFG3
      generic map(INIT => x"20")

      port map(A => \mac_2_byte_3_reg_en\, B => 
        \mac_2_byte_2_reg_en\, C => N_420, Y => 
        un13_mac_2_byte_3_reg_en);
    
    mac_2_byte_4_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_350, ALn => N_480_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_2_byte_4_reg_en\);
    
    \APB3_RDATA_1_18_0_wmux_0[5]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_18_0_0_y0[5]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_5_reg[5]_net_1\, D => 
        \mac_4_byte_6_reg[5]_net_1\, FCI => 
        \APB3_RDATA_1_18_0_0_co0[5]\, S => OPEN, Y => N_121, FCO
         => OPEN);
    
    \APB3_RDATA_1_22_1_0[7]\ : CFG3
      generic map(INIT => x"47")

      port map(A => \consumer_type3_reg[7]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \scratch_pad_reg[7]_net_1\, Y => 
        \APB3_RDATA_1_22_1_0[7]_net_1\);
    
    \mac_4_byte_3_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_3_reg[3]_net_1\);
    
    \mac_4_byte_2_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_2_reg[4]_net_1\);
    
    \APB3_RDATA_1[0]\ : CFG4
      generic map(INIT => x"0C5D")

      port map(A => APB3_RDATA_1_sn_N_33_mux, B => 
        \APB3_RDATA_1_d_0[0]_net_1\, C => 
        \APB3_RDATA_1_1[0]_net_1\, D => 
        \APB3_RDATA_1_1_0[0]_net_1\, Y => \APB3_RDATA_1[0]_net_1\);
    
    APB3_RDATA_1_sn_m24 : CFG4
      generic map(INIT => x"DD50")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        APB3_RDATA_1_sn_N_23, C => CoreAPB3_0_APBmslave0_PADDR(4), 
        D => CoreAPB3_0_APBmslave0_PADDR(6), Y => 
        APB3_RDATA_1_sn_N_25);
    
    \REG_WRITE_PROC.un13_mac_2_byte_1_reg_en_0_a2_2_a2\ : CFG3
      generic map(INIT => x"80")

      port map(A => N_414, B => \mac_2_byte_1_reg_en\, C => N_413, 
        Y => un13_mac_2_byte_1_reg_en);
    
    \mac_1_byte_1_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type1_reg[9]\);
    
    \mac_1_byte_5_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type3_reg[9]\);
    
    \APB3_RDATA_1_21_0_0_wmux[7]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_2_byte_4_reg[7]_net_1\, D => 
        \mac_2_byte_6_reg[7]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_21_0_0_y0[7]\, FCO => 
        \APB3_RDATA_1_21_0_0_co0[7]\);
    
    \mac_2_byte_6_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_6_reg[2]_net_1\);
    
    \APB3_RDATA_1_25_0_wmux_0[5]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_25_0_0_y0[5]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_1_reg[5]_net_1\, D => 
        \mac_3_byte_3_reg[5]_net_1\, FCI => 
        \APB3_RDATA_1_25_0_0_co0[5]\, S => OPEN, Y => 
        \APB3_RDATA_1_25_0_wmux_0_Y[5]\, FCO => OPEN);
    
    APB3_RDATA_1_sn_m19_4_1_0_wmux : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \APB3_RDATA_1_sn_m19_0\, D => 
        CoreAPB3_0_APBmslave0_PADDR(7), FCI => VCC_net_1, S => 
        OPEN, Y => APB3_RDATA_1_sn_m19_4_1_0_y0, FCO => 
        APB3_RDATA_1_sn_m19_4_1_0_co0);
    
    \scratch_pad_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \write_scratch_reg_en\, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \scratch_pad_reg[5]_net_1\);
    
    APB3_RDATA_1_sn_m22 : CFG3
      generic map(INIT => x"2E")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => APB3_RDATA_1_sn_N_23);
    
    \APB3_RDATA_1_18_0_wmux_0[3]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_18_0_0_y0[3]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_5_reg[3]_net_1\, D => 
        \mac_4_byte_6_reg[3]_net_1\, FCI => 
        \APB3_RDATA_1_18_0_0_co0[3]\, S => OPEN, Y => N_119, FCO
         => OPEN);
    
    \APB3_RDATA_1_18_0_wmux_0[2]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_18_0_0_y0[2]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_5_reg[2]_net_1\, D => 
        \mac_4_byte_6_reg[2]_net_1\, FCI => 
        \APB3_RDATA_1_18_0_0_co0[2]\, S => OPEN, Y => N_118, FCO
         => OPEN);
    
    \APB3_RDATA_1_18_0_wmux_0[4]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_18_0_0_y0[4]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_5_reg[4]_net_1\, D => 
        \mac_4_byte_6_reg[4]_net_1\, FCI => 
        \APB3_RDATA_1_18_0_0_co0[4]\, S => OPEN, Y => N_120, FCO
         => OPEN);
    
    \mac_4_byte_2_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_2_reg[2]_net_1\);
    
    \mac_3_byte_5_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_5_reg[0]_net_1\);
    
    \APB3_RDATA_1_d_bm_RNO[3]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \APB3_RDATA_1_25_0_wmux_0_Y[3]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \APB3_RDATA_1_25_3[3]_net_1\, Y => N_1748);
    
    \mac_4_byte_3_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_3_reg[2]_net_1\);
    
    \APB3_RDATA_1_21_0_wmux_0[3]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_21_0_0_y0[3]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \consumer_type1_reg[3]\, D => \consumer_type2_reg[3]\, 
        FCI => \APB3_RDATA_1_21_0_0_co0[3]\, S => OPEN, Y => 
        N_1715, FCO => OPEN);
    
    APB3_RDATA_1_sn_m9 : CFG3
      generic map(INIT => x"47")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => APB3_RDATA_1_sn_N_10);
    
    \APB3_RDATA_1_18_0_wmux_0[6]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_18_0_0_y0[6]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_5_reg[6]_net_1\, D => 
        \mac_4_byte_6_reg[6]_net_1\, FCI => 
        \APB3_RDATA_1_18_0_0_co0[6]\, S => OPEN, Y => N_122, FCO
         => OPEN);
    
    \mac_1_byte_4_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type2_reg[7]\);
    
    \mac_1_byte_4_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type2_reg[6]\);
    
    \REG_WRITE_PROC.un13_int_mask_reg_en_i_i_a2\ : CFG2
      generic map(INIT => x"2")

      port map(A => \int_mask_reg_en\, B => N_813, Y => 
        un13_int_mask_reg_en_i_i_a2);
    
    \mac_2_byte_2_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type4_reg[6]\);
    
    \mac_1_byte_3_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_3_reg[6]_net_1\);
    
    \mac_2_byte_2_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type4_reg[1]\);
    
    mac_1_byte_6_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_346, ALn => N_480_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_1_byte_6_reg_en\);
    
    \APB3_RDATA_1_25_3[0]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_558, B => CoreAPB3_0_APBmslave0_PADDR(3), C
         => N_1564, Y => \APB3_RDATA_1_25_3[0]_net_1\);
    
    \APB3_RDATA_1_ns[4]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \APB3_RDATA_1_s[7]_net_1\, B => 
        \APB3_RDATA_1_am[4]_net_1\, C => 
        \APB3_RDATA_1_bm[4]_net_1\, Y => \APB3_RDATA_1[4]\);
    
    \APB3_RDATA_1_18_0_0_wmux[7]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_3_reg[7]_net_1\, D => 
        \mac_4_byte_4_reg[7]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_18_0_0_y0[7]\, FCO => 
        \APB3_RDATA_1_18_0_0_co0[7]\);
    
    \N_480_i\ : CFG4
      generic map(INIT => x"0080")

      port map(A => CoreAPB3_0_APBmslave0_PWRITE, B => 
        CoreAPB3_0_APBmslave0_PSELx, C => 
        CoreAPB3_0_APBmslave0_PENABLE, D => long_reset, Y => 
        N_480_i);
    
    \RX_PACKET_DEPTH_STATUS_PROC.un1_RX_packet_depthlto7_4\ : 
        CFG4
      generic map(INIT => x"0001")

      port map(A => \RX_packet_depth[7]_net_1\, B => 
        \RX_packet_depth[6]_net_1\, C => 
        \RX_packet_depth[5]_net_1\, D => 
        \RX_packet_depth[4]_net_1\, Y => 
        un1_RX_packet_depthlto7_4);
    
    \mac_4_byte_5_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_5_reg[2]_net_1\);
    
    \APB3_RDATA_1_22_ns[1]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        \APB3_RDATA_1_22_am[1]_net_1\, C => 
        \APB3_RDATA_1_22_bm[1]_net_1\, Y => N_1721);
    
    \mac_2_byte_1_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_1_reg[3]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_2_byte_5_reg_en_0_a2_1_a2\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_420, B => \mac_2_byte_5_reg_en\, C => N_129, 
        Y => un13_mac_2_byte_5_reg_en);
    
    \APB3_RDATA_1_21_0_0_wmux[5]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_2_byte_4_reg[5]_net_1\, D => 
        \mac_2_byte_6_reg[5]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_21_0_0_y0[5]\, FCO => 
        \APB3_RDATA_1_21_0_0_co0[5]\);
    
    \APB3_RDATA_1_25_3[5]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_55, B => CoreAPB3_0_APBmslave0_PADDR(3), C
         => N_1569, Y => \APB3_RDATA_1_25_3[5]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un41_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_199, D => N_201, Y
         => N_348);
    
    \mac_1_byte_4_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type2_reg[3]\);
    
    \APB3_RDATA_1_24[3]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_1683, B => CoreAPB3_0_APBmslave0_PADDR(3), 
        C => N_1699, Y => N_1740);
    
    \mac_1_byte_3_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_3_reg[4]_net_1\);
    
    \mac_1_byte_2_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type1_reg[3]\);
    
    \APB3_RDATA_1_29_d_am[5]\ : CFG4
      generic map(INIT => x"2075")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => RX_FIFO_DOUT(5), D
         => \APB3_RDATA_1_29_d_am_1_0[5]_net_1\, Y => 
        \APB3_RDATA_1_29_d_am[5]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_1_byte_6_reg_en_0_a2_1_a2_0\ : CFG3
      generic map(INIT => x"01")

      port map(A => \mac_1_byte_5_reg_en\, B => 
        \mac_1_byte_4_reg_en\, C => \mac_1_byte_3_reg_en\, Y => 
        N_412);
    
    \APB3_RDATA_1_26[2]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_1714, B => N_118, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_1755);
    
    mac_2_byte_1_reg_en_ret_4 : SLE
      port map(D => un12_mac_2_byte_1_reg_en_16_2, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        N_480_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        un12_mac_2_byte_1_reg_en_16_2_reto);
    
    \APB3_RDATA_1_18_0_0_wmux[4]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_3_reg[4]_net_1\, D => 
        \mac_4_byte_4_reg[4]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_18_0_0_y0[4]\, FCO => 
        \APB3_RDATA_1_18_0_0_co0[4]\);
    
    \RX_packet_depth[5]\ : SLE
      port map(D => \RX_packet_depth_s[5]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_1528_i, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RX_packet_depth[5]_net_1\);
    
    \REG_WRITE_PROC.un12_mac_1_byte_1_reg_en_20\ : CFG4
      generic map(INIT => x"FCFA")

      port map(A => mac_1_byte_1_reg_en_reto, B => 
        mac_4_byte_6_reg_en_1_reto_0, C => N_803_reto, D => 
        N_341_reto, Y => N_802);
    
    \mac_3_byte_5_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_5_reg[7]_net_1\);
    
    mac_4_byte_4_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_362, ALn => N_480_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_4_byte_4_reg_en\);
    
    \mac_2_byte_6_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_6_reg[5]_net_1\);
    
    \APB3_RDATA_1_29_d_am_1_0[5]\ : CFG3
      generic map(INIT => x"47")

      port map(A => \consumer_type3_reg[5]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \scratch_pad_reg[5]_net_1\, Y => 
        \APB3_RDATA_1_29_d_am_1_0[5]_net_1\);
    
    \RX_packet_depth_cry[6]\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \RX_packet_depth[6]_net_1\, B => 
        rx_packet_complt, C => GND_net_1, D => GND_net_1, FCI => 
        \RX_packet_depth_cry[5]_net_1\, S => 
        \RX_packet_depth_s[6]\, Y => OPEN, FCO => 
        \RX_packet_depth_cry[6]_net_1\);
    
    \mac_1_byte_3_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_3_reg[3]_net_1\);
    
    \mac_1_byte_2_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type1_reg[4]\);
    
    \mac_3_byte_5_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_5_reg[4]_net_1\);
    
    \mac_2_byte_4_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_4_reg[4]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un5_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"0008")

      port map(A => APB3_RDATA_1_sn_N_18, B => N_200, C => 
        CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => N_337);
    
    \REG_WRITE_PROC.un13_mac_3_byte_4_reg_en_0_a2_1_o2\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \mac_3_byte_2_reg_en\, B => 
        \mac_3_byte_1_reg_en\, C => N_131, Y => N_141);
    
    \mac_2_byte_6_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_6_reg[0]_net_1\);
    
    \APB3_RDATA_1_27[3]\ : CFG4
      generic map(INIT => x"FFB1")

      port map(A => APB3_RDATA_1_sn_m8_out, B => \read_reg_en\, C
         => \APB3_RDATA_1_27_d_0_wmux_0_Y[3]\, D => \N_455_i\, Y
         => N_1765);
    
    \REG_WRITE_PROC.un13_mac_1_byte_4_reg_en_0_a2_0_a2\ : CFG3
      generic map(INIT => x"20")

      port map(A => \mac_1_byte_4_reg_en\, B => 
        \mac_1_byte_3_reg_en\, C => N_414, Y => 
        un13_mac_1_byte_4_reg_en);
    
    \APB3_RDATA_1_24[7]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_1687, B => CoreAPB3_0_APBmslave0_PADDR(3), 
        C => N_1703, Y => N_1744);
    
    \APB3_RDATA_1_15[7]\ : CFG4
      generic map(INIT => x"C5C0")

      port map(A => \i_int_mask_reg[7]_net_1\, B => 
        \mac_4_byte_2_reg[7]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(3), D => tx_packet_complt_int, 
        Y => N_1671);
    
    \mac_2_byte_1_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_1_reg[5]_net_1\);
    
    \scratch_pad_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \write_scratch_reg_en\, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \scratch_pad_reg[7]_net_1\);
    
    \APB3_RDATA_1_25_0_0_wmux[6]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_1_byte_5_reg[6]_net_1\, D => 
        \mac_2_byte_1_reg[6]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_25_0_0_y0[6]\, FCO => 
        \APB3_RDATA_1_25_0_0_co0[6]\);
    
    \mac_4_byte_1_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_1_reg[4]_net_1\);
    
    \APB3_RDATA_1_25_0_0_wmux[0]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \consumer_type3_reg[8]\, D => \consumer_type4_reg[8]\, 
        FCI => VCC_net_1, S => OPEN, Y => 
        \APB3_RDATA_1_25_0_0_y0[0]\, FCO => 
        \APB3_RDATA_1_25_0_0_co0[0]\);
    
    \mac_3_byte_6_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_6_reg[6]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_4_byte_2_reg_en_0_a2_3_o2_0\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \mac_4_byte_1_reg_en\, B => 
        \mac_3_byte_6_reg_en\, C => \mac_3_byte_5_reg_en\, Y => 
        un13_mac_4_byte_2_reg_en_0_a2_3_o2_0);
    
    \APB3_RDATA_1_18_0_0_wmux[1]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_3_reg[1]_net_1\, D => 
        \mac_4_byte_4_reg[1]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_18_0_0_y0[1]\, FCO => 
        \APB3_RDATA_1_18_0_0_co0[1]\);
    
    \APB3_RDATA_1_21_0_wmux_0[7]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_21_0_0_y0[7]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \consumer_type1_reg[7]\, D => \consumer_type2_reg[7]\, 
        FCI => \APB3_RDATA_1_21_0_0_co0[7]\, S => OPEN, Y => 
        N_1719, FCO => OPEN);
    
    \mac_2_byte_1_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_1_reg[2]_net_1\);
    
    \mac_1_byte_2_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type1_reg[2]\);
    
    \APB3_RDATA_1_25_0_wmux_0[4]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_25_0_0_y0[4]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_1_reg[4]_net_1\, D => 
        \mac_3_byte_3_reg[4]_net_1\, FCI => 
        \APB3_RDATA_1_25_0_0_co0[4]\, S => OPEN, Y => 
        \APB3_RDATA_1_25_0_wmux_0_Y[4]\, FCO => OPEN);
    
    \mac_1_byte_3_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_3_reg[2]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un101_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"0800")

      port map(A => N_201, B => un105_apb3_addr_0_a2_0_1, C => 
        CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => N_363);
    
    \APB3_RDATA_1_27_d_1[6]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        \APB3_RDATA_1_27_d_0[6]_net_1\, C => 
        \mac_4_byte_2_reg[6]_net_1\, Y => 
        \APB3_RDATA_1_27_d_1[6]_net_1\);
    
    \mac_4_byte_6_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_6_reg[1]_net_1\);
    
    \mac_4_byte_1_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_1_reg[0]_net_1\);
    
    \APB3_RDATA_1_23[1]\ : CFG3
      generic map(INIT => x"EF")

      port map(A => \N_455_i\, B => N_1665, C => 
        APB3_RDATA_1_sn_m8_out, Y => N_1730);
    
    \mac_3_byte_4_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_4_reg[2]_net_1\);
    
    \mac_2_byte_4_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_4_reg[1]_net_1\);
    
    \APB3_RDATA_1_17_0_0_wmux[3]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => \control_reg_3\, D
         => \mac_2_byte_3_reg[3]_net_1\, FCI => VCC_net_1, S => 
        OPEN, Y => \APB3_RDATA_1_17_0_0_y0[3]\, FCO => 
        \APB3_RDATA_1_17_0_0_co0[3]\);
    
    \mac_2_byte_4_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_4_reg[0]_net_1\);
    
    \APB3_RDATA_1_17_0_0_wmux[0]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => \control_reg_0\, D
         => \mac_2_byte_3_reg[0]_net_1\, FCI => VCC_net_1, S => 
        OPEN, Y => \APB3_RDATA_1_17_0_0_y0[0]\, FCO => 
        \APB3_RDATA_1_17_0_0_co0[0]\);
    
    \mac_4_byte_6_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_6_reg[7]_net_1\);
    
    \APB3_RDATA_1_27_d_0_0_wmux[3]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        APB3_RDATA_1_sn_N_31_mux, C => \int_reg[3]\, D => 
        \mac_4_byte_2_reg[3]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_27_d_0_0_y0[3]\, FCO => 
        \APB3_RDATA_1_27_d_0_0_co0[3]\);
    
    \RX_packet_depth[1]\ : SLE
      port map(D => \RX_packet_depth_s[1]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_1528_i, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RX_packet_depth[1]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_4_byte_6_reg_en_0_a2_4_o2_RNI16D31\ : 
        CFG4
      generic map(INIT => x"FFFE")

      port map(A => un1_control_reg_en_2_i_0_0_o2_0, B => N_146, 
        C => un13_mac_4_byte_2_reg_en_0_a2_3_o2_0, D => N_157, Y
         => N_160);
    
    \mac_3_byte_3_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_3_reg[5]_net_1\);
    
    \APB3_RDATA_1_d_bm[3]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => N_1740, B => APB3_RDATA_1_sn_N_14, C => 
        N_1748, Y => \APB3_RDATA_1_d_bm[3]_net_1\);
    
    \APB3_RDATA_1_28_RNO[6]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \APB3_RDATA_1_25_0_wmux_0_Y[6]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \APB3_RDATA_1_25_3[6]_net_1\, Y => N_1751);
    
    \APB3_RDATA_1_4[4]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \consumer_type3_reg[4]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \scratch_pad_reg[4]_net_1\, Y => N_1578);
    
    \REG_WRITE_PROC.un13_mac_2_byte_1_reg_en_0_a2_2_a2_0\ : CFG4
      generic map(INIT => x"0001")

      port map(A => \mac_1_byte_6_reg_en\, B => 
        \mac_1_byte_5_reg_en\, C => \mac_1_byte_4_reg_en\, D => 
        \mac_1_byte_3_reg_en\, Y => N_413);
    
    \mac_1_byte_5_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_5_reg[2]_net_1\);
    
    APB3_RDATA_1_sn_m19_2 : CFG4
      generic map(INIT => x"EE50")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        CoreAPB3_0_APBmslave0_PADDR(7), D => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => 
        \APB3_RDATA_1_sn_m19_2\);
    
    \APB3_RDATA_1_3[5]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \consumer_type4_reg[5]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_4_reg[5]_net_1\, Y => N_1569);
    
    mac_2_byte_1_reg_en_ret_8 : SLE
      port map(D => \mac_1_byte_1_reg_en\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        N_480_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        mac_1_byte_1_reg_en_reto);
    
    \mac_2_byte_4_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_4_reg[5]_net_1\);
    
    \mac_4_byte_2_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_2_reg[5]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_4_byte_3_reg_en_0_a2_4_a2\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \mac_1_byte_2_reg_en\, B => 
        \mac_1_byte_1_reg_en\, C => N_553, D => 
        un13_mac_4_byte_3_reg_en_0_a2_4_a2_2, Y => 
        un13_mac_4_byte_3_reg_en);
    
    \APB3_RDATA_1_3[7]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \consumer_type4_reg[7]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_4_reg[7]_net_1\, Y => N_1571);
    
    mac_2_byte_1_reg_en_ret_5 : SLE
      port map(D => N_341, CLK => m2s010_som_sb_0_CCC_71MHz, EN
         => VCC_net_1, ALn => N_480_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        N_341_reto);
    
    \mac_3_byte_5_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_5_reg[5]_net_1\);
    
    \APB3_RDATA_1_bm[1]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_1754, B => N_1721, C => 
        APB3_RDATA_1_sn_N_32_mux, Y => \APB3_RDATA_1_bm[1]_net_1\);
    
    \APB3_RDATA_1_27_d_3_1[6]\ : CFG3
      generic map(INIT => x"47")

      port map(A => \consumer_type3_reg[6]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \scratch_pad_reg[6]_net_1\, Y => 
        \APB3_RDATA_1_27_d_3_1[6]_net_1\);
    
    \mac_2_byte_6_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_6_reg[3]_net_1\);
    
    \mac_4_byte_1_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_1_reg[6]_net_1\);
    
    mac_2_byte_2_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_348, ALn => N_480_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_2_byte_2_reg_en\);
    
    \iAPB3_READY_RNIKLOT[1]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => CoreAPB3_0_APBmslave0_PREADYrs, B => 
        un5_apb3_rst_rs, C => long_reset_set, Y => 
        \CoreAPB3_0_APBmslave0_PREADY\);
    
    \REG_WRITE_PROC.un13_mac_4_byte_5_reg_en_0_a2_0_a2_0\ : CFG2
      generic map(INIT => x"4")

      port map(A => N_802, B => \mac_4_byte_5_reg_en\, Y => 
        un13_mac_4_byte_5_reg_en_0_a2_0_a2_0);
    
    \APB3_RDATA_1_3[0]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \consumer_type4_reg[0]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_4_reg[0]_net_1\, Y => N_1564);
    
    \APB3_RDATA[4]\ : SLE
      port map(D => \APB3_RDATA_1[4]\, CLK => 
        \APB3_RDATA_31_sqmuxa_i\, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => VCC_net_1, Q => 
        CoreAPB3_0_APBmslave0_PRDATA(4));
    
    \APB3_RDATA_1_14[2]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => RX_FIFO_DOUT(2), B => TX_FIFO_Empty, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_1658);
    
    mac_3_byte_4_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_356, ALn => N_480_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_3_byte_4_reg_en\);
    
    RX_packet_depth_s_914 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => rx_packet_complt, C => 
        GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => OPEN, Y
         => OPEN, FCO => RX_packet_depth_s_914_FCO);
    
    \APB3_RDATA_1_25_3[4]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_562, B => CoreAPB3_0_APBmslave0_PADDR(3), C
         => N_1568, Y => \APB3_RDATA_1_25_3[4]_net_1\);
    
    control_reg_en_ret : SLE
      port map(D => N_804, CLK => m2s010_som_sb_0_CCC_71MHz, EN
         => VCC_net_1, ALn => N_480_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        N_813);
    
    \APB3_RDATA_1_25_3[1]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_559, B => CoreAPB3_0_APBmslave0_PADDR(3), C
         => N_1565, Y => \APB3_RDATA_1_25_3[1]_net_1\);
    
    \iup_EOP\ : SLE
      port map(D => un116_apb3_addr, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => iup_EOP_net_1);
    
    \APB3_RDATA_1_23[2]\ : CFG3
      generic map(INIT => x"EF")

      port map(A => \N_455_i\, B => N_1666, C => 
        APB3_RDATA_1_sn_m8_out, Y => N_1731);
    
    \mac_4_byte_6_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_6_reg[4]_net_1\);
    
    \mac_3_byte_1_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_1_reg[1]_net_1\);
    
    \mac_3_byte_5_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_5_reg[1]_net_1\);
    
    \APB3_RDATA_1_24[5]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_1685, B => CoreAPB3_0_APBmslave0_PADDR(3), 
        C => N_1701, Y => N_1742);
    
    \mac_1_byte_1_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_1_reg[4]_net_1\);
    
    \mac_2_byte_1_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_1_reg[7]_net_1\);
    
    \APB3_RDATA_1_24[1]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_1681, B => CoreAPB3_0_APBmslave0_PADDR(3), 
        C => N_1697, Y => N_1738);
    
    \APB3_RDATA_1_19_0_0_wmux[3]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \i_int_mask_reg[3]_net_1\, D => 
        \mac_1_byte_3_reg[3]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_19_0_0_y0[3]\, FCO => 
        \APB3_RDATA_1_19_0_0_co0[3]\);
    
    \APB3_RDATA_1_19_0_0_wmux[0]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \i_int_mask_reg[0]_net_1\, D => \consumer_type2_reg[8]\, 
        FCI => VCC_net_1, S => OPEN, Y => 
        \APB3_RDATA_1_19_0_0_y0[0]\, FCO => 
        \APB3_RDATA_1_19_0_0_co0[0]\);
    
    \REG_WRITE_PROC.un12_control_reg_en_0\ : CFG4
      generic map(INIT => x"FFCA")

      port map(A => \write_scratch_reg_en\, B => 
        mac_4_byte_6_reg_en_1, C => N_335, D => N_3, Y => N_804);
    
    APB3_RDATA_31_sqmuxa_1_a3_0_2 : CFG4
      generic map(INIT => x"0001")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(7), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        CoreAPB3_0_APBmslave0_PADDR(4), D => 
        CoreAPB3_0_APBmslave0_PADDR(2), Y => 
        \APB3_RDATA_31_sqmuxa_1_a3_0_2\);
    
    mac_2_byte_5_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_351, ALn => N_480_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_2_byte_5_reg_en\);
    
    \WRITE_REGISTER_ENABLE_PROC.un49_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"0080")

      port map(A => APB3_RDATA_1_sn_N_18, B => N_199, C => 
        CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => N_350);
    
    \PROCESSOR_EOP_READ_PROC.un116_apb3_addr\ : CFG4
      generic map(INIT => x"8000")

      port map(A => N_336, B => RX_FIFO_DOUT(8), C => 
        \read_reg_en\, D => \CoreAPB3_0_APBmslave0_PREADY\, Y => 
        un116_apb3_addr);
    
    APB3_RDATA_1_sn_m17 : CFG2
      generic map(INIT => x"4")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => APB3_RDATA_1_sn_N_18);
    
    \APB3_RDATA_1_25_0_wmux_0[0]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_25_0_0_y0[0]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_1_reg[0]_net_1\, D => 
        \mac_3_byte_3_reg[0]_net_1\, FCI => 
        \APB3_RDATA_1_25_0_0_co0[0]\, S => OPEN, Y => 
        \APB3_RDATA_1_25_0_wmux_0_Y[0]\, FCO => OPEN);
    
    \APB3_RDATA_1_14[4]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => RX_FIFO_DOUT(4), B => 
        RX_packet_depth_status_net_1, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_1660);
    
    \APB3_RDATA_1_21_0_wmux_0[5]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_21_0_0_y0[5]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \consumer_type1_reg[5]\, D => \consumer_type2_reg[5]\, 
        FCI => \APB3_RDATA_1_21_0_0_co0[5]\, S => OPEN, Y => 
        N_1717, FCO => OPEN);
    
    \RX_packet_depth[7]\ : SLE
      port map(D => \RX_packet_depth_s[7]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_1528_i, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RX_packet_depth[7]_net_1\);
    
    \mac_2_byte_2_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type4_reg[0]\);
    
    \mac_1_byte_6_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type3_reg[1]\);
    
    \mac_1_byte_1_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type1_reg[8]\);
    
    \mac_4_byte_6_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_6_reg[2]_net_1\);
    
    \i_int_mask_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_int_mask_reg_en_i_i_a2, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \i_int_mask_reg[5]_net_1\);
    
    \APB3_RDATA_1_25_4_wmux_3[7]\ : ARI1
      generic map(INIT => x"0EC2C")

      port map(A => \APB3_RDATA_1_25_4_0_y3[7]\, B => 
        \APB3_RDATA_1_25_4_0_y1[7]\, C => 
        CoreAPB3_0_APBmslave0_PADDR(2), D => VCC_net_1, FCI => 
        \APB3_RDATA_1_25_4_co1_0[7]\, S => OPEN, Y => N_1752, FCO
         => OPEN);
    
    read_reg_en_RNI5GHE2 : CFG3
      generic map(INIT => x"40")

      port map(A => \N_455_i\, B => \read_reg_en\, C => 
        APB3_RDATA_1_sn_N_25, Y => APB3_RDATA_1_sn_N_33_mux);
    
    \APB3_RDATA_1_18_0_0_wmux[6]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_3_reg[6]_net_1\, D => 
        \mac_4_byte_4_reg[6]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_18_0_0_y0[6]\, FCO => 
        \APB3_RDATA_1_18_0_0_co0[6]\);
    
    \mac_1_byte_6_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type3_reg[7]\);
    
    \WRITE_REGISTER_ENABLE_PROC.un45_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"0008")

      port map(A => APB3_RDATA_1_sn_N_18, B => N_199, C => 
        CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => N_349);
    
    \APB3_RDATA_1_3[1]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \consumer_type4_reg[1]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_4_reg[1]_net_1\, Y => N_1565);
    
    \mac_3_byte_4_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_4_reg[7]_net_1\);
    
    \mac_3_byte_4_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_4_reg[6]_net_1\);
    
    \mac_3_byte_3_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_3_reg[6]_net_1\);
    
    \APB3_RDATA_1_19_0_wmux_0[0]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_19_0_0_y0[0]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \mac_2_byte_5_reg[0]_net_1\, D => 
        \mac_4_byte_1_reg[0]_net_1\, FCI => 
        \APB3_RDATA_1_19_0_0_co0[0]\, S => OPEN, Y => N_1696, FCO
         => OPEN);
    
    \APB3_RDATA_1_28_RNO[5]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \APB3_RDATA_1_25_0_wmux_0_Y[5]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \APB3_RDATA_1_25_3[5]_net_1\, Y => N_1750);
    
    \APB3_RDATA_1_21_0_0_wmux[6]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_2_byte_4_reg[6]_net_1\, D => 
        \mac_2_byte_6_reg[6]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_21_0_0_y0[6]\, FCO => 
        \APB3_RDATA_1_21_0_0_co0[6]\);
    
    \APB3_RDATA[1]\ : SLE
      port map(D => \APB3_RDATA_1[1]\, CLK => 
        \APB3_RDATA_31_sqmuxa_i\, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => VCC_net_1, Q => 
        CoreAPB3_0_APBmslave0_PRDATA(1));
    
    \REG_WRITE_PROC.un13_mac_3_byte_6_reg_en_0_a2_1_a2\ : CFG4
      generic map(INIT => x"0020")

      port map(A => \mac_3_byte_6_reg_en\, B => 
        \mac_3_byte_5_reg_en\, C => N_420, D => N_146, Y => 
        un13_mac_3_byte_6_reg_en);
    
    \APB3_RDATA_1_22_am[0]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \consumer_type3_reg[0]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \scratch_pad_reg[0]_net_1\, Y => 
        \APB3_RDATA_1_22_am[0]_net_1\);
    
    \i_int_mask_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_int_mask_reg_en_i_i_a2, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \i_int_mask_reg[2]_net_1\);
    
    \APB3_RDATA_1_4[3]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \consumer_type3_reg[3]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \scratch_pad_reg[3]_net_1\, Y => N_1577);
    
    \mac_2_byte_3_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_3_reg[0]_net_1\);
    
    \APB3_RDATA_1_25_0_wmux_0[1]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_25_0_0_y0[1]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_1_reg[1]_net_1\, D => 
        \mac_3_byte_3_reg[1]_net_1\, FCI => 
        \APB3_RDATA_1_25_0_0_co0[1]\, S => OPEN, Y => 
        \APB3_RDATA_1_25_0_wmux_0_Y[1]\, FCO => OPEN);
    
    \APB3_RDATA_1_21_0_0_wmux[0]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_2_byte_4_reg[0]_net_1\, D => 
        \mac_2_byte_6_reg[0]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_21_0_0_y0[0]\, FCO => 
        \APB3_RDATA_1_21_0_0_co0[0]\);
    
    \WRITE_REGISTER_ENABLE_PROC.un65_apb3_addr_0_a2_0\ : CFG3
      generic map(INIT => x"40")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => N_199, C
         => CoreAPB3_0_APBmslave0_PADDR(2), Y => N_213);
    
    \mac_1_byte_2_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type1_reg[5]\);
    
    \APB3_RDATA_1_25_4_wmux_0[7]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_25_4_0_y0[7]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_1_reg[7]_net_1\, D => 
        \mac_3_byte_3_reg[7]_net_1\, FCI => 
        \APB3_RDATA_1_25_4_0_co0[7]\, S => OPEN, Y => 
        \APB3_RDATA_1_25_4_0_y1[7]\, FCO => 
        \APB3_RDATA_1_25_4_0_co1[7]\);
    
    \READY_DELAY_PROC.un5_apb3_rst_0_a2\ : CFG3
      generic map(INIT => x"F8")

      port map(A => CoreAPB3_0_APBmslave0_PSELx, B => 
        CoreAPB3_0_APBmslave0_PENABLE, C => long_reset, Y => 
        un5_apb3_rst_i);
    
    \APB3_RDATA_1_1_0[0]\ : CFG3
      generic map(INIT => x"54")

      port map(A => APB3_RDATA_1_sn_N_33_mux, B => 
        APB3_RDATA_1_sn_N_31_mux, C => APB3_RDATA_1_sn_N_32_mux, 
        Y => \APB3_RDATA_1_1[0]_net_1\);
    
    \APB3_RDATA_1[7]\ : CFG3
      generic map(INIT => x"AB")

      port map(A => \APB3_RDATA_1_4\, B => 
        APB3_RDATA_1_sn_N_33_mux, C => \APB3_RDATA_1_1[7]_net_1\, 
        Y => \APB3_RDATA_1[7]_net_1\);
    
    \mac_3_byte_4_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_4_reg[3]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un33_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"4000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_199, D => N_201, Y
         => N_346);
    
    \mac_4_byte_2_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_2_reg[6]_net_1\);
    
    \mac_4_byte_2_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_2_reg[1]_net_1\);
    
    mac_4_byte_2_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_360, ALn => N_480_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_4_byte_2_reg_en\);
    
    \mac_3_byte_3_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_3_reg[4]_net_1\);
    
    \mac_3_byte_2_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_2_reg[3]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.mac_4_byte_6_reg_en_1\ : CFG2
      generic map(INIT => x"4")

      port map(A => \CoreAPB3_0_APBmslave0_PREADY\, B => 
        \iAPB3_READY[0]_net_1\, Y => mac_4_byte_6_reg_en_1);
    
    read_reg_en_RNIICDH5 : CFG3
      generic map(INIT => x"40")

      port map(A => \N_455_i\, B => \read_reg_en\, C => 
        APB3_RDATA_1_sn_i6_mux, Y => APB3_RDATA_1_sn_N_32_mux);
    
    \APB3_RDATA_1_15[4]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \int_reg[4]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_2_reg[4]_net_1\, Y => N_1668);
    
    \mac_1_byte_1_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_1_reg[6]_net_1\);
    
    \RX_packet_depth[4]\ : SLE
      port map(D => \RX_packet_depth_s[4]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_1528_i, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RX_packet_depth[4]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un13_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"1000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_200, D => N_202, Y
         => N_341);
    
    \mac_4_byte_1_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_1_reg[3]_net_1\);
    
    \APB3_RDATA_1_25_0_0_wmux[1]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \consumer_type3_reg[9]\, D => \consumer_type4_reg[9]\, 
        FCI => VCC_net_1, S => OPEN, Y => 
        \APB3_RDATA_1_25_0_0_y0[1]\, FCO => 
        \APB3_RDATA_1_25_0_0_co0[1]\);
    
    \iAPB3_READY[1]\ : SLE
      port map(D => \iAPB3_READY[0]_net_1\, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        un5_apb3_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, SD
         => GND_net_1, LAT => GND_net_1, Q => 
        CoreAPB3_0_APBmslave0_PREADYrs);
    
    \mac_2_byte_5_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_5_reg[3]_net_1\);
    
    \control_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => control_reg_22, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \rx_FIFO_rst_reg\);
    
    \REG_WRITE_PROC.un13_mac_3_byte_1_reg_en_0_a2_1_a2\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_420, B => \mac_3_byte_1_reg_en\, C => N_131, 
        Y => un13_mac_3_byte_1_reg_en);
    
    \REG_WRITE_PROC.un13_mac_4_byte_6_reg_en_0_a2_4_a2\ : CFG4
      generic map(INIT => x"0040")

      port map(A => N_801, B => N_553, C => \mac_4_byte_6_reg_en\, 
        D => N_157, Y => un13_mac_4_byte_6_reg_en);
    
    \REG_WRITE_PROC.un13_mac_4_byte_4_reg_en_0_a2_0_a2_1\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \mac_4_byte_3_reg_en\, B => 
        \mac_4_byte_2_reg_en\, C => N_812, D => 
        \mac_4_byte_4_reg_en\, Y => 
        un13_mac_4_byte_4_reg_en_0_a2_0_a2_1);
    
    \APB3_RDATA_1_ns[1]\ : CFG4
      generic map(INIT => x"CCE2")

      port map(A => \APB3_RDATA_1_bm[1]_net_1\, B => 
        \APB3_RDATA_1_ns_1[1]_net_1\, C => N_1730, D => 
        APB3_RDATA_1_sn_N_33_mux, Y => \APB3_RDATA_1[1]\);
    
    \mac_3_byte_3_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_3_reg[3]_net_1\);
    
    \mac_3_byte_2_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_2_reg[4]_net_1\);
    
    iRX_FIFO_rd_en_RNO : CFG1
      generic map(INIT => "01")

      port map(A => \iAPB3_READY[0]_net_1\, Y => 
        \iAPB3_READY_i[0]\);
    
    \mac_1_byte_6_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type3_reg[4]\);
    
    \APB3_RDATA_1_25_0_wmux_0[6]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_25_0_0_y0[6]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_1_reg[6]_net_1\, D => 
        \mac_3_byte_3_reg[6]_net_1\, FCI => 
        \APB3_RDATA_1_25_0_0_co0[6]\, S => OPEN, Y => 
        \APB3_RDATA_1_25_0_wmux_0_Y[6]\, FCO => OPEN);
    
    \APB3_RDATA_1_am_1_RNO[1]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \APB3_RDATA_1_25_0_wmux_0_Y[1]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \APB3_RDATA_1_25_3[1]_net_1\, Y => N_1746);
    
    \mac_2_byte_5_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_5_reg[6]_net_1\);
    
    \RX_packet_depth_cry[2]\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \RX_packet_depth[2]_net_1\, B => 
        rx_packet_complt, C => GND_net_1, D => GND_net_1, FCI => 
        \RX_packet_depth_cry[1]_net_1\, S => 
        \RX_packet_depth_s[2]\, Y => OPEN, FCO => 
        \RX_packet_depth_cry[2]_net_1\);
    
    \APB3_RDATA_1_ns[2]\ : CFG3
      generic map(INIT => x"E4")

      port map(A => \APB3_RDATA_1_s[7]_net_1\, B => 
        \APB3_RDATA_1_am[2]_net_1\, C => 
        \APB3_RDATA_1_bm[2]_net_1\, Y => \APB3_RDATA_1[2]\);
    
    \RX_packet_depth[0]\ : SLE
      port map(D => \RX_packet_depth_s[0]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_1528_i, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RX_packet_depth[0]_net_1\);
    
    \mac_4_byte_6_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_6_reg[5]_net_1\);
    
    mac_1_byte_4_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_344, ALn => N_480_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_1_byte_4_reg_en\);
    
    read_reg_en_RNI3OAV1 : CFG4
      generic map(INIT => x"0800")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \read_reg_en\, C => \N_455_i\, D => APB3_RDATA_1_sn_N_10, 
        Y => APB3_RDATA_1_sn_N_31_mux);
    
    mac_4_byte_5_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_363, ALn => N_480_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_4_byte_5_reg_en\);
    
    \APB3_RDATA_1_19_0_wmux_0[1]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_19_0_0_y0[1]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \mac_2_byte_5_reg[1]_net_1\, D => 
        \mac_4_byte_1_reg[1]_net_1\, FCI => 
        \APB3_RDATA_1_19_0_0_co0[1]\, S => OPEN, Y => N_1697, FCO
         => OPEN);
    
    \mac_4_byte_4_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_4_reg[4]_net_1\);
    
    \mac_4_byte_6_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_6_reg[0]_net_1\);
    
    mac_1_byte_2_reg_en_ret_3 : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        N_480_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        mac_4_byte_6_reg_en_1_reto);
    
    \APB3_RDATA_1_25_4_wmux_2[7]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_25_4_y0_0[7]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => N_57, D => N_1571, 
        FCI => \APB3_RDATA_1_25_4_co0_0[7]\, S => OPEN, Y => 
        \APB3_RDATA_1_25_4_0_y3[7]\, FCO => 
        \APB3_RDATA_1_25_4_co1_0[7]\);
    
    \mac_3_byte_2_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_2_reg[2]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_3_byte_2_reg_en_0_a2_1_a2\ : CFG4
      generic map(INIT => x"0040")

      port map(A => \mac_3_byte_1_reg_en\, B => 
        \mac_3_byte_2_reg_en\, C => N_420, D => N_131, Y => 
        un13_mac_3_byte_2_reg_en);
    
    \mac_4_byte_1_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_1_reg[5]_net_1\);
    
    \mac_1_byte_6_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type3_reg[2]\);
    
    \mac_3_byte_3_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_3_reg[2]_net_1\);
    
    mac_2_byte_1_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_347, ALn => N_480_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_2_byte_1_reg_en\);
    
    \APB3_RDATA_1_27_d_0_wmux_0[3]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_27_d_0_0_y0[3]\, B => 
        APB3_RDATA_1_sn_N_31_mux, C => N_1577, D => N_1659, FCI
         => \APB3_RDATA_1_27_d_0_0_co0[3]\, S => OPEN, Y => 
        \APB3_RDATA_1_27_d_0_wmux_0_Y[3]\, FCO => OPEN);
    
    \WRITE_REGISTER_ENABLE_PROC.un61_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"1000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_199, D => N_212, Y
         => N_353);
    
    \APB3_RDATA_1_23[4]\ : CFG3
      generic map(INIT => x"EF")

      port map(A => \N_455_i\, B => N_1668, C => 
        APB3_RDATA_1_sn_m8_out, Y => N_1733);
    
    \APB3_RDATA_1_21_0_wmux_0[4]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_21_0_0_y0[4]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \consumer_type1_reg[4]\, D => \consumer_type2_reg[4]\, 
        FCI => \APB3_RDATA_1_21_0_0_co0[4]\, S => OPEN, Y => 
        N_1716, FCO => OPEN);
    
    \mac_4_byte_1_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_1_reg[2]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un81_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"4000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_199, D => N_202, Y
         => N_358);
    
    \mac_3_byte_5_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_5_reg[2]_net_1\);
    
    \mac_4_byte_4_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_4_reg[1]_net_1\);
    
    write_scratch_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_335, ALn => N_480_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \write_scratch_reg_en\);
    
    N_455_i : CFG4
      generic map(INIT => x"CC4C")

      port map(A => CoreAPB3_0_APBmslave0_PENABLE, B => 
        long_reset, C => CoreAPB3_0_APBmslave0_PSELx, D => 
        CoreAPB3_0_APBmslave0_PWRITE, Y => \N_455_i\);
    
    \mac_4_byte_4_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_4_reg[0]_net_1\);
    
    control_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_337, ALn => N_480_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \control_reg_en\);
    
    \mac_2_byte_2_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type4_reg[7]\);
    
    \mac_1_byte_2_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type1_reg[6]\);
    
    \mac_1_byte_2_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type1_reg[1]\);
    
    mac_2_byte_1_reg_en_0 : CFG3
      generic map(INIT => x"CA")

      port map(A => \mac_2_byte_1_reg_en\, B => 
        mac_4_byte_6_reg_en_1, C => N_347, Y => N_11);
    
    \REG_WRITE_PROC.un13_mac_1_byte_6_reg_en_0_a2_1_a2\ : CFG3
      generic map(INIT => x"80")

      port map(A => N_414, B => \mac_1_byte_6_reg_en\, C => N_412, 
        Y => un13_mac_1_byte_6_reg_en);
    
    \APB3_RDATA_1_bm[5]\ : CFG4
      generic map(INIT => x"CFEF")

      port map(A => APB3_RDATA_1_sn_m8_out, B => \N_455_i\, C => 
        \read_reg_en\, D => \APB3_RDATA_1_bm_1[5]_net_1\, Y => 
        \APB3_RDATA_1_bm[5]_net_1\);
    
    mac_3_byte_2_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_354, ALn => N_480_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_3_byte_2_reg_en\);
    
    write_reg_en : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => N_480_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \write_reg_en\);
    
    \APB3_RDATA_1_d_a1[0]\ : CFG4
      generic map(INIT => x"A280")

      port map(A => APB3_RDATA_1_sn_N_25, B => 
        APB3_RDATA_1_sn_N_14, C => N_1737, D => N_1745, Y => 
        \APB3_RDATA_1_d_a1[0]_net_1\);
    
    \APB3_RDATA_1_am_1[1]\ : CFG3
      generic map(INIT => x"47")

      port map(A => N_1738, B => APB3_RDATA_1_sn_N_14, C => 
        N_1746, Y => \APB3_RDATA_1_am_1[1]_net_1\);
    
    \mac_1_byte_1_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_1_reg[3]_net_1\);
    
    \APB3_RDATA_1_d_RNO[6]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \APB3_RDATA_1_27_d_3[6]_net_1\, B => 
        APB3_RDATA_1_sn_N_31_mux, C => 
        \APB3_RDATA_1_27_d_1[6]_net_1\, Y => 
        \APB3_RDATA_1_d_RNO[6]_net_1\);
    
    \mac_4_byte_4_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_4_reg[5]_net_1\);
    
    \RX_PACKET_DEPTH_STATUS_PROC.un1_RX_packet_depthlto7_5\ : 
        CFG4
      generic map(INIT => x"0001")

      port map(A => \RX_packet_depth[3]_net_1\, B => 
        \RX_packet_depth[2]_net_1\, C => 
        \RX_packet_depth[1]_net_1\, D => 
        \RX_packet_depth[0]_net_1\, Y => 
        un1_RX_packet_depthlto7_5);
    
    \REG_WRITE_PROC.un12_int_mask_reg_en\ : CFG4
      generic map(INIT => x"FAFC")

      port map(A => mac_4_byte_6_reg_en_1, B => \int_mask_reg_en\, 
        C => N_804, D => N_339, Y => N_803);
    
    \i_int_mask_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_int_mask_reg_en_i_i_a2, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \i_int_mask_reg[6]_net_1\);
    
    \mac_2_byte_3_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_3_reg[7]_net_1\);
    
    \APB3_RDATA_1_17_0_wmux_0[7]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_17_0_0_y0[7]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_1_byte_1_reg[7]_net_1\, D => 
        \mac_3_byte_5_reg[7]_net_1\, FCI => 
        \APB3_RDATA_1_17_0_0_co0[7]\, S => OPEN, Y => N_1687, FCO
         => OPEN);
    
    \mac_4_byte_6_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_6_reg[3]_net_1\);
    
    \mac_2_byte_3_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_3_reg[1]_net_1\);
    
    \RX_PACKET_DEPTH_STATUS_PROC.rx_packet_depth_status2\ : CFG4
      generic map(INIT => x"7707")

      port map(A => un1_RX_packet_depthlto7_5, B => 
        un1_RX_packet_depthlto7_4, C => iup_EOP_net_1, D => 
        RX_packet_depth_status_net_1, Y => 
        rx_packet_depth_status2);
    
    \iAPB3_READY_RNIJKOT[0]\ : CFG3
      generic map(INIT => x"EA")

      port map(A => \iAPB3_READYrs[0]\, B => un5_apb3_rst_rs, C
         => long_reset_set, Y => \iAPB3_READY[0]_net_1\);
    
    \APB3_RDATA_1_27_d_3[6]\ : CFG4
      generic map(INIT => x"2075")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => RX_FIFO_DOUT(6), D
         => \APB3_RDATA_1_27_d_3_1[6]_net_1\, Y => 
        \APB3_RDATA_1_27_d_3[6]_net_1\);
    
    APB3_RDATA_1_sn_m19_0 : CFG3
      generic map(INIT => x"E4")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CoreAPB3_0_APBmslave0_PADDR(7), C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => 
        \APB3_RDATA_1_sn_m19_0\);
    
    \APB3_RDATA_1_18_0_wmux_0[0]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_18_0_0_y0[0]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_5_reg[0]_net_1\, D => 
        \mac_4_byte_6_reg[0]_net_1\, FCI => 
        \APB3_RDATA_1_18_0_0_co0[0]\, S => OPEN, Y => N_116, FCO
         => OPEN);
    
    \mac_1_byte_6_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type3_reg[5]\);
    
    mac_2_byte_1_reg_en_ret_7 : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        N_480_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        mac_4_byte_6_reg_en_1_reto_0);
    
    \up_EOP_sync[1]\ : SLE
      port map(D => \up_EOP_sync[0]_net_1\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => VCC_net_1, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \up_EOP_sync[1]_net_1\);
    
    read_reg_en_RNIJAKE : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        \read_reg_en\, Y => APB3_RDATA_1_sn_m8_out);
    
    \mac_3_byte_1_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_1_reg[4]_net_1\);
    
    \i_int_mask_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_int_mask_reg_en_i_i_a2, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \i_int_mask_reg[0]_net_1\);
    
    \READ_FIFO_ENABLE_PROC.un109_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_200, D => N_201, Y
         => N_336);
    
    \APB3_RDATA_1_25_0_0_wmux[3]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_1_byte_5_reg[3]_net_1\, D => 
        \mac_2_byte_1_reg[3]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_25_0_0_y0[3]\, FCO => 
        \APB3_RDATA_1_25_0_0_co0[3]\);
    
    \APB3_RDATA_1_28_RNO[4]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \APB3_RDATA_1_25_0_wmux_0_Y[4]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \APB3_RDATA_1_25_3[4]_net_1\, Y => N_1749);
    
    \mac_1_byte_4_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type2_reg[4]\);
    
    \APB3_RDATA_1_21_0_0_wmux[1]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_2_byte_4_reg[1]_net_1\, D => 
        \mac_2_byte_6_reg[1]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_21_0_0_y0[1]\, FCO => 
        \APB3_RDATA_1_21_0_0_co0[1]\);
    
    mac_3_byte_5_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_357, ALn => N_480_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_3_byte_5_reg_en\);
    
    \APB3_RDATA_1_22[7]\ : CFG4
      generic map(INIT => x"2075")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), C => RX_FIFO_DOUT(7), D
         => \APB3_RDATA_1_22_1_0[7]_net_1\, Y => N_1727);
    
    \mac_1_byte_6_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type3_reg[0]\);
    
    \APB3_RDATA[0]\ : SLE
      port map(D => \APB3_RDATA_1[0]_net_1\, CLK => 
        \APB3_RDATA_31_sqmuxa_i\, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => VCC_net_1, Q => 
        CoreAPB3_0_APBmslave0_PRDATA(0));
    
    \mac_1_byte_1_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_1_reg[5]_net_1\);
    
    mac_4_byte_1_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_359, ALn => N_480_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_4_byte_1_reg_en\);
    
    \mac_3_byte_6_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_6_reg[1]_net_1\);
    
    \mac_3_byte_1_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_1_reg[0]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un37_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"2000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_199, D => N_201, Y
         => N_347);
    
    \scratch_pad_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \write_scratch_reg_en\, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \scratch_pad_reg[6]_net_1\);
    
    \mac_4_byte_1_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_1_reg[7]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_4_byte_5_reg_en_0_a2_0_o2\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \mac_4_byte_4_reg_en\, B => 
        \mac_4_byte_3_reg_en\, C => \mac_4_byte_2_reg_en\, Y => 
        N_156);
    
    \APB3_RDATA_1_bm_1[5]\ : CFG3
      generic map(INIT => x"1D")

      port map(A => \int_reg[5]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_2_reg[5]_net_1\, Y => 
        \APB3_RDATA_1_bm_1[5]_net_1\);
    
    \REG_WRITE_PROC.un12_mac_2_byte_1_reg_en_16_0\ : CFG4
      generic map(INIT => x"FFCA")

      port map(A => \mac_1_byte_2_reg_en\, B => 
        mac_4_byte_6_reg_en_1, C => N_342, D => N_7, Y => 
        un12_mac_2_byte_1_reg_en_16_0);
    
    \mac_3_byte_6_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_6_reg[7]_net_1\);
    
    \APB3_RDATA_1_25_0_0_wmux[4]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_1_byte_5_reg[4]_net_1\, D => 
        \mac_2_byte_1_reg[4]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_25_0_0_y0[4]\, FCO => 
        \APB3_RDATA_1_25_0_0_co0[4]\);
    
    \APB3_RDATA_1_25_4_wmux_1[7]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => N_57, D => N_1571, 
        FCI => \APB3_RDATA_1_25_4_0_co1[7]\, S => OPEN, Y => 
        \APB3_RDATA_1_25_4_y0_0[7]\, FCO => 
        \APB3_RDATA_1_25_4_co0_0[7]\);
    
    \APB3_RDATA_1_21_0_wmux_0[0]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_21_0_0_y0[0]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \consumer_type1_reg[0]\, D => \consumer_type2_reg[0]\, 
        FCI => \APB3_RDATA_1_21_0_0_co0[0]\, S => OPEN, Y => 
        N_1712, FCO => OPEN);
    
    \WRITE_REGISTER_ENABLE_PROC.un17_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"4000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_200, D => N_202, Y
         => N_342);
    
    \mac_1_byte_1_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_1_reg[2]_net_1\);
    
    \APB3_RDATA_1_26[0]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_1712, B => N_116, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_1753);
    
    \mac_4_byte_2_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_2_reg[0]_net_1\);
    
    \APB3_RDATA_1_0_0[7]\ : CFG4
      generic map(INIT => x"2F0F")

      port map(A => N_1671, B => APB3_RDATA_1_sn_N_10, C => 
        \read_reg_en\, D => CoreAPB3_0_APBmslave0_PADDR(2), Y => 
        \APB3_RDATA_1_0_0[7]_net_1\);
    
    \APB3_RDATA_1_25_4_0_wmux[7]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_1_byte_5_reg[7]_net_1\, D => 
        \mac_2_byte_1_reg[7]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_25_4_0_y0[7]\, FCO => 
        \APB3_RDATA_1_25_4_0_co0[7]\);
    
    \APB3_RDATA_1_1[3]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \mac_3_byte_6_reg[3]_net_1\, B => 
        \mac_3_byte_2_reg[3]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_561);
    
    \mac_1_byte_4_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type2_reg[1]\);
    
    \WRITE_REGISTER_ENABLE_PROC.un21_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"2000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_200, D => N_202, Y
         => N_343);
    
    \REG_WRITE_PROC.un13_mac_4_byte_2_reg_en_0_a2_3_a2_0\ : CFG3
      generic map(INIT => x"20")

      port map(A => N_414, B => \mac_2_byte_1_reg_en\, C => N_413, 
        Y => N_420);
    
    \REG_WRITE_PROC.un12_mac_2_byte_1_reg_en_16_RNIH70G\ : CFG2
      generic map(INIT => x"E")

      port map(A => N_796, B => \mac_4_byte_6_reg_en\, Y => 
        un1_control_reg_en_2_i_0_0_o2_0);
    
    \mac_3_byte_2_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_2_reg[5]_net_1\);
    
    \APB3_RDATA_1_22_bm[0]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => RX_FIFO_DOUT(0), B => RX_FIFO_Empty, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => 
        \APB3_RDATA_1_22_bm[0]_net_1\);
    
    \mac_1_byte_4_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type2_reg[0]\);
    
    \REG_WRITE_PROC.un13_mac_3_byte_4_reg_en_0_a2_1_a2\ : CFG4
      generic map(INIT => x"0040")

      port map(A => \mac_3_byte_3_reg_en\, B => 
        \mac_3_byte_4_reg_en\, C => N_420, D => N_141, Y => 
        un13_mac_3_byte_4_reg_en);
    
    \APB3_RDATA_1_18_0_wmux_0[1]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_18_0_0_y0[1]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_5_reg[1]_net_1\, D => 
        \mac_4_byte_6_reg[1]_net_1\, FCI => 
        \APB3_RDATA_1_18_0_0_co0[1]\, S => OPEN, Y => N_117, FCO
         => OPEN);
    
    \RX_packet_depth[6]\ : SLE
      port map(D => \RX_packet_depth_s[6]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_1528_i, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RX_packet_depth[6]_net_1\);
    
    mac_2_byte_1_reg_en_ret_3 : SLE
      port map(D => un12_mac_2_byte_1_reg_en_16_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        N_480_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        un12_mac_2_byte_1_reg_en_16_1_reto);
    
    \APB3_RDATA_1_21_0_wmux_0[1]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_21_0_0_y0[1]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \consumer_type1_reg[1]\, D => \consumer_type2_reg[1]\, 
        FCI => \APB3_RDATA_1_21_0_0_co0[1]\, S => OPEN, Y => 
        N_1713, FCO => OPEN);
    
    \mac_3_byte_1_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_1_reg[6]_net_1\);
    
    \APB3_RDATA_1_ns_1[1]\ : CFG4
      generic map(INIT => x"3305")

      port map(A => APB3_RDATA_1_sn_N_32_mux, B => 
        \APB3_RDATA_1_am_1[1]_net_1\, C => 
        APB3_RDATA_1_sn_N_31_mux, D => APB3_RDATA_1_sn_N_33_mux, 
        Y => \APB3_RDATA_1_ns_1[1]_net_1\);
    
    \mac_4_byte_3_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_3_reg[0]_net_1\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \mac_1_byte_4_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type2_reg[5]\);
    
    \APB3_RDATA_1_d_a0[0]\ : CFG4
      generic map(INIT => x"2000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        APB3_RDATA_1_sn_N_25, C => \mac_4_byte_2_reg[0]_net_1\, D
         => CoreAPB3_0_APBmslave0_PADDR(2), Y => 
        \APB3_RDATA_1_d_a0[0]_net_1\);
    
    \RX_packet_depth[2]\ : SLE
      port map(D => \RX_packet_depth_s[2]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_1528_i, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RX_packet_depth[2]_net_1\);
    
    \APB3_RDATA_1_18_0_0_wmux[3]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_3_reg[3]_net_1\, D => 
        \mac_4_byte_4_reg[3]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_18_0_0_y0[3]\, FCO => 
        \APB3_RDATA_1_18_0_0_co0[3]\);
    
    mac_2_byte_1_reg_en_ret_2 : SLE
      port map(D => un12_mac_2_byte_1_reg_en_16_0, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        N_480_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        un12_mac_2_byte_1_reg_en_16_0_reto);
    
    \APB3_RDATA_1_18_0_0_wmux[0]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        CoreAPB3_0_APBmslave0_PADDR(3), C => 
        \mac_4_byte_3_reg[0]_net_1\, D => 
        \mac_4_byte_4_reg[0]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_18_0_0_y0[0]\, FCO => 
        \APB3_RDATA_1_18_0_0_co0[0]\);
    
    \APB3_RDATA_1_17_0_wmux_0[5]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_17_0_0_y0[5]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_1_byte_1_reg[5]_net_1\, D => 
        \mac_3_byte_5_reg[5]_net_1\, FCI => 
        \APB3_RDATA_1_17_0_0_co0[5]\, S => OPEN, Y => N_1685, FCO
         => OPEN);
    
    mac_2_byte_3_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_349, ALn => N_480_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_2_byte_3_reg_en\);
    
    \iAPB3_READY[0]\ : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => un5_apb3_rst_i, ADn => VCC_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \iAPB3_READYrs[0]\);
    
    \mac_1_byte_6_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type3_reg[3]\);
    
    mac_1_byte_3_reg_en_0 : CFG3
      generic map(INIT => x"CA")

      port map(A => \mac_1_byte_3_reg_en\, B => 
        mac_4_byte_6_reg_en_1, C => N_343, Y => N_7);
    
    mac_1_byte_2_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_342, ALn => N_480_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_1_byte_2_reg_en\);
    
    \RX_packet_depth_cry[4]\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \RX_packet_depth[4]_net_1\, B => 
        rx_packet_complt, C => GND_net_1, D => GND_net_1, FCI => 
        \RX_packet_depth_cry[3]_net_1\, S => 
        \RX_packet_depth_s[4]\, Y => OPEN, FCO => 
        \RX_packet_depth_cry[4]_net_1\);
    
    \APB3_RDATA_1_s[7]\ : CFG4
      generic map(INIT => x"CFDF")

      port map(A => APB3_RDATA_1_sn_i6_mux, B => \N_455_i\, C => 
        \read_reg_en\, D => APB3_RDATA_1_sn_N_25, Y => 
        \APB3_RDATA_1_s[7]_net_1\);
    
    \mac_3_byte_6_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_6_reg[4]_net_1\);
    
    \APB3_RDATA_1_1[1]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \mac_3_byte_6_reg[1]_net_1\, B => 
        \mac_3_byte_2_reg[1]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_559);
    
    \REG_WRITE_PROC.un13_mac_4_byte_4_reg_en_0_a2_0_a2\ : CFG4
      generic map(INIT => x"1000")

      port map(A => \mac_1_byte_2_reg_en\, B => 
        \mac_1_byte_1_reg_en\, C => N_553, D => 
        un13_mac_4_byte_4_reg_en_0_a2_0_a2_1, Y => 
        un13_mac_4_byte_4_reg_en);
    
    \mac_2_byte_5_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_5_reg[0]_net_1\);
    
    \control_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => control_reg_22, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \control_reg_3\);
    
    \control_reg_RNO[5]\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PWDATA(5), B => 
        \control_reg_en\, Y => N_456_i);
    
    \WRITE_REGISTER_ENABLE_PROC.un69_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"2000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_199, D => N_212, Y
         => N_355);
    
    \mac_4_byte_5_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_5_reg[3]_net_1\);
    
    \i_int_mask_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => 
        un13_int_mask_reg_en_i_i_a2, ALn => long_reset_i, ADn => 
        VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \i_int_mask_reg[1]_net_1\);
    
    APB3_RDATA_1_4 : CFG4
      generic map(INIT => x"B080")

      port map(A => N_1744, B => APB3_RDATA_1_sn_N_14, C => 
        APB3_RDATA_1_sn_N_33_mux, D => N_1752, Y => 
        \APB3_RDATA_1_4\);
    
    \APB3_RDATA_1_17_0_wmux_0[3]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_17_0_0_y0[3]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_1_byte_1_reg[3]_net_1\, D => 
        \mac_3_byte_5_reg[3]_net_1\, FCI => 
        \APB3_RDATA_1_17_0_0_co0[3]\, S => OPEN, Y => N_1683, FCO
         => OPEN);
    
    \APB3_RDATA_1_21_0_wmux_0[6]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_21_0_0_y0[6]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \consumer_type1_reg[6]\, D => \consumer_type2_reg[6]\, 
        FCI => \APB3_RDATA_1_21_0_0_co0[6]\, S => OPEN, Y => 
        N_1718, FCO => OPEN);
    
    \WRITE_REGISTER_ENABLE_PROC.un89_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_199, D => N_202, Y
         => N_360);
    
    \APB3_RDATA_1_17_0_wmux_0[2]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_17_0_0_y0[2]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_1_byte_1_reg[2]_net_1\, D => 
        \mac_3_byte_5_reg[2]_net_1\, FCI => 
        \APB3_RDATA_1_17_0_0_co0[2]\, S => OPEN, Y => N_1682, FCO
         => OPEN);
    
    \WRITE_REGISTER_ENABLE_PROC.un65_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"4000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_199, D => N_212, Y
         => N_354);
    
    \mac_4_byte_5_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_5_reg[6]_net_1\);
    
    \APB3_RDATA_1_17_0_wmux_0[4]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_17_0_0_y0[4]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_1_byte_1_reg[4]_net_1\, D => 
        \mac_3_byte_5_reg[4]_net_1\, FCI => 
        \APB3_RDATA_1_17_0_0_co0[4]\, S => OPEN, Y => N_1684, FCO
         => OPEN);
    
    \APB3_RDATA[3]\ : SLE
      port map(D => \APB3_RDATA_1[3]_net_1\, CLK => 
        \APB3_RDATA_31_sqmuxa_i\, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => VCC_net_1, Q => 
        CoreAPB3_0_APBmslave0_PRDATA(3));
    
    \WRITE_REGISTER_ENABLE_PROC.un89_apb3_addr_0_a2_0\ : CFG2
      generic map(INIT => x"8")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_202);
    
    \APB3_RDATA_1_1_0[7]\ : CFG4
      generic map(INIT => x"3035")

      port map(A => \N_455_i\, B => N_1760, C => 
        APB3_RDATA_1_sn_N_32_mux, D => 
        \APB3_RDATA_1_0_1[7]_net_1\, Y => 
        \APB3_RDATA_1_1[7]_net_1\);
    
    \mac_3_byte_6_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_6_reg[2]_net_1\);
    
    APB3_RDATA_31_sqmuxa_i : CFG4
      generic map(INIT => x"F7F5")

      port map(A => \read_reg_en\, B => N_1805, C => \N_455_i\, D
         => \APB3_RDATA_31_sqmuxa_i_1\, Y => 
        \APB3_RDATA_31_sqmuxa_i\);
    
    \APB3_RDATA_1_17_0_wmux_0[6]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_17_0_0_y0[6]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_1_byte_1_reg[6]_net_1\, D => 
        \mac_3_byte_5_reg[6]_net_1\, FCI => 
        \APB3_RDATA_1_17_0_0_co0[6]\, S => OPEN, Y => N_1686, FCO
         => OPEN);
    
    \mac_1_byte_1_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_1_reg[7]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un85_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"2000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_199, D => N_202, Y
         => N_359);
    
    \REG_WRITE_PROC.un12_mac_2_byte_1_reg_en_16\ : CFG4
      generic map(INIT => x"FFFE")

      port map(A => un12_mac_2_byte_1_reg_en_16_2_reto, B => 
        un12_mac_2_byte_1_reg_en_16_1_reto, C => 
        un12_mac_2_byte_1_reg_en_16_0_reto, D => N_802, Y => 
        N_796);
    
    \REG_WRITE_PROC.un13_mac_4_byte_1_reg_en_0_a2_0_a2_1\ : CFG4
      generic map(INIT => x"0200")

      port map(A => \mac_4_byte_1_reg_en\, B => 
        \mac_3_byte_6_reg_en\, C => \mac_3_byte_5_reg_en\, D => 
        N_420, Y => un13_mac_4_byte_1_reg_en_0_a2_0_a2_1);
    
    mac_3_byte_1_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_353, ALn => N_480_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_3_byte_1_reg_en\);
    
    mac_1_byte_5_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_345, ALn => N_480_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_1_byte_5_reg_en\);
    
    \APB3_RDATA_1_24[2]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_1682, B => CoreAPB3_0_APBmslave0_PADDR(3), 
        C => N_1698, Y => N_1739);
    
    \APB3_RDATA_1_28[6]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => N_1743, B => APB3_RDATA_1_sn_N_14, C => 
        N_1751, Y => N_1778);
    
    \APB3_RDATA[6]\ : SLE
      port map(D => \APB3_RDATA_1[6]_net_1\, CLK => 
        \APB3_RDATA_31_sqmuxa_i\, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => VCC_net_1, Q => 
        CoreAPB3_0_APBmslave0_PRDATA(6));
    
    \mac_1_byte_2_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type1_reg[0]\);
    
    \APB3_RDATA_1_29_d_1[6]\ : CFG3
      generic map(INIT => x"53")

      port map(A => N_1718, B => N_122, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => 
        \APB3_RDATA_1_29_d_1[6]_net_1\);
    
    \mac_2_byte_5_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_5_reg[7]_net_1\);
    
    \APB3_RDATA_1_21_0_0_wmux[3]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_2_byte_4_reg[3]_net_1\, D => 
        \mac_2_byte_6_reg[3]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_21_0_0_y0[3]\, FCO => 
        \APB3_RDATA_1_21_0_0_co0[3]\);
    
    \APB3_RDATA_1_17_0_0_wmux[5]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => \start_tx_FIFO\, D
         => \mac_2_byte_3_reg[5]_net_1\, FCI => VCC_net_1, S => 
        OPEN, Y => \APB3_RDATA_1_17_0_0_y0[5]\, FCO => 
        \APB3_RDATA_1_17_0_0_co0[5]\);
    
    \scratch_pad_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \write_scratch_reg_en\, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \scratch_pad_reg[1]_net_1\);
    
    \APB3_RDATA_1_26[1]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_1713, B => N_117, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_1754);
    
    \WRITE_REGISTER_ENABLE_PROC.un73_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_199, D => N_212, Y
         => N_356);
    
    \REG_WRITE_PROC.un13_mac_1_byte_2_reg_en_0_a2_0_a2\ : CFG3
      generic map(INIT => x"08")

      port map(A => \mac_1_byte_2_reg_en\, B => N_407, C => 
        \mac_1_byte_1_reg_en\, Y => un13_mac_1_byte_2_reg_en);
    
    N_479_i : CFG4
      generic map(INIT => x"0040")

      port map(A => CoreAPB3_0_APBmslave0_PWRITE, B => 
        CoreAPB3_0_APBmslave0_PSELx, C => 
        CoreAPB3_0_APBmslave0_PENABLE, D => long_reset, Y => 
        N_479_i_i);
    
    \RX_packet_depth_s[7]\ : ARI1
      generic map(INIT => x"49900")

      port map(A => VCC_net_1, B => \RX_packet_depth[7]_net_1\, C
         => rx_packet_complt, D => GND_net_1, FCI => 
        \RX_packet_depth_cry[6]_net_1\, S => 
        \RX_packet_depth_s[7]_net_1\, Y => OPEN, FCO => OPEN);
    
    \control_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => control_reg_22, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \TX_FIFO_RST\);
    
    \mac_2_byte_5_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_5_reg[4]_net_1\);
    
    \APB3_RDATA_1_1[2]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \mac_3_byte_6_reg[2]_net_1\, B => 
        \mac_3_byte_2_reg[2]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_560);
    
    \mac_3_byte_2_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_2_reg[6]_net_1\);
    
    \mac_3_byte_2_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_2_reg[1]_net_1\);
    
    \mac_1_byte_3_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type2_reg[8]\);
    
    \APB3_RDATA_1_1[4]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \mac_3_byte_6_reg[4]_net_1\, B => 
        \mac_3_byte_2_reg[4]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_562);
    
    \APB3_RDATA_1_28_RNO[2]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \APB3_RDATA_1_25_0_wmux_0_Y[2]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \APB3_RDATA_1_25_3[2]_net_1\, Y => N_1747);
    
    \mac_3_byte_1_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_1_reg[3]_net_1\);
    
    mac_4_byte_3_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_361, ALn => N_480_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_4_byte_3_reg_en\);
    
    \APB3_RDATA_1_21_0_0_wmux[4]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_2_byte_4_reg[4]_net_1\, D => 
        \mac_2_byte_6_reg[4]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_21_0_0_y0[4]\, FCO => 
        \APB3_RDATA_1_21_0_0_co0[4]\);
    
    \APB3_RDATA_1_d_am[3]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_1715, B => N_119, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => 
        \APB3_RDATA_1_d_am[3]_net_1\);
    
    \APB3_RDATA_1_25_3[6]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_56, B => CoreAPB3_0_APBmslave0_PADDR(3), C
         => N_1570, Y => \APB3_RDATA_1_25_3[6]_net_1\);
    
    \APB3_RDATA_1_24[4]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_1684, B => CoreAPB3_0_APBmslave0_PADDR(3), 
        C => N_1700, Y => N_1741);
    
    \mac_4_byte_2_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_2_reg[7]_net_1\);
    
    \APB3_RDATA_1_3[2]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \consumer_type4_reg[2]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_4_reg[2]_net_1\, Y => N_1566);
    
    \mac_2_byte_6_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_6_reg[6]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un93_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"0008")

      port map(A => N_201, B => un105_apb3_addr_0_a2_0_1, C => 
        CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => N_361);
    
    int_mask_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_339, ALn => N_480_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \int_mask_reg_en\);
    
    \APB3_RDATA_1_24[0]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_1680, B => CoreAPB3_0_APBmslave0_PADDR(3), 
        C => N_1696, Y => N_1737);
    
    \APB3_RDATA_1_0_1[7]\ : CFG4
      generic map(INIT => x"F8F0")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(2), B => 
        APB3_RDATA_1_sn_N_10, C => \APB3_RDATA_1_0_0[7]_net_1\, D
         => N_1727, Y => \APB3_RDATA_1_0_1[7]_net_1\);
    
    \READY_DELAY_PROC.un5_apb3_rst_rs\ : SLE
      port map(D => VCC_net_1, CLK => long_reset, EN => VCC_net_1, 
        ALn => un5_apb3_rst_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => VCC_net_1, Q => un5_apb3_rst_rs);
    
    \APB3_RDATA_1_d_ns[3]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \APB3_RDATA_1_d_bm[3]_net_1\, B => 
        APB3_RDATA_1_sn_N_33_mux, C => 
        \APB3_RDATA_1_d_am[3]_net_1\, Y => 
        \APB3_RDATA_1_d_ns[3]_net_1\);
    
    \scratch_pad_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \write_scratch_reg_en\, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \scratch_pad_reg[0]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_1_byte_2_reg_en_0_a2_0_a2_0\ : CFG3
      generic map(INIT => x"01")

      port map(A => \control_reg_en\, B => \write_scratch_reg_en\, 
        C => \int_mask_reg_en\, Y => N_407);
    
    \mac_1_byte_5_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_5_reg[3]_net_1\);
    
    \mac_3_byte_6_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_6_reg[5]_net_1\);
    
    \mac_2_byte_4_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_4_reg[2]_net_1\);
    
    \control_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => control_reg_22, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \control_reg_0\);
    
    \APB3_RDATA_1_25_0_0_wmux[2]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_1_byte_5_reg[2]_net_1\, D => 
        \mac_2_byte_1_reg[2]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_25_0_0_y0[2]\, FCO => 
        \APB3_RDATA_1_25_0_0_co0[2]\);
    
    \mac_4_byte_3_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_3_reg[7]_net_1\);
    
    \APB3_RDATA_1_1[5]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \mac_3_byte_6_reg[5]_net_1\, B => 
        \mac_3_byte_2_reg[5]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_55);
    
    iTX_FIFO_wr_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un1_apb3_addr, ALn => 
        N_480_i_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => TX_FIFO_wr_en);
    
    \APB3_RDATA_1_d_0[0]\ : CFG4
      generic map(INIT => x"FFEF")

      port map(A => \N_455_i\, B => \APB3_RDATA_1_d_a1[0]_net_1\, 
        C => \read_reg_en\, D => \APB3_RDATA_1_d_a0[0]_net_1\, Y
         => \APB3_RDATA_1_d_0[0]_net_1\);
    
    \control_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => control_reg_22, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \external_loopback\);
    
    \RX_packet_depth_cry[3]\ : ARI1
      generic map(INIT => x"5AA55")

      port map(A => \RX_packet_depth[3]_net_1\, B => 
        rx_packet_complt, C => GND_net_1, D => GND_net_1, FCI => 
        \RX_packet_depth_cry[2]_net_1\, S => 
        \RX_packet_depth_s[3]\, Y => OPEN, FCO => 
        \RX_packet_depth_cry[3]_net_1\);
    
    \mac_4_byte_3_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_3_reg[1]_net_1\);
    
    \APB3_RDATA_1[6]\ : CFG4
      generic map(INIT => x"F1E0")

      port map(A => APB3_RDATA_1_sn_N_33_mux, B => 
        \APB3_RDATA_1_29_s[6]_net_1\, C => 
        \APB3_RDATA_1_d[6]_net_1\, D => 
        \APB3_RDATA_1_29_d[6]_net_1\, Y => 
        \APB3_RDATA_1[6]_net_1\);
    
    \control_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => control_reg_22, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \control_reg_2\);
    
    \APB3_RDATA_1_17_0_0_wmux[2]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => \control_reg_2\, D
         => \mac_2_byte_3_reg[2]_net_1\, FCI => VCC_net_1, S => 
        OPEN, Y => \APB3_RDATA_1_17_0_0_y0[2]\, FCO => 
        \APB3_RDATA_1_17_0_0_co0[2]\);
    
    \mac_2_byte_3_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_3_reg[5]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un105_apb3_addr_0_a2_0_1\ : CFG4
      generic map(INIT => x"0004")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CoreAPB3_0_APBmslave0_PADDR(7), C => 
        CoreAPB3_0_APBmslave0_PADDR(1), D => 
        CoreAPB3_0_APBmslave0_PADDR(0), Y => 
        un105_apb3_addr_0_a2_0_1);
    
    \mac_3_byte_4_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_4_reg[4]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un29_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"1000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_199, D => N_201, Y
         => N_345);
    
    \mac_1_byte_5_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_5_reg[6]_net_1\);
    
    \mac_3_byte_6_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_6_reg[0]_net_1\);
    
    \APB3_RDATA_1_3[4]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \consumer_type4_reg[4]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_4_reg[4]_net_1\, Y => N_1568);
    
    \APB3_RDATA_1_d_a1_RNO[0]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => \APB3_RDATA_1_25_0_wmux_0_Y[0]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => 
        \APB3_RDATA_1_25_3[0]_net_1\, Y => N_1745);
    
    \APB3_RDATA_1_29_d_bm[5]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_1717, B => N_121, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => 
        \APB3_RDATA_1_29_d_bm[5]_net_1\);
    
    \mac_3_byte_1_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_1_reg[5]_net_1\);
    
    \APB3_RDATA_1_19_0_0_wmux[5]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \i_int_mask_reg[5]_net_1\, D => 
        \mac_1_byte_3_reg[5]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_19_0_0_y0[5]\, FCO => 
        \APB3_RDATA_1_19_0_0_co0[5]\);
    
    \mac_2_byte_5_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_5_reg[5]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un25_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"8000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_200, D => N_202, Y
         => N_344);
    
    \APB3_RDATA_1_25_0_wmux_0[2]\ : ARI1
      generic map(INIT => x"0F588")

      port map(A => \APB3_RDATA_1_25_0_0_y0[2]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => 
        \mac_3_byte_1_reg[2]_net_1\, D => 
        \mac_3_byte_3_reg[2]_net_1\, FCI => 
        \APB3_RDATA_1_25_0_0_co0[2]\, S => OPEN, Y => 
        \APB3_RDATA_1_25_0_wmux_0_Y[2]\, FCO => OPEN);
    
    \APB3_RDATA_1_28[5]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => N_1742, B => APB3_RDATA_1_sn_N_14, C => 
        N_1750, Y => N_1777);
    
    \REG_WRITE_PROC.un13_mac_4_byte_2_reg_en_0_a2_3_a2\ : CFG4
      generic map(INIT => x"0020")

      port map(A => \mac_4_byte_2_reg_en\, B => 
        un13_mac_4_byte_2_reg_en_0_a2_3_o2_0, C => N_420, D => 
        N_146, Y => un13_mac_4_byte_2_reg_en);
    
    \REG_WRITE_PROC.un13_mac_2_byte_6_reg_en_0_a2_1_a2\ : CFG4
      generic map(INIT => x"0040")

      port map(A => \mac_2_byte_5_reg_en\, B => 
        \mac_2_byte_6_reg_en\, C => N_420, D => N_129, Y => 
        un13_mac_2_byte_6_reg_en);
    
    \APB3_RDATA_1_1[6]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \mac_3_byte_6_reg[6]_net_1\, B => 
        \mac_3_byte_2_reg[6]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_56);
    
    \mac_3_byte_1_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_1_reg[2]_net_1\);
    
    \APB3_RDATA[2]\ : SLE
      port map(D => \APB3_RDATA_1[2]\, CLK => 
        \APB3_RDATA_31_sqmuxa_i\, EN => VCC_net_1, ALn => 
        VCC_net_1, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => VCC_net_1, Q => 
        CoreAPB3_0_APBmslave0_PRDATA(2));
    
    \mac_3_byte_4_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_4_reg[1]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_3_byte_5_reg_en_0_a2_1_a2\ : CFG3
      generic map(INIT => x"08")

      port map(A => \mac_3_byte_5_reg_en\, B => N_420, C => N_146, 
        Y => un13_mac_3_byte_5_reg_en);
    
    mac_1_byte_1_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_341, ALn => N_480_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_1_byte_1_reg_en\);
    
    \mac_3_byte_4_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_4_reg[0]_net_1\);
    
    control_reg_22_0_0_a2_0 : CFG4
      generic map(INIT => x"0C88")

      port map(A => TX_PreAmble, B => \control_reg_en\, C => 
        \write_scratch_reg_en\, D => N_160, Y => control_reg_22);
    
    \APB3_RDATA_1_4[2]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => \consumer_type3_reg[2]\, B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \scratch_pad_reg[2]_net_1\, Y => N_1576);
    
    \scratch_pad_reg[2]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(2), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \write_scratch_reg_en\, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \scratch_pad_reg[2]_net_1\);
    
    \APB3_RDATA_1_bm_1[2]\ : CFG3
      generic map(INIT => x"1B")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => N_1576, 
        C => N_1658, Y => \APB3_RDATA_1_bm_1[2]_net_1\);
    
    \up_EOP_sync_RNIOGPQ[2]\ : CFG3
      generic map(INIT => x"9C")

      port map(A => \up_EOP_sync[1]_net_1\, B => rx_packet_complt, 
        C => \up_EOP_sync[2]_net_1\, Y => N_1528_i);
    
    \RX_packet_depth[3]\ : SLE
      port map(D => \RX_packet_depth_s[3]\, CLK => 
        CommsFPGA_CCC_0_GL0, EN => N_1528_i, ALn => long_reset_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \RX_packet_depth[3]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un1_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"2000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_200, D => N_201, Y
         => un1_apb3_addr);
    
    \mac_2_byte_1_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_1_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type4_reg[9]\);
    
    \REG_WRITE_PROC.un13_mac_4_byte_6_reg_en_0_a2_4_a2_0\ : CFG4
      generic map(INIT => x"0010")

      port map(A => \mac_2_byte_1_reg_en\, B => 
        un13_mac_4_byte_2_reg_en_0_a2_3_o2_0, C => N_413, D => 
        N_146, Y => N_553);
    
    read_reg_en : SLE
      port map(D => VCC_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => N_479_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \read_reg_en\);
    
    INTERRUPT_INST : Interrupts
      port map(CoreAPB3_0_APBmslave0_PADDR(3) => 
        CoreAPB3_0_APBmslave0_PADDR(3), 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        CoreAPB3_0_APBmslave0_PADDR(2), 
        CoreAPB3_0_APBmslave0_PWDATA(7) => 
        CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), int_reg(7) => int_reg(7), 
        int_reg(6) => int_reg(6), int_reg(5) => \int_reg[5]\, 
        int_reg(4) => \int_reg[4]\, int_reg(3) => \int_reg[3]\, 
        int_reg(2) => \int_reg[2]\, int_reg(1) => \int_reg[1]\, 
        i_int_mask_reg(7) => \i_int_mask_reg[7]_net_1\, 
        i_int_mask_reg(6) => \i_int_mask_reg[6]_net_1\, 
        i_int_mask_reg(5) => \i_int_mask_reg[5]_net_1\, 
        i_int_mask_reg(4) => \i_int_mask_reg[4]_net_1\, 
        i_int_mask_reg(3) => \i_int_mask_reg[3]_net_1\, 
        i_int_mask_reg(2) => \i_int_mask_reg[2]_net_1\, 
        i_int_mask_reg(1) => \i_int_mask_reg[1]_net_1\, 
        up_EOP_del(5) => up_EOP_del(5), up_EOP_del(4) => 
        up_EOP_del(4), up_EOP_del(3) => up_EOP_del(3), 
        up_EOP_del(2) => up_EOP_del(2), up_EOP_del(1) => 
        up_EOP_del(1), up_EOP_del(0) => up_EOP_del(0), N_218 => 
        N_218, write_reg_en => \write_reg_en\, 
        CommsFPGA_top_0_INT => CommsFPGA_top_0_INT, RESET => 
        RESET, int_reg_clr => int_reg_clr, long_reset => 
        long_reset, RX_packet_depth_status => 
        RX_packet_depth_status_net_1, tx_packet_complt_int => 
        tx_packet_complt_int, TX_FIFO_UNDERRUN => 
        TX_FIFO_UNDERRUN, un15_int_reg_clr => un15_int_reg_clr, 
        TX_FIFO_UNDERRUN_set => TX_FIFO_UNDERRUN_set, 
        TX_FIFO_OVERFLOW => TX_FIFO_OVERFLOW, un19_int_reg_clr
         => un19_int_reg_clr, TX_FIFO_OVERFLOW_set => 
        TX_FIFO_OVERFLOW_set, RX_FIFO_UNDERRUN => 
        RX_FIFO_UNDERRUN, un23_int_reg_clr => un23_int_reg_clr, 
        rx_FIFO_UNDERRUN_int => rx_FIFO_UNDERRUN_int, 
        RX_FIFO_UNDERRUN_set => RX_FIFO_UNDERRUN_set, 
        RX_FIFO_OVERFLOW => RX_FIFO_OVERFLOW, un27_int_reg_clr
         => un27_int_reg_clr, rx_FIFO_OVERFLOW_int => 
        rx_FIFO_OVERFLOW_int, RX_FIFO_OVERFLOW_set => 
        RX_FIFO_OVERFLOW_set, rx_CRC_error => rx_CRC_error, 
        un31_int_reg_clr => un31_int_reg_clr, rx_CRC_error_int
         => rx_CRC_error_int, rx_CRC_error_set => 
        rx_CRC_error_set, rx_packet_avail_int => 
        \rx_packet_avail_int\, tx_packet_complt => 
        tx_packet_complt, iup_EOP => iup_EOP_net_1, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, RESET_i => 
        RESET_i, block_int_until_rd => block_int_until_rd);
    
    \mac_2_byte_5_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_5_reg[1]_net_1\);
    
    \mac_3_byte_4_reg[5]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(5), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_4_reg[5]_net_1\);
    
    mac_3_byte_3_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_355, ALn => N_480_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_3_byte_3_reg_en\);
    
    \mac_1_byte_2_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_2_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type1_reg[7]\);
    
    \RX_packet_depth_status\ : SLE
      port map(D => rx_packet_depth_status2, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => VCC_net_1, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => 
        RX_packet_depth_status_net_1);
    
    \WRITE_REGISTER_ENABLE_PROC.un53_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"0800")

      port map(A => APB3_RDATA_1_sn_N_18, B => N_199, C => 
        CoreAPB3_0_APBmslave0_PADDR(2), D => 
        CoreAPB3_0_APBmslave0_PADDR(3), Y => N_351);
    
    \REG_WRITE_PROC.un13_mac_4_byte_3_reg_en_0_a2_4_a2_2\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \int_mask_reg_en\, B => \mac_4_byte_2_reg_en\, 
        C => N_813, D => \mac_4_byte_3_reg_en\, Y => 
        un13_mac_4_byte_3_reg_en_0_a2_4_a2_2);
    
    \APB3_RDATA_1_1[7]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \mac_3_byte_6_reg[7]_net_1\, B => 
        \mac_3_byte_2_reg[7]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_57);
    
    \APB3_RDATA_1_19_0_0_wmux[2]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(6), C => 
        \i_int_mask_reg[2]_net_1\, D => 
        \mac_1_byte_3_reg[2]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_19_0_0_y0[2]\, FCO => 
        \APB3_RDATA_1_19_0_0_co0[2]\);
    
    \mac_3_byte_6_reg[3]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(3), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_3_byte_6_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_3_byte_6_reg[3]_net_1\);
    
    \APB3_RDATA_1_1[0]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => \mac_3_byte_6_reg[0]_net_1\, B => 
        \mac_3_byte_2_reg[0]_net_1\, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_558);
    
    \APB3_RDATA_1_17_0_0_wmux[7]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => \TX_FIFO_RST\, D => 
        \mac_2_byte_3_reg[7]_net_1\, FCI => VCC_net_1, S => OPEN, 
        Y => \APB3_RDATA_1_17_0_0_y0[7]\, FCO => 
        \APB3_RDATA_1_17_0_0_co0[7]\);
    
    \REG_WRITE_PROC.un13_mac_1_byte_3_reg_en_0_a2_0_a2\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_414, B => \mac_1_byte_3_reg_en\, Y => 
        un13_mac_1_byte_3_reg_en);
    
    \scratch_pad_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => \write_scratch_reg_en\, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \scratch_pad_reg[4]_net_1\);
    
    \APB3_RDATA_1_14[3]\ : CFG3
      generic map(INIT => x"CA")

      port map(A => RX_FIFO_DOUT(3), B => TX_FIFO_Full, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_1659);
    
    \APB3_RDATA_1_25_3[2]\ : CFG3
      generic map(INIT => x"E2")

      port map(A => N_560, B => CoreAPB3_0_APBmslave0_PADDR(3), C
         => N_1566, Y => \APB3_RDATA_1_25_3[2]_net_1\);
    
    \mac_1_byte_3_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_1_byte_3_reg[7]_net_1\);
    
    \control_reg[4]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(4), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => control_reg_22, ALn => 
        long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, SD => 
        GND_net_1, LAT => GND_net_1, Q => \internal_loopback\);
    
    \mac_1_byte_3_reg[1]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(1), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_1_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \consumer_type2_reg[9]\);
    
    \REG_WRITE_PROC.un13_mac_3_byte_1_reg_en_0_a2_1_o2\ : CFG3
      generic map(INIT => x"FE")

      port map(A => \mac_2_byte_6_reg_en\, B => 
        \mac_2_byte_5_reg_en\, C => N_129, Y => N_131);
    
    \APB3_RDATA_1_29_d[6]\ : CFG4
      generic map(INIT => x"AFEF")

      port map(A => \N_455_i\, B => APB3_RDATA_1_sn_N_32_mux, C
         => \read_reg_en\, D => \APB3_RDATA_1_29_d_1[6]_net_1\, Y
         => \APB3_RDATA_1_29_d[6]_net_1\);
    
    \APB3_RDATA_1_26[7]\ : CFG3
      generic map(INIT => x"AC")

      port map(A => N_1719, B => N_123, C => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_1760);
    
    \mac_2_byte_4_reg[7]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(7), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_4_reg[7]_net_1\);
    
    \REG_WRITE_PROC.un13_mac_1_byte_1_reg_en_0_a2_2_a2\ : CFG2
      generic map(INIT => x"8")

      port map(A => N_407, B => \mac_1_byte_1_reg_en\, Y => 
        un13_mac_1_byte_1_reg_en);
    
    \mac_2_byte_4_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_4_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_4_reg[6]_net_1\);
    
    mac_2_byte_1_reg_en_ret_6 : SLE
      port map(D => N_803, CLK => m2s010_som_sb_0_CCC_71MHz, EN
         => VCC_net_1, ALn => N_480_i_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        N_803_reto);
    
    \APB3_RDATA_1_am[2]\ : CFG3
      generic map(INIT => x"B8")

      port map(A => N_1774, B => APB3_RDATA_1_sn_N_33_mux, C => 
        N_1755, Y => \APB3_RDATA_1_am[2]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un41_apb3_addr_0_a2_0\ : CFG2
      generic map(INIT => x"1")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(5), B => 
        CoreAPB3_0_APBmslave0_PADDR(4), Y => N_201);
    
    \mac_2_byte_3_reg[6]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(6), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_2_byte_3_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_2_byte_3_reg[6]_net_1\);
    
    mac_2_byte_6_reg_en : SLE
      port map(D => mac_4_byte_6_reg_en_1, CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => N_352, ALn => N_480_i_i, 
        ADn => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT
         => GND_net_1, Q => \mac_2_byte_6_reg_en\);
    
    \up_EOP_sync[0]\ : SLE
      port map(D => iup_EOP_net_1, CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => long_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \up_EOP_sync[0]_net_1\);
    
    \APB3_RDATA_1_17_0_0_wmux[4]\ : ARI1
      generic map(INIT => x"0FA44")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(6), B => 
        CoreAPB3_0_APBmslave0_PADDR(5), C => \internal_loopback\, 
        D => \mac_2_byte_3_reg[4]_net_1\, FCI => VCC_net_1, S => 
        OPEN, Y => \APB3_RDATA_1_17_0_0_y0[4]\, FCO => 
        \APB3_RDATA_1_17_0_0_co0[4]\);
    
    \mac_4_byte_5_reg[0]\ : SLE
      port map(D => CoreAPB3_0_APBmslave0_PWDATA(0), CLK => 
        m2s010_som_sb_0_CCC_71MHz, EN => un13_mac_4_byte_5_reg_en, 
        ALn => long_reset_i, ADn => VCC_net_1, SLn => VCC_net_1, 
        SD => GND_net_1, LAT => GND_net_1, Q => 
        \mac_4_byte_5_reg[0]_net_1\);
    
    \WRITE_REGISTER_ENABLE_PROC.un77_apb3_addr_0_a2\ : CFG4
      generic map(INIT => x"1000")

      port map(A => CoreAPB3_0_APBmslave0_PADDR(3), B => 
        CoreAPB3_0_APBmslave0_PADDR(2), C => N_199, D => N_202, Y
         => N_357);
    
    \REG_WRITE_PROC.un13_mac_3_byte_3_reg_en_0_a2_1_a2\ : CFG3
      generic map(INIT => x"08")

      port map(A => N_420, B => \mac_3_byte_3_reg_en\, C => N_141, 
        Y => un13_mac_3_byte_3_reg_en);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity CommsFPGA_top is

    port( packet_available_clear_reg         : out   std_logic_vector(2 downto 0);
          ReadFIFO_Read_Ptr                  : out   std_logic_vector(1 downto 0);
          ReadFIFO_Write_Ptr                 : out   std_logic_vector(1 downto 0);
          iRX_FIFO_Empty                     : out   std_logic_vector(3 downto 0);
          iRX_FIFO_UNDERRUN                  : out   std_logic_vector(3 downto 0);
          iRX_FIFO_Full                      : out   std_logic_vector(3 downto 0);
          CoreAPB3_0_APBmslave0_PRDATA_m     : out   std_logic_vector(7 downto 0);
          un15                               : out   std_logic_vector(10 downto 0);
          RX_FIFO_DIN                        : out   std_logic_vector(7 downto 0);
          RX_FIFO_DIN_pipe                   : out   std_logic_vector(8 downto 0);
          clkdiv                             : out   std_logic_vector(3 downto 0);
          un6                                : out   std_logic_vector(5 downto 0);
          p2s_data                           : out   std_logic_vector(7 downto 0);
          manches_in_dly                     : out   std_logic_vector(1 downto 0);
          CoreAPB3_0_APBmslave0_PWDATA       : in    std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PRDATA       : out   std_logic_vector(7 downto 0);
          RX_packet_depth                    : out   std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PADDR        : in    std_logic_vector(7 downto 0);
          RX_FIFO_DOUT                       : out   std_logic_vector(8 downto 0);
          int_reg                            : out   std_logic_vector(7 downto 1);
          up_EOP_del                         : out   std_logic_vector(5 downto 0);
          DEBOUNCE_IN_c                      : in    std_logic_vector(2 downto 0);
          Y_net_0                            : in    std_logic_vector(3 downto 1);
          control_reg_0                      : out   std_logic;
          control_reg_2                      : out   std_logic;
          control_reg_3                      : out   std_logic;
          DEBOUNCE_OUT_net_0_0               : out   std_logic;
          CoreAPB3_0_APBmslave0_PREADY_i_m_i : out   std_logic;
          MANCHESTER_IN_c                    : in    std_logic;
          irx_center_sample                  : out   std_logic;
          iNRZ_data                          : out   std_logic;
          MANCH_OUT_P_c                      : out   std_logic;
          MANCH_OUT_P_c_i                    : out   std_logic;
          DRVR_EN_c                          : out   std_logic;
          iup_EOP                            : out   std_logic;
          long_reset_set                     : in    std_logic;
          CoreAPB3_0_APBmslave0_PREADY       : out   std_logic;
          external_loopback                  : out   std_logic;
          internal_loopback                  : out   std_logic;
          start_tx_FIFO                      : out   std_logic;
          TX_FIFO_RST                        : out   std_logic;
          N_480_i_i                          : in    std_logic;
          RX_FIFO_rd_en                      : out   std_logic;
          TX_FIFO_wr_en                      : out   std_logic;
          RX_packet_depth_status             : out   std_logic;
          rx_packet_complt                   : out   std_logic;
          rx_packet_avail_int                : out   std_logic;
          TX_FIFO_Full                       : out   std_logic;
          TX_FIFO_Empty                      : out   std_logic;
          CoreAPB3_0_APBmslave0_PSELx        : in    std_logic;
          CoreAPB3_0_APBmslave0_PENABLE      : in    std_logic;
          RX_FIFO_Full                       : out   std_logic;
          RX_FIFO_Empty                      : out   std_logic;
          CoreAPB3_0_APBmslave0_PWRITE       : in    std_logic;
          N_480_i                            : out   std_logic;
          CommsFPGA_top_0_INT                : out   std_logic;
          int_reg_clr                        : out   std_logic;
          rx_FIFO_UNDERRUN_int               : out   std_logic;
          rx_FIFO_OVERFLOW_int               : out   std_logic;
          rx_CRC_error_int                   : out   std_logic;
          tx_packet_complt                   : out   std_logic;
          block_int_until_rd                 : out   std_logic;
          RESET_set                          : in    std_logic;
          DEBOUNCE_OUT_1_c                   : out   std_logic;
          DEBOUNCE_OUT_2_c                   : out   std_logic;
          CommsFPGA_top_0_CAMERA_NODE        : out   std_logic;
          CommsFPGA_CCC_0_LOCK               : in    std_logic;
          m2s010_som_sb_0_POWER_ON_RESET_N   : in    std_logic;
          m2s010_som_sb_0_GPIO_28_SW_RESET   : in    std_logic;
          rx_FIFO_rst_reg                    : out   std_logic;
          CommsFPGA_CCC_0_GL1                : in    std_logic;
          CommsFPGA_CCC_0_GL0                : in    std_logic;
          m2s010_som_sb_0_CCC_71MHz          : in    std_logic;
          long_reset_i                       : out   std_logic;
          RESET_i                            : out   std_logic;
          RESET                              : out   std_logic;
          BIT_CLK                            : out   std_logic;
          long_reset                         : out   std_logic;
          bd_reset                           : out   std_logic
        );

end CommsFPGA_top;

architecture DEF_ARCH of CommsFPGA_top is 

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG3
    generic (INIT:std_logic_vector(7 downto 0) := x"00");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CFG2
    generic (INIT:std_logic_vector(3 downto 0) := x"0");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CFG4
    generic (INIT:std_logic_vector(15 downto 0) := x"0000");

    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          D : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ARI1
    generic (INIT:std_logic_vector(19 downto 0) := x"00000");

    port( A   : in    std_logic := 'U';
          B   : in    std_logic := 'U';
          C   : in    std_logic := 'U';
          D   : in    std_logic := 'U';
          FCI : in    std_logic := 'U';
          S   : out   std_logic;
          Y   : out   std_logic;
          FCO : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component CFG1
    generic (INIT:std_logic_vector(1 downto 0) := "00");

    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component TriDebounce
    port( DEBOUNCE_IN_c        : in    std_logic_vector(2 downto 0) := (others => 'U');
          DEBOUNCE_OUT_net_0_0 : out   std_logic;
          DEBOUNCE_OUT_2_c     : out   std_logic;
          DEBOUNCE_OUT_1_c     : out   std_logic;
          BIT_CLK              : in    std_logic := 'U';
          RESET_set            : in    std_logic := 'U';
          RESET                : in    std_logic := 'U'
        );
  end component;

  component ManchesEncoder
    port( manches_in_dly      : in    std_logic_vector(1 downto 0) := (others => 'U');
          TX_FIFO_DOUT        : in    std_logic_vector(7 downto 0) := (others => 'U');
          p2s_data            : out   std_logic_vector(7 downto 0);
          start_tx_FIFO       : in    std_logic := 'U';
          TX_FIFO_Empty       : in    std_logic := 'U';
          N_114               : out   std_logic;
          idle_line5          : out   std_logic;
          tx_col_detect_en    : out   std_logic;
          CommsFPGA_CCC_0_GL0 : in    std_logic := 'U';
          DRVR_EN_c           : out   std_logic;
          internal_loopback   : in    std_logic := 'U';
          external_loopback   : in    std_logic := 'U';
          tx_packet_complt    : out   std_logic;
          RESET               : in    std_logic := 'U';
          TX_PreAmble         : out   std_logic;
          CommsFPGA_CCC_0_GL1 : in    std_logic := 'U';
          byte_clk_en         : in    std_logic := 'U';
          BIT_CLK             : in    std_logic := 'U';
          RESET_i             : in    std_logic := 'U';
          MANCH_OUT_P_c_i     : out   std_logic;
          MANCH_OUT_P_c       : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component ManchesDecoder
    port( un6                                : out   std_logic_vector(5 downto 0);
          manches_in_dly                     : out   std_logic_vector(1 downto 0);
          clkdiv                             : out   std_logic_vector(3 downto 0);
          RX_FIFO_DIN_pipe                   : out   std_logic_vector(8 downto 0);
          RX_FIFO_DIN                        : out   std_logic_vector(7 downto 0);
          un15                               : out   std_logic_vector(10 downto 0);
          CoreAPB3_0_APBmslave0_PRDATA       : in    std_logic_vector(7 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PRDATA_m     : out   std_logic_vector(7 downto 0);
          consumer_type2_reg                 : in    std_logic_vector(9 downto 0) := (others => 'U');
          consumer_type1_reg                 : in    std_logic_vector(9 downto 0) := (others => 'U');
          consumer_type3_reg                 : in    std_logic_vector(9 downto 0) := (others => 'U');
          consumer_type4_reg                 : in    std_logic_vector(9 downto 0) := (others => 'U');
          iNRZ_data                          : out   std_logic;
          irx_center_sample                  : out   std_logic;
          internal_loopback                  : in    std_logic := 'U';
          MANCH_OUT_P_c                      : in    std_logic := 'U';
          MANCHESTER_IN_c                    : in    std_logic := 'U';
          idle_line5                         : in    std_logic := 'U';
          rx_CRC_error                       : out   std_logic;
          rx_CRC_error_i                     : out   std_logic;
          CommsFPGA_CCC_0_GL0                : in    std_logic := 'U';
          RESET_i                            : in    std_logic := 'U';
          RX_EarlyTerm                       : out   std_logic;
          rx_packet_complt                   : out   std_logic;
          CoreAPB3_0_APBmslave0_PSELx        : in    std_logic := 'U';
          tx_col_detect_en                   : in    std_logic := 'U';
          RX_FIFO_TxColDetDis_wr_en          : out   std_logic;
          RESET                              : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PREADY       : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PREADY_i_m_i : out   std_logic;
          DRVR_EN_c                          : in    std_logic := 'U'
        );
  end component;

  component FIFOs
    port( RX_FIFO_DIN_pipe             : in    std_logic_vector(8 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PWDATA : in    std_logic_vector(7 downto 0) := (others => 'U');
          TX_FIFO_DOUT                 : out   std_logic_vector(7 downto 0);
          up_EOP_sync                  : in    std_logic_vector(2 downto 1) := (others => 'U');
          RX_FIFO_DOUT                 : out   std_logic_vector(8 downto 0);
          iRX_FIFO_Full                : out   std_logic_vector(3 downto 0);
          iRX_FIFO_UNDERRUN            : out   std_logic_vector(3 downto 0);
          iRX_FIFO_Empty               : out   std_logic_vector(3 downto 0);
          ReadFIFO_Write_Ptr           : out   std_logic_vector(1 downto 0);
          ReadFIFO_Read_Ptr            : out   std_logic_vector(1 downto 0);
          packet_available_clear_reg   : out   std_logic_vector(2 downto 0);
          RX_FIFO_TxColDetDis_wr_en    : in    std_logic := 'U';
          TX_FIFO_UNDERRUN             : out   std_logic;
          TX_FIFO_UNDERRUN_i           : out   std_logic;
          TX_FIFO_OVERFLOW             : out   std_logic;
          TX_FIFO_OVERFLOW_i           : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz    : in    std_logic := 'U';
          TX_FIFO_Full                 : out   std_logic;
          TX_FIFO_wr_en                : in    std_logic := 'U';
          TX_FIFO_Empty                : out   std_logic;
          N_114                        : in    std_logic := 'U';
          BIT_CLK                      : in    std_logic := 'U';
          RX_FIFO_RST                  : in    std_logic := 'U';
          TX_FIFO_RST                  : in    std_logic := 'U';
          RESET                        : in    std_logic := 'U';
          RX_FIFO_rd_en                : in    std_logic := 'U';
          rx_packet_complt             : in    std_logic := 'U';
          RX_FIFO_Full                 : out   std_logic;
          RX_FIFO_Empty                : out   std_logic;
          rx_packet_avail_int          : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0          : in    std_logic := 'U';
          RX_FIFO_OVERFLOW_i           : out   std_logic;
          RX_FIFO_OVERFLOW             : out   std_logic;
          RX_FIFO_UNDERRUN_i           : out   std_logic;
          RX_FIFO_UNDERRUN             : out   std_logic
        );
  end component;

  component uP_if
    port( up_EOP_del                    : out   std_logic_vector(5 downto 0);
          int_reg                       : out   std_logic_vector(7 downto 1);
          RX_FIFO_DOUT                  : in    std_logic_vector(8 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PADDR   : in    std_logic_vector(7 downto 0) := (others => 'U');
          RX_packet_depth               : out   std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PRDATA  : out   std_logic_vector(7 downto 0);
          consumer_type4_reg            : out   std_logic_vector(9 downto 0);
          consumer_type3_reg            : out   std_logic_vector(9 downto 0);
          consumer_type2_reg            : out   std_logic_vector(9 downto 0);
          consumer_type1_reg            : out   std_logic_vector(9 downto 0);
          CoreAPB3_0_APBmslave0_PWDATA  : in    std_logic_vector(7 downto 0) := (others => 'U');
          up_EOP_sync                   : out   std_logic_vector(2 downto 1);
          control_reg_0                 : out   std_logic;
          control_reg_2                 : out   std_logic;
          control_reg_3                 : out   std_logic;
          block_int_until_rd            : out   std_logic;
          RESET_i                       : in    std_logic := 'U';
          tx_packet_complt              : in    std_logic := 'U';
          rx_CRC_error_set              : in    std_logic := 'U';
          rx_CRC_error_int              : out   std_logic;
          un31_int_reg_clr              : out   std_logic;
          rx_CRC_error                  : in    std_logic := 'U';
          RX_FIFO_OVERFLOW_set          : in    std_logic := 'U';
          rx_FIFO_OVERFLOW_int          : out   std_logic;
          un27_int_reg_clr              : out   std_logic;
          RX_FIFO_OVERFLOW              : in    std_logic := 'U';
          RX_FIFO_UNDERRUN_set          : in    std_logic := 'U';
          rx_FIFO_UNDERRUN_int          : out   std_logic;
          un23_int_reg_clr              : out   std_logic;
          RX_FIFO_UNDERRUN              : in    std_logic := 'U';
          TX_FIFO_OVERFLOW_set          : in    std_logic := 'U';
          un19_int_reg_clr              : out   std_logic;
          TX_FIFO_OVERFLOW              : in    std_logic := 'U';
          TX_FIFO_UNDERRUN_set          : in    std_logic := 'U';
          un15_int_reg_clr              : out   std_logic;
          TX_FIFO_UNDERRUN              : in    std_logic := 'U';
          int_reg_clr                   : out   std_logic;
          RESET                         : in    std_logic := 'U';
          CommsFPGA_top_0_INT           : out   std_logic;
          TX_PreAmble                   : in    std_logic := 'U';
          N_480_i                       : out   std_logic;
          CoreAPB3_0_APBmslave0_PWRITE  : in    std_logic := 'U';
          RX_FIFO_Empty                 : in    std_logic := 'U';
          RX_FIFO_Full                  : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PENABLE : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PSELx   : in    std_logic := 'U';
          TX_FIFO_Empty                 : in    std_logic := 'U';
          TX_FIFO_Full                  : in    std_logic := 'U';
          rx_packet_avail_int           : out   std_logic;
          rx_packet_complt              : in    std_logic := 'U';
          RX_packet_depth_status        : out   std_logic;
          TX_FIFO_wr_en                 : out   std_logic;
          RX_FIFO_rd_en                 : out   std_logic;
          N_480_i_i                     : in    std_logic := 'U';
          TX_FIFO_RST                   : out   std_logic;
          rx_FIFO_rst_reg               : out   std_logic;
          start_tx_FIFO                 : out   std_logic;
          internal_loopback             : out   std_logic;
          external_loopback             : out   std_logic;
          long_reset                    : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PREADY  : out   std_logic;
          m2s010_som_sb_0_CCC_71MHz     : in    std_logic := 'U';
          long_reset_set                : in    std_logic := 'U';
          iup_EOP                       : out   std_logic;
          CommsFPGA_CCC_0_GL0           : in    std_logic := 'U';
          long_reset_i                  : in    std_logic := 'U'
        );
  end component;

    signal bd_reset_net_1, bd_reset_0, long_reset_net_1, 
        long_reset_0, BIT_CLK_net_1, BIT_CLK_0, RESET_net_1, 
        RESET_0, \ClkDivider[0]_net_1\, \ClkDivider_i[0]\, 
        BIT_CLK_i_i, \RESET_i\, \long_reset_i\, bd_reset_i, 
        \rx_CRC_error_set\, GND_net_1, rx_CRC_error_i, 
        un31_int_reg_clr, VCC_net_1, \RX_FIFO_OVERFLOW_set\, 
        RX_FIFO_OVERFLOW_i, un27_int_reg_clr, 
        \RX_FIFO_UNDERRUN_set\, RX_FIFO_UNDERRUN_i, 
        un23_int_reg_clr, \TX_FIFO_OVERFLOW_set\, 
        TX_FIFO_OVERFLOW_i, un19_int_reg_clr, 
        \TX_FIFO_UNDERRUN_set\, TX_FIFO_UNDERRUN_i, 
        un15_int_reg_clr, \long_reset_cntr[0]_net_1\, 
        \long_reset_cntr_3[0]_net_1\, \long_reset_cntr[1]_net_1\, 
        \long_reset_cntr_3[1]_net_1\, \long_reset_cntr[2]_net_1\, 
        \long_reset_cntr_3[2]_net_1\, \long_reset_cntr[3]_net_1\, 
        \long_reset_cntr_3[3]_net_1\, \long_reset_cntr[4]_net_1\, 
        \long_reset_cntr_3[4]_net_1\, \long_reset_cntr[5]_net_1\, 
        \long_reset_cntr_3[5]_net_1\, \long_reset_cntr[6]_net_1\, 
        un4_long_reset_cntr_cry_6_S, \long_reset_cntr[7]_net_1\, 
        un4_long_reset_cntr_s_7_S, \ClkDivider[1]_net_1\, 
        \ClkDivider_RNO[1]_net_1\, \ClkDivider[2]_net_1\, 
        \ClkDivider_RNO[2]_net_1\, \RX_FIFO_RST\, RX_FIFO_RST_1, 
        \byte_clk_en\, byte_clk_en_1, un2_long_reset_cntr_i, 
        un4_long_reset_cntr_s_1_920_FCO, 
        \un4_long_reset_cntr_cry_1\, un4_long_reset_cntr_cry_1_S, 
        \un4_long_reset_cntr_cry_2\, un4_long_reset_cntr_cry_2_S, 
        \un4_long_reset_cntr_cry_3\, un4_long_reset_cntr_cry_3_S, 
        \un4_long_reset_cntr_cry_4\, un4_long_reset_cntr_cry_4_S, 
        \un4_long_reset_cntr_cry_5\, un4_long_reset_cntr_cry_5_S, 
        \un4_long_reset_cntr_cry_6\, RX_EarlyTerm, 
        \rx_FIFO_rst_reg\, un2_long_reset_cntr_5, 
        un2_long_reset_cntr_4, \RX_FIFO_DOUT[0]\, 
        \RX_FIFO_DOUT[1]\, \RX_FIFO_DOUT[2]\, \RX_FIFO_DOUT[3]\, 
        \RX_FIFO_DOUT[4]\, \RX_FIFO_DOUT[5]\, \RX_FIFO_DOUT[6]\, 
        \RX_FIFO_DOUT[7]\, \RX_FIFO_DOUT[8]\, 
        \CoreAPB3_0_APBmslave0_PRDATA[0]\, 
        \CoreAPB3_0_APBmslave0_PRDATA[1]\, 
        \CoreAPB3_0_APBmslave0_PRDATA[2]\, 
        \CoreAPB3_0_APBmslave0_PRDATA[3]\, 
        \CoreAPB3_0_APBmslave0_PRDATA[4]\, 
        \CoreAPB3_0_APBmslave0_PRDATA[5]\, 
        \CoreAPB3_0_APBmslave0_PRDATA[6]\, 
        \CoreAPB3_0_APBmslave0_PRDATA[7]\, 
        \consumer_type4_reg[0]\, \consumer_type4_reg[1]\, 
        \consumer_type4_reg[2]\, \consumer_type4_reg[3]\, 
        \consumer_type4_reg[4]\, \consumer_type4_reg[5]\, 
        \consumer_type4_reg[6]\, \consumer_type4_reg[7]\, 
        \consumer_type4_reg[8]\, \consumer_type4_reg[9]\, 
        \consumer_type3_reg[0]\, \consumer_type3_reg[1]\, 
        \consumer_type3_reg[2]\, \consumer_type3_reg[3]\, 
        \consumer_type3_reg[4]\, \consumer_type3_reg[5]\, 
        \consumer_type3_reg[6]\, \consumer_type3_reg[7]\, 
        \consumer_type3_reg[8]\, \consumer_type3_reg[9]\, 
        \consumer_type2_reg[0]\, \consumer_type2_reg[1]\, 
        \consumer_type2_reg[2]\, \consumer_type2_reg[3]\, 
        \consumer_type2_reg[4]\, \consumer_type2_reg[5]\, 
        \consumer_type2_reg[6]\, \consumer_type2_reg[7]\, 
        \consumer_type2_reg[8]\, \consumer_type2_reg[9]\, 
        \consumer_type1_reg[0]\, \consumer_type1_reg[1]\, 
        \consumer_type1_reg[2]\, \consumer_type1_reg[3]\, 
        \consumer_type1_reg[4]\, \consumer_type1_reg[5]\, 
        \consumer_type1_reg[6]\, \consumer_type1_reg[7]\, 
        \consumer_type1_reg[8]\, \consumer_type1_reg[9]\, 
        \up_EOP_sync[1]\, \up_EOP_sync[2]\, \tx_packet_complt\, 
        rx_CRC_error, RX_FIFO_OVERFLOW, RX_FIFO_UNDERRUN, 
        TX_FIFO_OVERFLOW, TX_FIFO_UNDERRUN, TX_PreAmble, 
        \RX_FIFO_Empty\, \RX_FIFO_Full\, \TX_FIFO_Empty\, 
        \TX_FIFO_Full\, \rx_packet_avail_int\, \rx_packet_complt\, 
        \TX_FIFO_wr_en\, \RX_FIFO_rd_en\, \TX_FIFO_RST\, 
        \start_tx_FIFO\, \internal_loopback\, \external_loopback\, 
        \CoreAPB3_0_APBmslave0_PREADY\, \manches_in_dly[0]\, 
        \manches_in_dly[1]\, \TX_FIFO_DOUT[0]\, \TX_FIFO_DOUT[1]\, 
        \TX_FIFO_DOUT[2]\, \TX_FIFO_DOUT[3]\, \TX_FIFO_DOUT[4]\, 
        \TX_FIFO_DOUT[5]\, \TX_FIFO_DOUT[6]\, \TX_FIFO_DOUT[7]\, 
        N_114, idle_line5, tx_col_detect_en, \DRVR_EN_c\, 
        \MANCH_OUT_P_c\, \RX_FIFO_DIN_pipe[0]\, 
        \RX_FIFO_DIN_pipe[1]\, \RX_FIFO_DIN_pipe[2]\, 
        \RX_FIFO_DIN_pipe[3]\, \RX_FIFO_DIN_pipe[4]\, 
        \RX_FIFO_DIN_pipe[5]\, \RX_FIFO_DIN_pipe[6]\, 
        \RX_FIFO_DIN_pipe[7]\, \RX_FIFO_DIN_pipe[8]\, 
        RX_FIFO_TxColDetDis_wr_en : std_logic;
    signal nc2, nc1 : std_logic;

    for all : TriDebounce
	Use entity work.TriDebounce(DEF_ARCH);
    for all : ManchesEncoder
	Use entity work.ManchesEncoder(DEF_ARCH);
    for all : ManchesDecoder
	Use entity work.ManchesDecoder(DEF_ARCH);
    for all : FIFOs
	Use entity work.FIFOs(DEF_ARCH);
    for all : uP_if
	Use entity work.uP_if(DEF_ARCH);
begin 

    RX_FIFO_DIN_pipe(8) <= \RX_FIFO_DIN_pipe[8]\;
    RX_FIFO_DIN_pipe(7) <= \RX_FIFO_DIN_pipe[7]\;
    RX_FIFO_DIN_pipe(6) <= \RX_FIFO_DIN_pipe[6]\;
    RX_FIFO_DIN_pipe(5) <= \RX_FIFO_DIN_pipe[5]\;
    RX_FIFO_DIN_pipe(4) <= \RX_FIFO_DIN_pipe[4]\;
    RX_FIFO_DIN_pipe(3) <= \RX_FIFO_DIN_pipe[3]\;
    RX_FIFO_DIN_pipe(2) <= \RX_FIFO_DIN_pipe[2]\;
    RX_FIFO_DIN_pipe(1) <= \RX_FIFO_DIN_pipe[1]\;
    RX_FIFO_DIN_pipe(0) <= \RX_FIFO_DIN_pipe[0]\;
    manches_in_dly(1) <= \manches_in_dly[1]\;
    manches_in_dly(0) <= \manches_in_dly[0]\;
    CoreAPB3_0_APBmslave0_PRDATA(7) <= 
        \CoreAPB3_0_APBmslave0_PRDATA[7]\;
    CoreAPB3_0_APBmslave0_PRDATA(6) <= 
        \CoreAPB3_0_APBmslave0_PRDATA[6]\;
    CoreAPB3_0_APBmslave0_PRDATA(5) <= 
        \CoreAPB3_0_APBmslave0_PRDATA[5]\;
    CoreAPB3_0_APBmslave0_PRDATA(4) <= 
        \CoreAPB3_0_APBmslave0_PRDATA[4]\;
    CoreAPB3_0_APBmslave0_PRDATA(3) <= 
        \CoreAPB3_0_APBmslave0_PRDATA[3]\;
    CoreAPB3_0_APBmslave0_PRDATA(2) <= 
        \CoreAPB3_0_APBmslave0_PRDATA[2]\;
    CoreAPB3_0_APBmslave0_PRDATA(1) <= 
        \CoreAPB3_0_APBmslave0_PRDATA[1]\;
    CoreAPB3_0_APBmslave0_PRDATA(0) <= 
        \CoreAPB3_0_APBmslave0_PRDATA[0]\;
    RX_FIFO_DOUT(8) <= \RX_FIFO_DOUT[8]\;
    RX_FIFO_DOUT(7) <= \RX_FIFO_DOUT[7]\;
    RX_FIFO_DOUT(6) <= \RX_FIFO_DOUT[6]\;
    RX_FIFO_DOUT(5) <= \RX_FIFO_DOUT[5]\;
    RX_FIFO_DOUT(4) <= \RX_FIFO_DOUT[4]\;
    RX_FIFO_DOUT(3) <= \RX_FIFO_DOUT[3]\;
    RX_FIFO_DOUT(2) <= \RX_FIFO_DOUT[2]\;
    RX_FIFO_DOUT(1) <= \RX_FIFO_DOUT[1]\;
    RX_FIFO_DOUT(0) <= \RX_FIFO_DOUT[0]\;
    MANCH_OUT_P_c <= \MANCH_OUT_P_c\;
    DRVR_EN_c <= \DRVR_EN_c\;
    CoreAPB3_0_APBmslave0_PREADY <= 
        \CoreAPB3_0_APBmslave0_PREADY\;
    external_loopback <= \external_loopback\;
    internal_loopback <= \internal_loopback\;
    start_tx_FIFO <= \start_tx_FIFO\;
    TX_FIFO_RST <= \TX_FIFO_RST\;
    RX_FIFO_rd_en <= \RX_FIFO_rd_en\;
    TX_FIFO_wr_en <= \TX_FIFO_wr_en\;
    rx_packet_complt <= \rx_packet_complt\;
    rx_packet_avail_int <= \rx_packet_avail_int\;
    TX_FIFO_Full <= \TX_FIFO_Full\;
    TX_FIFO_Empty <= \TX_FIFO_Empty\;
    RX_FIFO_Full <= \RX_FIFO_Full\;
    RX_FIFO_Empty <= \RX_FIFO_Empty\;
    tx_packet_complt <= \tx_packet_complt\;
    rx_FIFO_rst_reg <= \rx_FIFO_rst_reg\;
    long_reset_i <= \long_reset_i\;
    RESET_i <= \RESET_i\;
    RESET <= RESET_net_1;
    BIT_CLK <= BIT_CLK_net_1;
    long_reset <= long_reset_net_1;
    bd_reset <= bd_reset_net_1;

    BIT_CLK_inferred_clock_RNIT9E2 : CLKINT
      port map(A => BIT_CLK_0, Y => BIT_CLK_net_1);
    
    \long_reset_cntr_3[3]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => un2_long_reset_cntr_4, B => 
        un2_long_reset_cntr_5, C => un4_long_reset_cntr_cry_3_S, 
        Y => \long_reset_cntr_3[3]_net_1\);
    
    \bd_reset\ : CFG2
      generic map(INIT => x"B")

      port map(A => m2s010_som_sb_0_GPIO_28_SW_RESET, B => 
        m2s010_som_sb_0_POWER_ON_RESET_N, Y => bd_reset_0);
    
    \long_reset_cntr[3]\ : SLE
      port map(D => \long_reset_cntr_3[3]_net_1\, CLK => 
        BIT_CLK_net_1, EN => VCC_net_1, ALn => bd_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \long_reset_cntr[3]_net_1\);
    
    \RESET_DELAY_PROC.un2_long_reset_cntr_4\ : CFG4
      generic map(INIT => x"8000")

      port map(A => \long_reset_cntr[4]_net_1\, B => 
        \long_reset_cntr[3]_net_1\, C => 
        \long_reset_cntr[2]_net_1\, D => 
        \long_reset_cntr[1]_net_1\, Y => un2_long_reset_cntr_4);
    
    \long_reset_cntr[6]\ : SLE
      port map(D => un4_long_reset_cntr_cry_6_S, CLK => 
        BIT_CLK_net_1, EN => VCC_net_1, ALn => bd_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \long_reset_cntr[6]_net_1\);
    
    \ClkDivider_RNO[2]\ : CFG3
      generic map(INIT => x"6A")

      port map(A => \ClkDivider[2]_net_1\, B => 
        \ClkDivider[1]_net_1\, C => \ClkDivider[0]_net_1\, Y => 
        \ClkDivider_RNO[2]_net_1\);
    
    byte_clk_en : SLE
      port map(D => byte_clk_en_1, CLK => BIT_CLK_net_1, EN => 
        VCC_net_1, ALn => \RESET_i\, ADn => VCC_net_1, SLn => 
        VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \byte_clk_en\);
    
    \ClkDivider_RNO[1]\ : CFG2
      generic map(INIT => x"6")

      port map(A => \ClkDivider[0]_net_1\, B => 
        \ClkDivider[1]_net_1\, Y => \ClkDivider_RNO[1]_net_1\);
    
    \RESET_DELAY_PROC.un2_long_reset_cntr_5\ : CFG4
      generic map(INIT => x"0100")

      port map(A => \long_reset_cntr[7]_net_1\, B => 
        \long_reset_cntr[6]_net_1\, C => 
        \long_reset_cntr[5]_net_1\, D => 
        \long_reset_cntr[0]_net_1\, Y => un2_long_reset_cntr_5);
    
    un4_long_reset_cntr_cry_2 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \long_reset_cntr[2]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un4_long_reset_cntr_cry_1\, S => 
        un4_long_reset_cntr_cry_2_S, Y => OPEN, FCO => 
        \un4_long_reset_cntr_cry_2\);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    \ID_RES_DECODE_PROC.un4_id_res\ : CFG3
      generic map(INIT => x"08")

      port map(A => Y_net_0(3), B => Y_net_0(2), C => Y_net_0(1), 
        Y => CommsFPGA_top_0_CAMERA_NODE);
    
    un4_long_reset_cntr_s_1_920 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \long_reset_cntr[0]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => VCC_net_1, S => 
        OPEN, Y => OPEN, FCO => un4_long_reset_cntr_s_1_920_FCO);
    
    RESET_RNIFEG6 : CLKINT
      port map(A => RESET_0, Y => RESET_net_1);
    
    \ClkDivider_RNO[0]\ : CFG1
      generic map(INIT => "01")

      port map(A => \ClkDivider[0]_net_1\, Y => \ClkDivider_i[0]\);
    
    \long_reset_cntr[5]\ : SLE
      port map(D => \long_reset_cntr_3[5]_net_1\, CLK => 
        BIT_CLK_net_1, EN => VCC_net_1, ALn => bd_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \long_reset_cntr[5]_net_1\);
    
    TRIPLE_DEBOUNCE_INST : TriDebounce
      port map(DEBOUNCE_IN_c(2) => DEBOUNCE_IN_c(2), 
        DEBOUNCE_IN_c(1) => DEBOUNCE_IN_c(1), DEBOUNCE_IN_c(0)
         => DEBOUNCE_IN_c(0), DEBOUNCE_OUT_net_0_0 => 
        DEBOUNCE_OUT_net_0_0, DEBOUNCE_OUT_2_c => 
        DEBOUNCE_OUT_2_c, DEBOUNCE_OUT_1_c => DEBOUNCE_OUT_1_c, 
        BIT_CLK => BIT_CLK_net_1, RESET_set => RESET_set, RESET
         => RESET_net_1);
    
    un4_long_reset_cntr_cry_3 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \long_reset_cntr[3]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un4_long_reset_cntr_cry_2\, S => 
        un4_long_reset_cntr_cry_3_S, Y => OPEN, FCO => 
        \un4_long_reset_cntr_cry_3\);
    
    MANCHESTER_ENCODER_INST : ManchesEncoder
      port map(manches_in_dly(1) => \manches_in_dly[1]\, 
        manches_in_dly(0) => \manches_in_dly[0]\, TX_FIFO_DOUT(7)
         => \TX_FIFO_DOUT[7]\, TX_FIFO_DOUT(6) => 
        \TX_FIFO_DOUT[6]\, TX_FIFO_DOUT(5) => \TX_FIFO_DOUT[5]\, 
        TX_FIFO_DOUT(4) => \TX_FIFO_DOUT[4]\, TX_FIFO_DOUT(3) => 
        \TX_FIFO_DOUT[3]\, TX_FIFO_DOUT(2) => \TX_FIFO_DOUT[2]\, 
        TX_FIFO_DOUT(1) => \TX_FIFO_DOUT[1]\, TX_FIFO_DOUT(0) => 
        \TX_FIFO_DOUT[0]\, p2s_data(7) => p2s_data(7), 
        p2s_data(6) => p2s_data(6), p2s_data(5) => p2s_data(5), 
        p2s_data(4) => p2s_data(4), p2s_data(3) => p2s_data(3), 
        p2s_data(2) => p2s_data(2), p2s_data(1) => p2s_data(1), 
        p2s_data(0) => p2s_data(0), start_tx_FIFO => 
        \start_tx_FIFO\, TX_FIFO_Empty => \TX_FIFO_Empty\, N_114
         => N_114, idle_line5 => idle_line5, tx_col_detect_en => 
        tx_col_detect_en, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, DRVR_EN_c => \DRVR_EN_c\, 
        internal_loopback => \internal_loopback\, 
        external_loopback => \external_loopback\, 
        tx_packet_complt => \tx_packet_complt\, RESET => 
        RESET_net_1, TX_PreAmble => TX_PreAmble, 
        CommsFPGA_CCC_0_GL1 => CommsFPGA_CCC_0_GL1, byte_clk_en
         => \byte_clk_en\, BIT_CLK => BIT_CLK_net_1, RESET_i => 
        \RESET_i\, MANCH_OUT_P_c_i => MANCH_OUT_P_c_i, 
        MANCH_OUT_P_c => \MANCH_OUT_P_c\);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \SAMPLE_5MHZ_EN_PROC.byte_clk_en_1\ : CFG3
      generic map(INIT => x"08")

      port map(A => \ClkDivider[2]_net_1\, B => 
        \ClkDivider[1]_net_1\, C => \ClkDivider[0]_net_1\, Y => 
        byte_clk_en_1);
    
    \long_reset_cntr[7]\ : SLE
      port map(D => un4_long_reset_cntr_s_7_S, CLK => 
        BIT_CLK_net_1, EN => VCC_net_1, ALn => bd_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \long_reset_cntr[7]_net_1\);
    
    \long_reset\ : SLE
      port map(D => un2_long_reset_cntr_i, CLK => BIT_CLK_net_1, 
        EN => VCC_net_1, ALn => bd_reset_i, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        long_reset_0);
    
    TX_FIFO_OVERFLOW_set : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => un19_int_reg_clr, ALn => TX_FIFO_OVERFLOW_i, ADn
         => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \TX_FIFO_OVERFLOW_set\);
    
    RX_FIFO_OVERFLOW_set : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => un27_int_reg_clr, ALn => RX_FIFO_OVERFLOW_i, ADn
         => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_OVERFLOW_set\);
    
    un4_long_reset_cntr_cry_4 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \long_reset_cntr[4]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un4_long_reset_cntr_cry_3\, S => 
        un4_long_reset_cntr_cry_4_S, Y => OPEN, FCO => 
        \un4_long_reset_cntr_cry_4\);
    
    long_reset_RNO : CFG2
      generic map(INIT => x"7")

      port map(A => un2_long_reset_cntr_5, B => 
        un2_long_reset_cntr_4, Y => un2_long_reset_cntr_i);
    
    \BIT_CLK\ : SLE
      port map(D => BIT_CLK_i_i, CLK => CommsFPGA_CCC_0_GL1, EN
         => VCC_net_1, ALn => bd_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        BIT_CLK_0);
    
    MANCHESTER_DECODER_INST : ManchesDecoder
      port map(un6(5) => un6(5), un6(4) => un6(4), un6(3) => 
        un6(3), un6(2) => un6(2), un6(1) => nc2, un6(0) => un6(0), 
        manches_in_dly(1) => \manches_in_dly[1]\, 
        manches_in_dly(0) => \manches_in_dly[0]\, clkdiv(3) => 
        clkdiv(3), clkdiv(2) => clkdiv(2), clkdiv(1) => clkdiv(1), 
        clkdiv(0) => clkdiv(0), RX_FIFO_DIN_pipe(8) => 
        \RX_FIFO_DIN_pipe[8]\, RX_FIFO_DIN_pipe(7) => 
        \RX_FIFO_DIN_pipe[7]\, RX_FIFO_DIN_pipe(6) => 
        \RX_FIFO_DIN_pipe[6]\, RX_FIFO_DIN_pipe(5) => 
        \RX_FIFO_DIN_pipe[5]\, RX_FIFO_DIN_pipe(4) => 
        \RX_FIFO_DIN_pipe[4]\, RX_FIFO_DIN_pipe(3) => 
        \RX_FIFO_DIN_pipe[3]\, RX_FIFO_DIN_pipe(2) => 
        \RX_FIFO_DIN_pipe[2]\, RX_FIFO_DIN_pipe(1) => 
        \RX_FIFO_DIN_pipe[1]\, RX_FIFO_DIN_pipe(0) => 
        \RX_FIFO_DIN_pipe[0]\, RX_FIFO_DIN(7) => RX_FIFO_DIN(7), 
        RX_FIFO_DIN(6) => RX_FIFO_DIN(6), RX_FIFO_DIN(5) => 
        RX_FIFO_DIN(5), RX_FIFO_DIN(4) => RX_FIFO_DIN(4), 
        RX_FIFO_DIN(3) => RX_FIFO_DIN(3), RX_FIFO_DIN(2) => 
        RX_FIFO_DIN(2), RX_FIFO_DIN(1) => RX_FIFO_DIN(1), 
        RX_FIFO_DIN(0) => RX_FIFO_DIN(0), un15(10) => un15(10), 
        un15(9) => un15(9), un15(8) => un15(8), un15(7) => 
        un15(7), un15(6) => nc1, un15(5) => un15(5), un15(4) => 
        un15(4), un15(3) => un15(3), un15(2) => un15(2), un15(1)
         => un15(1), un15(0) => un15(0), 
        CoreAPB3_0_APBmslave0_PRDATA(7) => 
        \CoreAPB3_0_APBmslave0_PRDATA[7]\, 
        CoreAPB3_0_APBmslave0_PRDATA(6) => 
        \CoreAPB3_0_APBmslave0_PRDATA[6]\, 
        CoreAPB3_0_APBmslave0_PRDATA(5) => 
        \CoreAPB3_0_APBmslave0_PRDATA[5]\, 
        CoreAPB3_0_APBmslave0_PRDATA(4) => 
        \CoreAPB3_0_APBmslave0_PRDATA[4]\, 
        CoreAPB3_0_APBmslave0_PRDATA(3) => 
        \CoreAPB3_0_APBmslave0_PRDATA[3]\, 
        CoreAPB3_0_APBmslave0_PRDATA(2) => 
        \CoreAPB3_0_APBmslave0_PRDATA[2]\, 
        CoreAPB3_0_APBmslave0_PRDATA(1) => 
        \CoreAPB3_0_APBmslave0_PRDATA[1]\, 
        CoreAPB3_0_APBmslave0_PRDATA(0) => 
        \CoreAPB3_0_APBmslave0_PRDATA[0]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(7) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(7), 
        CoreAPB3_0_APBmslave0_PRDATA_m(6) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(6), 
        CoreAPB3_0_APBmslave0_PRDATA_m(5) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(5), 
        CoreAPB3_0_APBmslave0_PRDATA_m(4) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(4), 
        CoreAPB3_0_APBmslave0_PRDATA_m(3) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(3), 
        CoreAPB3_0_APBmslave0_PRDATA_m(2) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(2), 
        CoreAPB3_0_APBmslave0_PRDATA_m(1) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(1), 
        CoreAPB3_0_APBmslave0_PRDATA_m(0) => 
        CoreAPB3_0_APBmslave0_PRDATA_m(0), consumer_type2_reg(9)
         => \consumer_type2_reg[9]\, consumer_type2_reg(8) => 
        \consumer_type2_reg[8]\, consumer_type2_reg(7) => 
        \consumer_type2_reg[7]\, consumer_type2_reg(6) => 
        \consumer_type2_reg[6]\, consumer_type2_reg(5) => 
        \consumer_type2_reg[5]\, consumer_type2_reg(4) => 
        \consumer_type2_reg[4]\, consumer_type2_reg(3) => 
        \consumer_type2_reg[3]\, consumer_type2_reg(2) => 
        \consumer_type2_reg[2]\, consumer_type2_reg(1) => 
        \consumer_type2_reg[1]\, consumer_type2_reg(0) => 
        \consumer_type2_reg[0]\, consumer_type1_reg(9) => 
        \consumer_type1_reg[9]\, consumer_type1_reg(8) => 
        \consumer_type1_reg[8]\, consumer_type1_reg(7) => 
        \consumer_type1_reg[7]\, consumer_type1_reg(6) => 
        \consumer_type1_reg[6]\, consumer_type1_reg(5) => 
        \consumer_type1_reg[5]\, consumer_type1_reg(4) => 
        \consumer_type1_reg[4]\, consumer_type1_reg(3) => 
        \consumer_type1_reg[3]\, consumer_type1_reg(2) => 
        \consumer_type1_reg[2]\, consumer_type1_reg(1) => 
        \consumer_type1_reg[1]\, consumer_type1_reg(0) => 
        \consumer_type1_reg[0]\, consumer_type3_reg(9) => 
        \consumer_type3_reg[9]\, consumer_type3_reg(8) => 
        \consumer_type3_reg[8]\, consumer_type3_reg(7) => 
        \consumer_type3_reg[7]\, consumer_type3_reg(6) => 
        \consumer_type3_reg[6]\, consumer_type3_reg(5) => 
        \consumer_type3_reg[5]\, consumer_type3_reg(4) => 
        \consumer_type3_reg[4]\, consumer_type3_reg(3) => 
        \consumer_type3_reg[3]\, consumer_type3_reg(2) => 
        \consumer_type3_reg[2]\, consumer_type3_reg(1) => 
        \consumer_type3_reg[1]\, consumer_type3_reg(0) => 
        \consumer_type3_reg[0]\, consumer_type4_reg(9) => 
        \consumer_type4_reg[9]\, consumer_type4_reg(8) => 
        \consumer_type4_reg[8]\, consumer_type4_reg(7) => 
        \consumer_type4_reg[7]\, consumer_type4_reg(6) => 
        \consumer_type4_reg[6]\, consumer_type4_reg(5) => 
        \consumer_type4_reg[5]\, consumer_type4_reg(4) => 
        \consumer_type4_reg[4]\, consumer_type4_reg(3) => 
        \consumer_type4_reg[3]\, consumer_type4_reg(2) => 
        \consumer_type4_reg[2]\, consumer_type4_reg(1) => 
        \consumer_type4_reg[1]\, consumer_type4_reg(0) => 
        \consumer_type4_reg[0]\, iNRZ_data => iNRZ_data, 
        irx_center_sample => irx_center_sample, internal_loopback
         => \internal_loopback\, MANCH_OUT_P_c => \MANCH_OUT_P_c\, 
        MANCHESTER_IN_c => MANCHESTER_IN_c, idle_line5 => 
        idle_line5, rx_CRC_error => rx_CRC_error, rx_CRC_error_i
         => rx_CRC_error_i, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, RESET_i => \RESET_i\, RX_EarlyTerm
         => RX_EarlyTerm, rx_packet_complt => \rx_packet_complt\, 
        CoreAPB3_0_APBmslave0_PSELx => 
        CoreAPB3_0_APBmslave0_PSELx, tx_col_detect_en => 
        tx_col_detect_en, RX_FIFO_TxColDetDis_wr_en => 
        RX_FIFO_TxColDetDis_wr_en, RESET => RESET_net_1, 
        CoreAPB3_0_APBmslave0_PREADY => 
        \CoreAPB3_0_APBmslave0_PREADY\, 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i => 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i, DRVR_EN_c => 
        \DRVR_EN_c\);
    
    \RESET\ : CFG2
      generic map(INIT => x"D")

      port map(A => CommsFPGA_CCC_0_LOCK, B => long_reset_net_1, 
        Y => RESET_0);
    
    \long_reset_cntr_3[2]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => un2_long_reset_cntr_4, B => 
        un2_long_reset_cntr_5, C => un4_long_reset_cntr_cry_2_S, 
        Y => \long_reset_cntr_3[2]_net_1\);
    
    \long_reset_cntr_3[1]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => un2_long_reset_cntr_4, B => 
        un2_long_reset_cntr_5, C => un4_long_reset_cntr_cry_1_S, 
        Y => \long_reset_cntr_3[1]_net_1\);
    
    un4_long_reset_cntr_cry_5 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \long_reset_cntr[5]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un4_long_reset_cntr_cry_4\, S => 
        un4_long_reset_cntr_cry_5_S, Y => OPEN, FCO => 
        \un4_long_reset_cntr_cry_5\);
    
    un4_long_reset_cntr_cry_6 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \long_reset_cntr[6]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un4_long_reset_cntr_cry_5\, S => 
        un4_long_reset_cntr_cry_6_S, Y => OPEN, FCO => 
        \un4_long_reset_cntr_cry_6\);
    
    rx_CRC_error_set : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => un31_int_reg_clr, ALn => rx_CRC_error_i, ADn => 
        GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \rx_CRC_error_set\);
    
    BIT_CLK_RNO : CFG1
      generic map(INIT => "01")

      port map(A => BIT_CLK_0, Y => BIT_CLK_i_i);
    
    un4_long_reset_cntr_s_7 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \long_reset_cntr[7]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        \un4_long_reset_cntr_cry_6\, S => 
        un4_long_reset_cntr_s_7_S, Y => OPEN, FCO => OPEN);
    
    long_reset_RNIUA27 : CLKINT
      port map(A => long_reset_0, Y => long_reset_net_1);
    
    bd_reset_RNIK1J6_0 : CFG1
      generic map(INIT => "01")

      port map(A => bd_reset_net_1, Y => bd_reset_i);
    
    \SYNC2_APB3_CLK_PROC.RX_FIFO_RST_1\ : CFG2
      generic map(INIT => x"E")

      port map(A => RX_EarlyTerm, B => \rx_FIFO_rst_reg\, Y => 
        RX_FIFO_RST_1);
    
    \ClkDivider[2]\ : SLE
      port map(D => \ClkDivider_RNO[2]_net_1\, CLK => 
        BIT_CLK_net_1, EN => VCC_net_1, ALn => bd_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \ClkDivider[2]_net_1\);
    
    un4_long_reset_cntr_cry_1 : ARI1
      generic map(INIT => x"4AA00")

      port map(A => VCC_net_1, B => \long_reset_cntr[1]_net_1\, C
         => GND_net_1, D => GND_net_1, FCI => 
        un4_long_reset_cntr_s_1_920_FCO, S => 
        un4_long_reset_cntr_cry_1_S, Y => OPEN, FCO => 
        \un4_long_reset_cntr_cry_1\);
    
    \long_reset_cntr_3[5]\ : CFG3
      generic map(INIT => x"70")

      port map(A => un2_long_reset_cntr_4, B => 
        un2_long_reset_cntr_5, C => un4_long_reset_cntr_cry_5_S, 
        Y => \long_reset_cntr_3[5]_net_1\);
    
    RX_FIFO_RST : SLE
      port map(D => RX_FIFO_RST_1, CLK => CommsFPGA_CCC_0_GL0, EN
         => VCC_net_1, ALn => bd_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RX_FIFO_RST\);
    
    \ClkDivider[0]\ : SLE
      port map(D => \ClkDivider_i[0]\, CLK => BIT_CLK_net_1, EN
         => VCC_net_1, ALn => bd_reset_i, ADn => VCC_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \ClkDivider[0]_net_1\);
    
    long_reset_RNIUA27_0 : CFG1
      generic map(INIT => "01")

      port map(A => long_reset_net_1, Y => \long_reset_i\);
    
    \long_reset_cntr[2]\ : SLE
      port map(D => \long_reset_cntr_3[2]_net_1\, CLK => 
        BIT_CLK_net_1, EN => VCC_net_1, ALn => bd_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \long_reset_cntr[2]_net_1\);
    
    \long_reset_cntr[1]\ : SLE
      port map(D => \long_reset_cntr_3[1]_net_1\, CLK => 
        BIT_CLK_net_1, EN => VCC_net_1, ALn => bd_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \long_reset_cntr[1]_net_1\);
    
    \long_reset_cntr_3[0]\ : CFG3
      generic map(INIT => x"B3")

      port map(A => un2_long_reset_cntr_5, B => 
        \long_reset_cntr[0]_net_1\, C => un2_long_reset_cntr_4, Y
         => \long_reset_cntr_3[0]_net_1\);
    
    \long_reset_cntr[0]\ : SLE
      port map(D => \long_reset_cntr_3[0]_net_1\, CLK => 
        BIT_CLK_net_1, EN => VCC_net_1, ALn => bd_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \long_reset_cntr[0]_net_1\);
    
    TX_FIFO_UNDERRUN_set : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => un15_int_reg_clr, ALn => TX_FIFO_UNDERRUN_i, ADn
         => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \TX_FIFO_UNDERRUN_set\);
    
    \long_reset_cntr_3[4]\ : CFG3
      generic map(INIT => x"F8")

      port map(A => un2_long_reset_cntr_4, B => 
        un2_long_reset_cntr_5, C => un4_long_reset_cntr_cry_4_S, 
        Y => \long_reset_cntr_3[4]_net_1\);
    
    FIFOS_INST : FIFOs
      port map(RX_FIFO_DIN_pipe(8) => \RX_FIFO_DIN_pipe[8]\, 
        RX_FIFO_DIN_pipe(7) => \RX_FIFO_DIN_pipe[7]\, 
        RX_FIFO_DIN_pipe(6) => \RX_FIFO_DIN_pipe[6]\, 
        RX_FIFO_DIN_pipe(5) => \RX_FIFO_DIN_pipe[5]\, 
        RX_FIFO_DIN_pipe(4) => \RX_FIFO_DIN_pipe[4]\, 
        RX_FIFO_DIN_pipe(3) => \RX_FIFO_DIN_pipe[3]\, 
        RX_FIFO_DIN_pipe(2) => \RX_FIFO_DIN_pipe[2]\, 
        RX_FIFO_DIN_pipe(1) => \RX_FIFO_DIN_pipe[1]\, 
        RX_FIFO_DIN_pipe(0) => \RX_FIFO_DIN_pipe[0]\, 
        CoreAPB3_0_APBmslave0_PWDATA(7) => 
        CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), TX_FIFO_DOUT(7) => 
        \TX_FIFO_DOUT[7]\, TX_FIFO_DOUT(6) => \TX_FIFO_DOUT[6]\, 
        TX_FIFO_DOUT(5) => \TX_FIFO_DOUT[5]\, TX_FIFO_DOUT(4) => 
        \TX_FIFO_DOUT[4]\, TX_FIFO_DOUT(3) => \TX_FIFO_DOUT[3]\, 
        TX_FIFO_DOUT(2) => \TX_FIFO_DOUT[2]\, TX_FIFO_DOUT(1) => 
        \TX_FIFO_DOUT[1]\, TX_FIFO_DOUT(0) => \TX_FIFO_DOUT[0]\, 
        up_EOP_sync(2) => \up_EOP_sync[2]\, up_EOP_sync(1) => 
        \up_EOP_sync[1]\, RX_FIFO_DOUT(8) => \RX_FIFO_DOUT[8]\, 
        RX_FIFO_DOUT(7) => \RX_FIFO_DOUT[7]\, RX_FIFO_DOUT(6) => 
        \RX_FIFO_DOUT[6]\, RX_FIFO_DOUT(5) => \RX_FIFO_DOUT[5]\, 
        RX_FIFO_DOUT(4) => \RX_FIFO_DOUT[4]\, RX_FIFO_DOUT(3) => 
        \RX_FIFO_DOUT[3]\, RX_FIFO_DOUT(2) => \RX_FIFO_DOUT[2]\, 
        RX_FIFO_DOUT(1) => \RX_FIFO_DOUT[1]\, RX_FIFO_DOUT(0) => 
        \RX_FIFO_DOUT[0]\, iRX_FIFO_Full(3) => iRX_FIFO_Full(3), 
        iRX_FIFO_Full(2) => iRX_FIFO_Full(2), iRX_FIFO_Full(1)
         => iRX_FIFO_Full(1), iRX_FIFO_Full(0) => 
        iRX_FIFO_Full(0), iRX_FIFO_UNDERRUN(3) => 
        iRX_FIFO_UNDERRUN(3), iRX_FIFO_UNDERRUN(2) => 
        iRX_FIFO_UNDERRUN(2), iRX_FIFO_UNDERRUN(1) => 
        iRX_FIFO_UNDERRUN(1), iRX_FIFO_UNDERRUN(0) => 
        iRX_FIFO_UNDERRUN(0), iRX_FIFO_Empty(3) => 
        iRX_FIFO_Empty(3), iRX_FIFO_Empty(2) => iRX_FIFO_Empty(2), 
        iRX_FIFO_Empty(1) => iRX_FIFO_Empty(1), iRX_FIFO_Empty(0)
         => iRX_FIFO_Empty(0), ReadFIFO_Write_Ptr(1) => 
        ReadFIFO_Write_Ptr(1), ReadFIFO_Write_Ptr(0) => 
        ReadFIFO_Write_Ptr(0), ReadFIFO_Read_Ptr(1) => 
        ReadFIFO_Read_Ptr(1), ReadFIFO_Read_Ptr(0) => 
        ReadFIFO_Read_Ptr(0), packet_available_clear_reg(2) => 
        packet_available_clear_reg(2), 
        packet_available_clear_reg(1) => 
        packet_available_clear_reg(1), 
        packet_available_clear_reg(0) => 
        packet_available_clear_reg(0), RX_FIFO_TxColDetDis_wr_en
         => RX_FIFO_TxColDetDis_wr_en, TX_FIFO_UNDERRUN => 
        TX_FIFO_UNDERRUN, TX_FIFO_UNDERRUN_i => 
        TX_FIFO_UNDERRUN_i, TX_FIFO_OVERFLOW => TX_FIFO_OVERFLOW, 
        TX_FIFO_OVERFLOW_i => TX_FIFO_OVERFLOW_i, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz, 
        TX_FIFO_Full => \TX_FIFO_Full\, TX_FIFO_wr_en => 
        \TX_FIFO_wr_en\, TX_FIFO_Empty => \TX_FIFO_Empty\, N_114
         => N_114, BIT_CLK => BIT_CLK_net_1, RX_FIFO_RST => 
        \RX_FIFO_RST\, TX_FIFO_RST => \TX_FIFO_RST\, RESET => 
        RESET_net_1, RX_FIFO_rd_en => \RX_FIFO_rd_en\, 
        rx_packet_complt => \rx_packet_complt\, RX_FIFO_Full => 
        \RX_FIFO_Full\, RX_FIFO_Empty => \RX_FIFO_Empty\, 
        rx_packet_avail_int => \rx_packet_avail_int\, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0, 
        RX_FIFO_OVERFLOW_i => RX_FIFO_OVERFLOW_i, 
        RX_FIFO_OVERFLOW => RX_FIFO_OVERFLOW, RX_FIFO_UNDERRUN_i
         => RX_FIFO_UNDERRUN_i, RX_FIFO_UNDERRUN => 
        RX_FIFO_UNDERRUN);
    
    PROCESSOR_INTERFACE_INST : uP_if
      port map(up_EOP_del(5) => up_EOP_del(5), up_EOP_del(4) => 
        up_EOP_del(4), up_EOP_del(3) => up_EOP_del(3), 
        up_EOP_del(2) => up_EOP_del(2), up_EOP_del(1) => 
        up_EOP_del(1), up_EOP_del(0) => up_EOP_del(0), int_reg(7)
         => int_reg(7), int_reg(6) => int_reg(6), int_reg(5) => 
        int_reg(5), int_reg(4) => int_reg(4), int_reg(3) => 
        int_reg(3), int_reg(2) => int_reg(2), int_reg(1) => 
        int_reg(1), RX_FIFO_DOUT(8) => \RX_FIFO_DOUT[8]\, 
        RX_FIFO_DOUT(7) => \RX_FIFO_DOUT[7]\, RX_FIFO_DOUT(6) => 
        \RX_FIFO_DOUT[6]\, RX_FIFO_DOUT(5) => \RX_FIFO_DOUT[5]\, 
        RX_FIFO_DOUT(4) => \RX_FIFO_DOUT[4]\, RX_FIFO_DOUT(3) => 
        \RX_FIFO_DOUT[3]\, RX_FIFO_DOUT(2) => \RX_FIFO_DOUT[2]\, 
        RX_FIFO_DOUT(1) => \RX_FIFO_DOUT[1]\, RX_FIFO_DOUT(0) => 
        \RX_FIFO_DOUT[0]\, CoreAPB3_0_APBmslave0_PADDR(7) => 
        CoreAPB3_0_APBmslave0_PADDR(7), 
        CoreAPB3_0_APBmslave0_PADDR(6) => 
        CoreAPB3_0_APBmslave0_PADDR(6), 
        CoreAPB3_0_APBmslave0_PADDR(5) => 
        CoreAPB3_0_APBmslave0_PADDR(5), 
        CoreAPB3_0_APBmslave0_PADDR(4) => 
        CoreAPB3_0_APBmslave0_PADDR(4), 
        CoreAPB3_0_APBmslave0_PADDR(3) => 
        CoreAPB3_0_APBmslave0_PADDR(3), 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        CoreAPB3_0_APBmslave0_PADDR(2), 
        CoreAPB3_0_APBmslave0_PADDR(1) => 
        CoreAPB3_0_APBmslave0_PADDR(1), 
        CoreAPB3_0_APBmslave0_PADDR(0) => 
        CoreAPB3_0_APBmslave0_PADDR(0), RX_packet_depth(7) => 
        RX_packet_depth(7), RX_packet_depth(6) => 
        RX_packet_depth(6), RX_packet_depth(5) => 
        RX_packet_depth(5), RX_packet_depth(4) => 
        RX_packet_depth(4), RX_packet_depth(3) => 
        RX_packet_depth(3), RX_packet_depth(2) => 
        RX_packet_depth(2), RX_packet_depth(1) => 
        RX_packet_depth(1), RX_packet_depth(0) => 
        RX_packet_depth(0), CoreAPB3_0_APBmslave0_PRDATA(7) => 
        \CoreAPB3_0_APBmslave0_PRDATA[7]\, 
        CoreAPB3_0_APBmslave0_PRDATA(6) => 
        \CoreAPB3_0_APBmslave0_PRDATA[6]\, 
        CoreAPB3_0_APBmslave0_PRDATA(5) => 
        \CoreAPB3_0_APBmslave0_PRDATA[5]\, 
        CoreAPB3_0_APBmslave0_PRDATA(4) => 
        \CoreAPB3_0_APBmslave0_PRDATA[4]\, 
        CoreAPB3_0_APBmslave0_PRDATA(3) => 
        \CoreAPB3_0_APBmslave0_PRDATA[3]\, 
        CoreAPB3_0_APBmslave0_PRDATA(2) => 
        \CoreAPB3_0_APBmslave0_PRDATA[2]\, 
        CoreAPB3_0_APBmslave0_PRDATA(1) => 
        \CoreAPB3_0_APBmslave0_PRDATA[1]\, 
        CoreAPB3_0_APBmslave0_PRDATA(0) => 
        \CoreAPB3_0_APBmslave0_PRDATA[0]\, consumer_type4_reg(9)
         => \consumer_type4_reg[9]\, consumer_type4_reg(8) => 
        \consumer_type4_reg[8]\, consumer_type4_reg(7) => 
        \consumer_type4_reg[7]\, consumer_type4_reg(6) => 
        \consumer_type4_reg[6]\, consumer_type4_reg(5) => 
        \consumer_type4_reg[5]\, consumer_type4_reg(4) => 
        \consumer_type4_reg[4]\, consumer_type4_reg(3) => 
        \consumer_type4_reg[3]\, consumer_type4_reg(2) => 
        \consumer_type4_reg[2]\, consumer_type4_reg(1) => 
        \consumer_type4_reg[1]\, consumer_type4_reg(0) => 
        \consumer_type4_reg[0]\, consumer_type3_reg(9) => 
        \consumer_type3_reg[9]\, consumer_type3_reg(8) => 
        \consumer_type3_reg[8]\, consumer_type3_reg(7) => 
        \consumer_type3_reg[7]\, consumer_type3_reg(6) => 
        \consumer_type3_reg[6]\, consumer_type3_reg(5) => 
        \consumer_type3_reg[5]\, consumer_type3_reg(4) => 
        \consumer_type3_reg[4]\, consumer_type3_reg(3) => 
        \consumer_type3_reg[3]\, consumer_type3_reg(2) => 
        \consumer_type3_reg[2]\, consumer_type3_reg(1) => 
        \consumer_type3_reg[1]\, consumer_type3_reg(0) => 
        \consumer_type3_reg[0]\, consumer_type2_reg(9) => 
        \consumer_type2_reg[9]\, consumer_type2_reg(8) => 
        \consumer_type2_reg[8]\, consumer_type2_reg(7) => 
        \consumer_type2_reg[7]\, consumer_type2_reg(6) => 
        \consumer_type2_reg[6]\, consumer_type2_reg(5) => 
        \consumer_type2_reg[5]\, consumer_type2_reg(4) => 
        \consumer_type2_reg[4]\, consumer_type2_reg(3) => 
        \consumer_type2_reg[3]\, consumer_type2_reg(2) => 
        \consumer_type2_reg[2]\, consumer_type2_reg(1) => 
        \consumer_type2_reg[1]\, consumer_type2_reg(0) => 
        \consumer_type2_reg[0]\, consumer_type1_reg(9) => 
        \consumer_type1_reg[9]\, consumer_type1_reg(8) => 
        \consumer_type1_reg[8]\, consumer_type1_reg(7) => 
        \consumer_type1_reg[7]\, consumer_type1_reg(6) => 
        \consumer_type1_reg[6]\, consumer_type1_reg(5) => 
        \consumer_type1_reg[5]\, consumer_type1_reg(4) => 
        \consumer_type1_reg[4]\, consumer_type1_reg(3) => 
        \consumer_type1_reg[3]\, consumer_type1_reg(2) => 
        \consumer_type1_reg[2]\, consumer_type1_reg(1) => 
        \consumer_type1_reg[1]\, consumer_type1_reg(0) => 
        \consumer_type1_reg[0]\, CoreAPB3_0_APBmslave0_PWDATA(7)
         => CoreAPB3_0_APBmslave0_PWDATA(7), 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        CoreAPB3_0_APBmslave0_PWDATA(6), 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        CoreAPB3_0_APBmslave0_PWDATA(5), 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        CoreAPB3_0_APBmslave0_PWDATA(4), 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        CoreAPB3_0_APBmslave0_PWDATA(3), 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        CoreAPB3_0_APBmslave0_PWDATA(2), 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        CoreAPB3_0_APBmslave0_PWDATA(1), 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        CoreAPB3_0_APBmslave0_PWDATA(0), up_EOP_sync(2) => 
        \up_EOP_sync[2]\, up_EOP_sync(1) => \up_EOP_sync[1]\, 
        control_reg_0 => control_reg_0, control_reg_2 => 
        control_reg_2, control_reg_3 => control_reg_3, 
        block_int_until_rd => block_int_until_rd, RESET_i => 
        \RESET_i\, tx_packet_complt => \tx_packet_complt\, 
        rx_CRC_error_set => \rx_CRC_error_set\, rx_CRC_error_int
         => rx_CRC_error_int, un31_int_reg_clr => 
        un31_int_reg_clr, rx_CRC_error => rx_CRC_error, 
        RX_FIFO_OVERFLOW_set => \RX_FIFO_OVERFLOW_set\, 
        rx_FIFO_OVERFLOW_int => rx_FIFO_OVERFLOW_int, 
        un27_int_reg_clr => un27_int_reg_clr, RX_FIFO_OVERFLOW
         => RX_FIFO_OVERFLOW, RX_FIFO_UNDERRUN_set => 
        \RX_FIFO_UNDERRUN_set\, rx_FIFO_UNDERRUN_int => 
        rx_FIFO_UNDERRUN_int, un23_int_reg_clr => 
        un23_int_reg_clr, RX_FIFO_UNDERRUN => RX_FIFO_UNDERRUN, 
        TX_FIFO_OVERFLOW_set => \TX_FIFO_OVERFLOW_set\, 
        un19_int_reg_clr => un19_int_reg_clr, TX_FIFO_OVERFLOW
         => TX_FIFO_OVERFLOW, TX_FIFO_UNDERRUN_set => 
        \TX_FIFO_UNDERRUN_set\, un15_int_reg_clr => 
        un15_int_reg_clr, TX_FIFO_UNDERRUN => TX_FIFO_UNDERRUN, 
        int_reg_clr => int_reg_clr, RESET => RESET_net_1, 
        CommsFPGA_top_0_INT => CommsFPGA_top_0_INT, TX_PreAmble
         => TX_PreAmble, N_480_i => N_480_i, 
        CoreAPB3_0_APBmslave0_PWRITE => 
        CoreAPB3_0_APBmslave0_PWRITE, RX_FIFO_Empty => 
        \RX_FIFO_Empty\, RX_FIFO_Full => \RX_FIFO_Full\, 
        CoreAPB3_0_APBmslave0_PENABLE => 
        CoreAPB3_0_APBmslave0_PENABLE, 
        CoreAPB3_0_APBmslave0_PSELx => 
        CoreAPB3_0_APBmslave0_PSELx, TX_FIFO_Empty => 
        \TX_FIFO_Empty\, TX_FIFO_Full => \TX_FIFO_Full\, 
        rx_packet_avail_int => \rx_packet_avail_int\, 
        rx_packet_complt => \rx_packet_complt\, 
        RX_packet_depth_status => RX_packet_depth_status, 
        TX_FIFO_wr_en => \TX_FIFO_wr_en\, RX_FIFO_rd_en => 
        \RX_FIFO_rd_en\, N_480_i_i => N_480_i_i, TX_FIFO_RST => 
        \TX_FIFO_RST\, rx_FIFO_rst_reg => \rx_FIFO_rst_reg\, 
        start_tx_FIFO => \start_tx_FIFO\, internal_loopback => 
        \internal_loopback\, external_loopback => 
        \external_loopback\, long_reset => long_reset_net_1, 
        CoreAPB3_0_APBmslave0_PREADY => 
        \CoreAPB3_0_APBmslave0_PREADY\, m2s010_som_sb_0_CCC_71MHz
         => m2s010_som_sb_0_CCC_71MHz, long_reset_set => 
        long_reset_set, iup_EOP => iup_EOP, CommsFPGA_CCC_0_GL0
         => CommsFPGA_CCC_0_GL0, long_reset_i => \long_reset_i\);
    
    bd_reset_RNIK1J6 : CLKINT
      port map(A => bd_reset_0, Y => bd_reset_net_1);
    
    RX_FIFO_UNDERRUN_set : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => un23_int_reg_clr, ALn => RX_FIFO_UNDERRUN_i, ADn
         => GND_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \RX_FIFO_UNDERRUN_set\);
    
    \long_reset_cntr[4]\ : SLE
      port map(D => \long_reset_cntr_3[4]_net_1\, CLK => 
        BIT_CLK_net_1, EN => VCC_net_1, ALn => bd_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \long_reset_cntr[4]_net_1\);
    
    RESET_RNIFEG6_0 : CFG1
      generic map(INIT => "01")

      port map(A => RESET_net_1, Y => \RESET_i\);
    
    \ClkDivider[1]\ : SLE
      port map(D => \ClkDivider_RNO[1]_net_1\, CLK => 
        BIT_CLK_net_1, EN => VCC_net_1, ALn => bd_reset_i, ADn
         => VCC_net_1, SLn => VCC_net_1, SD => GND_net_1, LAT => 
        GND_net_1, Q => \ClkDivider[1]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity m2s010_som is

    port( DEBOUNCE_IN           : in    std_logic_vector(2 downto 0);
          ID_RES                : in    std_logic_vector(3 downto 0);
          MAC_MII_RXD           : in    std_logic_vector(3 downto 0);
          MAC_MII_TXD           : out   std_logic_vector(3 downto 0);
          MDDR_ADDR             : out   std_logic_vector(15 downto 0);
          MDDR_BA               : out   std_logic_vector(2 downto 0);
          GPIO_1_BI             : inout std_logic_vector(0 to 0) := (others => 'Z');
          GPIO_1_BIDI           : in    std_logic_vector(0 to 0);
          GPIO_6_PAD            : inout std_logic_vector(0 to 0) := (others => 'Z');
          GPIO_7_PADI           : inout std_logic_vector(0 to 0) := (others => 'Z');
          MDDR_DM_RDQS          : inout std_logic_vector(1 downto 0) := (others => 'Z');
          MDDR_DQ               : inout std_logic_vector(15 downto 0) := (others => 'Z');
          MDDR_DQS              : inout std_logic_vector(1 downto 0) := (others => 'Z');
          SPI_1_CLK             : inout std_logic_vector(0 to 0) := (others => 'Z');
          SPI_1_SS0_CAM         : inout std_logic_vector(0 to 0) := (others => 'Z');
          SPI_1_SS0_OTH         : inout std_logic_vector(0 to 0) := (others => 'Z');
          DEVRST_N              : in    std_logic;
          MAC_MII_COL           : in    std_logic;
          MAC_MII_CRS           : in    std_logic;
          MAC_MII_RX_CLK        : in    std_logic;
          MAC_MII_RX_DV         : in    std_logic;
          MAC_MII_RX_ER         : in    std_logic;
          MAC_MII_TX_CLK        : in    std_logic;
          MANCHESTER_IN         : in    std_logic;
          MDDR_DQS_TMATCH_0_IN  : in    std_logic;
          MMUART_0_RXD_F2M      : in    std_logic;
          MMUART_1_RXD          : in    std_logic;
          PULLDOWN_R9           : in    std_logic;
          SPI_0_DI              : in    std_logic;
          SPI_1_DI_CAM          : in    std_logic;
          SPI_1_DI_OTH          : in    std_logic;
          XTL                   : in    std_logic;
          DEBOUNCE_OUT_1        : out   std_logic;
          DEBOUNCE_OUT_2        : out   std_logic;
          DRVR_EN               : out   std_logic;
          Data_FAIL             : out   std_logic;
          GPIO_11_M2F           : out   std_logic;
          GPIO_20_OUT           : out   std_logic;
          GPIO_21_M2F           : out   std_logic;
          GPIO_22_M2F           : out   std_logic;
          GPIO_24_M2F           : out   std_logic;
          GPIO_5_M2F            : out   std_logic;
          GPIO_8_M2F            : out   std_logic;
          MAC_MII_MDC           : out   std_logic;
          MAC_MII_TX_EN         : out   std_logic;
          MANCH_OUT_N           : out   std_logic;
          MANCH_OUT_P           : out   std_logic;
          MDDR_CAS_N            : out   std_logic;
          MDDR_CKE              : out   std_logic;
          MDDR_CLK              : out   std_logic;
          MDDR_CLK_N            : out   std_logic;
          MDDR_CS_N             : out   std_logic;
          MDDR_DQS_TMATCH_0_OUT : out   std_logic;
          MDDR_ODT              : out   std_logic;
          MDDR_RAS_N            : out   std_logic;
          MDDR_RESET_N          : out   std_logic;
          MDDR_WE_N             : out   std_logic;
          MMUART_0_TXD_M2F      : out   std_logic;
          MMUART_1_TXD          : out   std_logic;
          RCVR_EN               : out   std_logic;
          SPI_0_DO              : out   std_logic;
          SPI_0_SS1             : out   std_logic;
          SPI_1_DO_CAM          : out   std_logic;
          SPI_1_DO_OTH          : out   std_logic;
          GPIO_0_BI             : inout std_logic := 'Z';
          GPIO_12_BI            : inout std_logic := 'Z';
          GPIO_14_BI            : inout std_logic := 'Z';
          GPIO_15_BI            : inout std_logic := 'Z';
          GPIO_16_BI            : inout std_logic := 'Z';
          GPIO_17_BI            : inout std_logic := 'Z';
          GPIO_18_BI            : inout std_logic := 'Z';
          GPIO_25_BI            : inout std_logic := 'Z';
          GPIO_26_BI            : inout std_logic := 'Z';
          GPIO_31_BI            : inout std_logic := 'Z';
          GPIO_3_BI             : inout std_logic := 'Z';
          GPIO_4_BI             : inout std_logic := 'Z';
          I2C_1_SCL             : inout std_logic := 'Z';
          I2C_1_SDA             : inout std_logic := 'Z';
          MAC_MII_MDIO          : inout std_logic := 'Z';
          SPI_0_CLK             : inout std_logic := 'Z';
          SPI_0_SS0             : inout std_logic := 'Z';
          atck                  : in    std_logic;
          atdi                  : in    std_logic;
          atdo                  : out   std_logic;
          atms                  : in    std_logic;
          atrstb                : in    std_logic
        );

end m2s010_som;

architecture DEF_ARCH of m2s010_som is 

  component syn_identify_core0_0
    port( un6                              : in    std_logic_vector(5 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PRDATA     : in    std_logic_vector(7 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PADDR      : in    std_logic_vector(7 downto 0) := (others => 'U');
          clkdiv                           : in    std_logic_vector(3 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PWDATA     : in    std_logic_vector(7 downto 0) := (others => 'U');
          manches_in_dly                   : in    std_logic_vector(1 downto 0) := (others => 'U');
          iRX_FIFO_Full                    : in    std_logic_vector(3 downto 0) := (others => 'U');
          iRX_FIFO_Empty                   : in    std_logic_vector(3 downto 0) := (others => 'U');
          int_reg                          : in    std_logic_vector(7 downto 1) := (others => 'U');
          iRX_FIFO_UNDERRUN                : in    std_logic_vector(3 downto 0) := (others => 'U');
          ReadFIFO_Read_Ptr                : in    std_logic_vector(1 downto 0) := (others => 'U');
          packet_available_clear_reg       : in    std_logic_vector(2 downto 0) := (others => 'U');
          p2s_data                         : in    std_logic_vector(7 downto 0) := (others => 'U');
          RX_FIFO_DIN_pipe                 : in    std_logic_vector(8 downto 0) := (others => 'U');
          ReadFIFO_Write_Ptr               : in    std_logic_vector(1 downto 0) := (others => 'U');
          un15                             : in    std_logic_vector(10 downto 0) := (others => 'U');
          RX_FIFO_DOUT                     : in    std_logic_vector(8 downto 0) := (others => 'U');
          RX_packet_depth                  : in    std_logic_vector(7 downto 0) := (others => 'U');
          RX_FIFO_DIN                      : in    std_logic_vector(7 downto 0) := (others => 'U');
          up_EOP_del                       : in    std_logic_vector(5 downto 0) := (others => 'U');
          control_reg_0                    : in    std_logic := 'U';
          control_reg_2                    : in    std_logic := 'U';
          control_reg_3                    : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0              : in    std_logic := 'U';
          long_reset                       : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PREADY     : in    std_logic := 'U';
          block_int_until_rd               : in    std_logic := 'U';
          m2s010_som_sb_0_POWER_ON_RESET_N : in    std_logic := 'U';
          bd_reset                         : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PWRITE     : in    std_logic := 'U';
          iNRZ_data                        : in    std_logic := 'U';
          external_loopback                : in    std_logic := 'U';
          internal_loopback                : in    std_logic := 'U';
          start_tx_FIFO                    : in    std_logic := 'U';
          rx_FIFO_rst_reg                  : in    std_logic := 'U';
          TX_FIFO_RST                      : in    std_logic := 'U';
          irx_center_sample                : in    std_logic := 'U';
          int_reg_clr                      : in    std_logic := 'U';
          MANCHESTER_IN_c                  : in    std_logic := 'U';
          MANCH_OUT_P_c                    : in    std_logic := 'U';
          CommsFPGA_CCC_0_LOCK             : in    std_logic := 'U';
          TX_FIFO_Empty                    : in    std_logic := 'U';
          rx_packet_avail_int              : in    std_logic := 'U';
          rx_CRC_error_int                 : in    std_logic := 'U';
          RESET                            : in    std_logic := 'U';
          rx_packet_complt                 : in    std_logic := 'U';
          rx_FIFO_UNDERRUN_int             : in    std_logic := 'U';
          RX_FIFO_rd_en                    : in    std_logic := 'U';
          rx_FIFO_OVERFLOW_int             : in    std_logic := 'U';
          RX_FIFO_Full                     : in    std_logic := 'U';
          RX_FIFO_Empty                    : in    std_logic := 'U';
          RX_packet_depth_status           : in    std_logic := 'U';
          tx_packet_complt                 : in    std_logic := 'U';
          TX_FIFO_wr_en                    : in    std_logic := 'U';
          TX_FIFO_Full                     : in    std_logic := 'U';
          m2s010_som_sb_0_GPIO_28_SW_RESET : in    std_logic := 'U';
          iup_EOP                          : in    std_logic := 'U';
          atrstb                           : in    std_logic := 'U';
          atms                             : in    std_logic := 'U';
          atdo                             : out   std_logic;
          atdi                             : in    std_logic := 'U';
          atck                             : in    std_logic := 'U'
        );
  end component;

  component OUTBUF
    generic (IOSTD:string := "");

    port( D   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component INBUF
    generic (IOSTD:string := "");

    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component SLE
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          EN  : in    std_logic := 'U';
          ALn : in    std_logic := 'U';
          ADn : in    std_logic := 'U';
          SLn : in    std_logic := 'U';
          SD  : in    std_logic := 'U';
          LAT : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component CoreAPB3
    port( m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR : in    std_logic_vector(15 downto 12) := (others => 'U');
          CoreAPB3_0_APBmslave0_PSELx            : out   std_logic;
          m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx : in    std_logic := 'U'
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component m2s010_som_CommsFPGA_CCC_0_FCCC
    port( m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC : in    std_logic := 'U';
          CommsFPGA_CCC_0_LOCK                      : out   std_logic;
          CommsFPGA_CCC_0_GL1                       : out   std_logic;
          CommsFPGA_CCC_0_GL0                       : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component m2s010_som_ID_RES_0_IO
    port( ID_RES  : in    std_logic_vector(3 downto 0) := (others => 'U');
          Y_net_0 : out   std_logic_vector(3 downto 0)
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component m2s010_som_sb
    port( MDDR_DQS                                  : inout   std_logic_vector(1 downto 0);
          MDDR_DQ                                   : inout   std_logic_vector(15 downto 0);
          MDDR_DM_RDQS                              : inout   std_logic_vector(1 downto 0);
          MDDR_BA                                   : out   std_logic_vector(2 downto 0);
          MDDR_ADDR                                 : out   std_logic_vector(15 downto 0);
          CoreAPB3_0_APBmslave0_PADDR               : out   std_logic_vector(7 downto 0);
          m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR    : out   std_logic_vector(15 downto 12);
          CoreAPB3_0_APBmslave0_PWDATA              : out   std_logic_vector(7 downto 0);
          MAC_MII_TXD_c                             : out   std_logic_vector(3 downto 0);
          CoreAPB3_0_APBmslave0_PRDATA_m            : in    std_logic_vector(7 downto 0) := (others => 'U');
          Y_net_0                                   : in    std_logic_vector(3 downto 0) := (others => 'U');
          MAC_MII_RXD_c                             : in    std_logic_vector(3 downto 0) := (others => 'U');
          SPI_1_SS0_OTH_0                           : inout   std_logic;
          DEBOUNCE_OUT_net_0_0                      : in    std_logic := 'U';
          GPIO_7_PADI_0                             : inout   std_logic;
          GPIO_6_PAD_0                              : inout   std_logic;
          GPIO_1_BI_0                               : inout   std_logic;
          SPI_1_SS0_CAM_0                           : inout   std_logic;
          SPI_1_CLK_0                               : inout   std_logic;
          SPI_0_SS1                                 : out   std_logic;
          SPI_0_SS0                                 : inout   std_logic;
          SPI_0_DO                                  : out   std_logic;
          SPI_0_DI                                  : in    std_logic := 'U';
          SPI_0_CLK                                 : inout   std_logic;
          MMUART_1_TXD                              : out   std_logic;
          MMUART_1_RXD                              : in    std_logic := 'U';
          MDDR_WE_N                                 : out   std_logic;
          MDDR_RESET_N                              : out   std_logic;
          MDDR_RAS_N                                : out   std_logic;
          MDDR_ODT                                  : out   std_logic;
          MDDR_DQS_TMATCH_0_OUT                     : out   std_logic;
          MDDR_DQS_TMATCH_0_IN                      : in    std_logic := 'U';
          MDDR_CS_N                                 : out   std_logic;
          MDDR_CKE                                  : out   std_logic;
          MDDR_CAS_N                                : out   std_logic;
          I2C_1_SDA                                 : inout   std_logic;
          I2C_1_SCL                                 : inout   std_logic;
          GPIO_31_BI                                : inout   std_logic;
          GPIO_26_BI                                : inout   std_logic;
          GPIO_25_BI                                : inout   std_logic;
          GPIO_20_OUT                               : out   std_logic;
          GPIO_18_BI                                : inout   std_logic;
          GPIO_17_BI                                : inout   std_logic;
          GPIO_16_BI                                : inout   std_logic;
          GPIO_15_BI                                : inout   std_logic;
          GPIO_14_BI                                : inout   std_logic;
          GPIO_12_BI                                : inout   std_logic;
          GPIO_4_BI                                 : inout   std_logic;
          GPIO_3_BI                                 : inout   std_logic;
          GPIO_0_BI                                 : inout   std_logic;
          CoreAPB3_0_APBmslave0_PENABLE             : out   std_logic;
          m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx    : out   std_logic;
          CoreAPB3_0_APBmslave0_PWRITE              : out   std_logic;
          MAC_MII_MDC_c                             : out   std_logic;
          GPIO_22_M2F_c                             : out   std_logic;
          GPIO_21_M2F_c                             : out   std_logic;
          m2s010_som_sb_0_GPIO_28_SW_RESET          : out   std_logic;
          MMUART_0_TXD_M2F_c                        : out   std_logic;
          GPIO_24_M2F_c                             : out   std_logic;
          GPIO_5_M2F_c                              : out   std_logic;
          GPIO_8_M2F_c                              : out   std_logic;
          GPIO_11_M2F_c                             : out   std_logic;
          MAC_MII_TX_EN_c                           : out   std_logic;
          MAC_MII_COL_c                             : in    std_logic := 'U';
          MAC_MII_CRS_c                             : in    std_logic := 'U';
          CommsFPGA_top_0_INT                       : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PREADY_i_m_i        : in    std_logic := 'U';
          DEBOUNCE_OUT_1_c                          : in    std_logic := 'U';
          DEBOUNCE_OUT_2_c                          : in    std_logic := 'U';
          MMUART_0_RXD_F2M_c                        : in    std_logic := 'U';
          MAC_MII_RX_CLK_c                          : in    std_logic := 'U';
          MAC_MII_RX_DV_c                           : in    std_logic := 'U';
          MAC_MII_RX_ER_c                           : in    std_logic := 'U';
          MAC_MII_TX_CLK_c                          : in    std_logic := 'U';
          MDDR_CLK_N                                : out   std_logic;
          MDDR_CLK                                  : out   std_logic;
          XTL                                       : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz                 : out   std_logic;
          m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC : inout   std_logic;
          SPI_1_DI_CAM_c                            : in    std_logic := 'U';
          SPI_1_DI_OTH_c                            : in    std_logic := 'U';
          CommsFPGA_top_0_CAMERA_NODE               : in    std_logic := 'U';
          DEVRST_N                                  : in    std_logic := 'U';
          m2s010_som_sb_0_POWER_ON_RESET_N          : out   std_logic;
          MAC_MII_MDIO                              : inout   std_logic;
          SPI_1_DO_CAM_c                            : inout   std_logic;
          SPI_1_DO_OTH                              : out   std_logic
        );
  end component;

  component CommsFPGA_top
    port( packet_available_clear_reg         : out   std_logic_vector(2 downto 0);
          ReadFIFO_Read_Ptr                  : out   std_logic_vector(1 downto 0);
          ReadFIFO_Write_Ptr                 : out   std_logic_vector(1 downto 0);
          iRX_FIFO_Empty                     : out   std_logic_vector(3 downto 0);
          iRX_FIFO_UNDERRUN                  : out   std_logic_vector(3 downto 0);
          iRX_FIFO_Full                      : out   std_logic_vector(3 downto 0);
          CoreAPB3_0_APBmslave0_PRDATA_m     : out   std_logic_vector(7 downto 0);
          un15                               : out   std_logic_vector(10 downto 0);
          RX_FIFO_DIN                        : out   std_logic_vector(7 downto 0);
          RX_FIFO_DIN_pipe                   : out   std_logic_vector(8 downto 0);
          clkdiv                             : out   std_logic_vector(3 downto 0);
          un6                                : out   std_logic_vector(5 downto 0);
          p2s_data                           : out   std_logic_vector(7 downto 0);
          manches_in_dly                     : out   std_logic_vector(1 downto 0);
          CoreAPB3_0_APBmslave0_PWDATA       : in    std_logic_vector(7 downto 0) := (others => 'U');
          CoreAPB3_0_APBmslave0_PRDATA       : out   std_logic_vector(7 downto 0);
          RX_packet_depth                    : out   std_logic_vector(7 downto 0);
          CoreAPB3_0_APBmslave0_PADDR        : in    std_logic_vector(7 downto 0) := (others => 'U');
          RX_FIFO_DOUT                       : out   std_logic_vector(8 downto 0);
          int_reg                            : out   std_logic_vector(7 downto 1);
          up_EOP_del                         : out   std_logic_vector(5 downto 0);
          DEBOUNCE_IN_c                      : in    std_logic_vector(2 downto 0) := (others => 'U');
          Y_net_0                            : in    std_logic_vector(3 downto 1) := (others => 'U');
          control_reg_0                      : out   std_logic;
          control_reg_2                      : out   std_logic;
          control_reg_3                      : out   std_logic;
          DEBOUNCE_OUT_net_0_0               : out   std_logic;
          CoreAPB3_0_APBmslave0_PREADY_i_m_i : out   std_logic;
          MANCHESTER_IN_c                    : in    std_logic := 'U';
          irx_center_sample                  : out   std_logic;
          iNRZ_data                          : out   std_logic;
          MANCH_OUT_P_c                      : out   std_logic;
          MANCH_OUT_P_c_i                    : out   std_logic;
          DRVR_EN_c                          : out   std_logic;
          iup_EOP                            : out   std_logic;
          long_reset_set                     : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PREADY       : out   std_logic;
          external_loopback                  : out   std_logic;
          internal_loopback                  : out   std_logic;
          start_tx_FIFO                      : out   std_logic;
          TX_FIFO_RST                        : out   std_logic;
          N_480_i_i                          : in    std_logic := 'U';
          RX_FIFO_rd_en                      : out   std_logic;
          TX_FIFO_wr_en                      : out   std_logic;
          RX_packet_depth_status             : out   std_logic;
          rx_packet_complt                   : out   std_logic;
          rx_packet_avail_int                : out   std_logic;
          TX_FIFO_Full                       : out   std_logic;
          TX_FIFO_Empty                      : out   std_logic;
          CoreAPB3_0_APBmslave0_PSELx        : in    std_logic := 'U';
          CoreAPB3_0_APBmslave0_PENABLE      : in    std_logic := 'U';
          RX_FIFO_Full                       : out   std_logic;
          RX_FIFO_Empty                      : out   std_logic;
          CoreAPB3_0_APBmslave0_PWRITE       : in    std_logic := 'U';
          N_480_i                            : out   std_logic;
          CommsFPGA_top_0_INT                : out   std_logic;
          int_reg_clr                        : out   std_logic;
          rx_FIFO_UNDERRUN_int               : out   std_logic;
          rx_FIFO_OVERFLOW_int               : out   std_logic;
          rx_CRC_error_int                   : out   std_logic;
          tx_packet_complt                   : out   std_logic;
          block_int_until_rd                 : out   std_logic;
          RESET_set                          : in    std_logic := 'U';
          DEBOUNCE_OUT_1_c                   : out   std_logic;
          DEBOUNCE_OUT_2_c                   : out   std_logic;
          CommsFPGA_top_0_CAMERA_NODE        : out   std_logic;
          CommsFPGA_CCC_0_LOCK               : in    std_logic := 'U';
          m2s010_som_sb_0_POWER_ON_RESET_N   : in    std_logic := 'U';
          m2s010_som_sb_0_GPIO_28_SW_RESET   : in    std_logic := 'U';
          rx_FIFO_rst_reg                    : out   std_logic;
          CommsFPGA_CCC_0_GL1                : in    std_logic := 'U';
          CommsFPGA_CCC_0_GL0                : in    std_logic := 'U';
          m2s010_som_sb_0_CCC_71MHz          : in    std_logic := 'U';
          long_reset_i                       : out   std_logic;
          RESET_i                            : out   std_logic;
          RESET                              : out   std_logic;
          BIT_CLK                            : out   std_logic;
          long_reset                         : out   std_logic;
          bd_reset                           : out   std_logic
        );
  end component;

    signal m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC, 
        CommsFPGA_CCC_0_LOCK, CommsFPGA_CCC_0_GL0, 
        CommsFPGA_CCC_0_GL1, m2s010_som_sb_0_GPIO_28_SW_RESET, 
        m2s010_som_sb_0_POWER_ON_RESET_N, 
        m2s010_som_sb_0_CCC_71MHz, 
        \CoreAPB3_0_APBmslave0_PRDATA[0]\, 
        \CoreAPB3_0_APBmslave0_PRDATA[1]\, 
        \CoreAPB3_0_APBmslave0_PRDATA[2]\, 
        \CoreAPB3_0_APBmslave0_PRDATA[3]\, 
        \CoreAPB3_0_APBmslave0_PRDATA[4]\, 
        \CoreAPB3_0_APBmslave0_PRDATA[5]\, 
        \CoreAPB3_0_APBmslave0_PRDATA[6]\, 
        \CoreAPB3_0_APBmslave0_PRDATA[7]\, 
        CoreAPB3_0_APBmslave0_PREADY, \Y_net_0[0]\, \Y_net_0[1]\, 
        \Y_net_0[2]\, \Y_net_0[3]\, CommsFPGA_top_0_CAMERA_NODE, 
        CommsFPGA_top_0_INT, \DEBOUNCE_OUT_net_0[0]\, GND_net_1, 
        \CoreAPB3_0_APBmslave0_PADDR[0]\, 
        \CoreAPB3_0_APBmslave0_PADDR[1]\, 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, 
        \CoreAPB3_0_APBmslave0_PADDR[4]\, 
        \CoreAPB3_0_APBmslave0_PADDR[5]\, 
        \CoreAPB3_0_APBmslave0_PADDR[6]\, 
        \CoreAPB3_0_APBmslave0_PADDR[7]\, 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[12]\, 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[13]\, 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[14]\, 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[15]\, 
        CoreAPB3_0_APBmslave0_PWRITE, 
        CoreAPB3_0_APBmslave0_PENABLE, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx, 
        \CoreAPB3_0_APBmslave0_PWDATA[0]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[1]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[2]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[3]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[4]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[5]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[6]\, 
        \CoreAPB3_0_APBmslave0_PWDATA[7]\, VCC_net_1, 
        \RX_FIFO_DIN_pipe[0]\, \RX_FIFO_DIN_pipe[1]\, 
        \RX_FIFO_DIN_pipe[2]\, \RX_FIFO_DIN_pipe[3]\, 
        \RX_FIFO_DIN_pipe[4]\, \RX_FIFO_DIN_pipe[5]\, 
        \RX_FIFO_DIN_pipe[6]\, \RX_FIFO_DIN_pipe[7]\, 
        \RX_FIFO_DIN_pipe[8]\, RESET, bd_reset, tx_packet_complt, 
        TX_FIFO_wr_en, TX_FIFO_Full, TX_FIFO_Empty, RX_FIFO_rd_en, 
        RX_FIFO_Full, RX_FIFO_Empty, \RX_FIFO_DOUT[0]\, 
        \RX_FIFO_DOUT[1]\, \RX_FIFO_DOUT[2]\, \RX_FIFO_DOUT[3]\, 
        \RX_FIFO_DOUT[4]\, \RX_FIFO_DOUT[5]\, \RX_FIFO_DOUT[6]\, 
        \RX_FIFO_DOUT[7]\, \RX_FIFO_DOUT[8]\, iup_EOP, 
        RX_packet_depth_status, \RX_packet_depth[0]\, 
        \RX_packet_depth[1]\, \RX_packet_depth[2]\, 
        \RX_packet_depth[3]\, \RX_packet_depth[4]\, 
        \RX_packet_depth[5]\, \RX_packet_depth[6]\, 
        \RX_packet_depth[7]\, \int_reg[1]\, \int_reg[2]\, 
        \int_reg[3]\, \int_reg[4]\, \int_reg[5]\, \int_reg[6]\, 
        \int_reg[7]\, \control_reg[0]\, external_loopback, 
        \control_reg[2]\, \control_reg[3]\, internal_loopback, 
        start_tx_FIFO, rx_FIFO_rst_reg, TX_FIFO_RST, 
        \up_EOP_del[0]\, \up_EOP_del[1]\, \up_EOP_del[2]\, 
        \up_EOP_del[3]\, \up_EOP_del[4]\, \up_EOP_del[5]\, 
        rx_FIFO_UNDERRUN_int, rx_FIFO_OVERFLOW_int, 
        rx_CRC_error_int, rx_packet_avail_int, int_reg_clr, 
        block_int_until_rd, long_reset, \p2s_data[0]\, 
        \p2s_data[1]\, \p2s_data[2]\, \p2s_data[3]\, 
        \p2s_data[4]\, \p2s_data[5]\, \p2s_data[6]\, 
        \p2s_data[7]\, \un15[10]\, \un15[5]\, \un15[4]\, 
        \un15[3]\, \un15[2]\, \un15[1]\, \un15[0]\, 
        \RX_FIFO_DIN[0]\, \RX_FIFO_DIN[1]\, \RX_FIFO_DIN[2]\, 
        \RX_FIFO_DIN[3]\, \RX_FIFO_DIN[4]\, \RX_FIFO_DIN[5]\, 
        \RX_FIFO_DIN[6]\, \RX_FIFO_DIN[7]\, irx_center_sample, 
        iNRZ_data, \manches_in_dly[0]\, \manches_in_dly[1]\, 
        \clkdiv[0]\, \clkdiv[1]\, \clkdiv[2]\, \clkdiv[3]\, 
        \un6[5]\, \un6[4]\, \un6[3]\, \un6[2]\, \un6[0]\, 
        \ReadFIFO_Write_Ptr[0]\, \ReadFIFO_Write_Ptr[1]\, 
        \packet_available_clear_reg[0]\, 
        \packet_available_clear_reg[1]\, 
        \packet_available_clear_reg[2]\, \iRX_FIFO_UNDERRUN[0]\, 
        \iRX_FIFO_UNDERRUN[1]\, \iRX_FIFO_UNDERRUN[2]\, 
        \iRX_FIFO_UNDERRUN[3]\, \iRX_FIFO_Full[0]\, 
        \iRX_FIFO_Full[1]\, \iRX_FIFO_Full[2]\, 
        \iRX_FIFO_Full[3]\, \iRX_FIFO_Empty[0]\, 
        \iRX_FIFO_Empty[1]\, \iRX_FIFO_Empty[2]\, 
        \iRX_FIFO_Empty[3]\, \CoreAPB3_0_APBmslave0_PRDATA_m[0]\, 
        \CoreAPB3_0_APBmslave0_PRDATA_m[1]\, 
        \CoreAPB3_0_APBmslave0_PRDATA_m[2]\, 
        \CoreAPB3_0_APBmslave0_PRDATA_m[3]\, 
        \CoreAPB3_0_APBmslave0_PRDATA_m[4]\, 
        \CoreAPB3_0_APBmslave0_PRDATA_m[5]\, 
        \CoreAPB3_0_APBmslave0_PRDATA_m[6]\, 
        \CoreAPB3_0_APBmslave0_PRDATA_m[7]\, 
        CoreAPB3_0_APBmslave0_PSELx, \CommsFPGA_top_0.BIT_CLK\, 
        \un15[9]\, \un15[7]\, \un15[8]\, \ReadFIFO_Read_Ptr[1]\, 
        \ReadFIFO_Read_Ptr[0]\, \DEBOUNCE_IN_c[0]\, 
        \DEBOUNCE_IN_c[1]\, \DEBOUNCE_IN_c[2]\, MAC_MII_COL_c, 
        MAC_MII_CRS_c, \MAC_MII_RXD_c[0]\, \MAC_MII_RXD_c[1]\, 
        \MAC_MII_RXD_c[2]\, \MAC_MII_RXD_c[3]\, MAC_MII_RX_CLK_c, 
        MAC_MII_RX_DV_c, MAC_MII_RX_ER_c, MAC_MII_TX_CLK_c, 
        MANCHESTER_IN_c, MMUART_0_RXD_F2M_c, Data_FAIL_c, 
        SPI_1_DI_CAM_c, SPI_1_DI_OTH_c, DEBOUNCE_OUT_1_c, 
        DEBOUNCE_OUT_2_c, DRVR_EN_c, GPIO_11_M2F_c, GPIO_21_M2F_c, 
        GPIO_22_M2F_c, GPIO_24_M2F_c, GPIO_5_M2F_c, GPIO_8_M2F_c, 
        MAC_MII_MDC_c, \MAC_MII_TXD_c[0]\, \MAC_MII_TXD_c[1]\, 
        \MAC_MII_TXD_c[2]\, \MAC_MII_TXD_c[3]\, MAC_MII_TX_EN_c, 
        MANCH_OUT_P_c, MMUART_0_TXD_M2F_c, SPI_1_DO_CAM_c, 
        rx_packet_complt, MANCH_OUT_P_c_i, 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i, 
        \CommsFPGA_top_0.N_480_i_i\, RESET_i, long_reset_i, 
        \long_reset_set\, \RESET_set\, N_480_i : std_logic;
    signal nc2, nc4, nc3, nc1 : std_logic;

    for all : syn_identify_core0_0
	Use entity work.syn_identify_core0_0(DEF_ARCH);
    for all : CoreAPB3
	Use entity work.CoreAPB3(DEF_ARCH);
    for all : m2s010_som_CommsFPGA_CCC_0_FCCC
	Use entity work.m2s010_som_CommsFPGA_CCC_0_FCCC(DEF_ARCH);
    for all : m2s010_som_ID_RES_0_IO
	Use entity work.m2s010_som_ID_RES_0_IO(DEF_ARCH);
    for all : m2s010_som_sb
	Use entity work.m2s010_som_sb(DEF_ARCH);
    for all : CommsFPGA_top
	Use entity work.CommsFPGA_top(DEF_ARCH);
begin 


    ident_coreinst : syn_identify_core0_0
      port map(un6(5) => \un6[5]\, un6(4) => \un6[4]\, un6(3) => 
        \un6[3]\, un6(2) => \un6[2]\, un6(1) => nc2, un6(0) => 
        \un6[0]\, CoreAPB3_0_APBmslave0_PRDATA(7) => 
        \CoreAPB3_0_APBmslave0_PRDATA[7]\, 
        CoreAPB3_0_APBmslave0_PRDATA(6) => 
        \CoreAPB3_0_APBmslave0_PRDATA[6]\, 
        CoreAPB3_0_APBmslave0_PRDATA(5) => 
        \CoreAPB3_0_APBmslave0_PRDATA[5]\, 
        CoreAPB3_0_APBmslave0_PRDATA(4) => 
        \CoreAPB3_0_APBmslave0_PRDATA[4]\, 
        CoreAPB3_0_APBmslave0_PRDATA(3) => 
        \CoreAPB3_0_APBmslave0_PRDATA[3]\, 
        CoreAPB3_0_APBmslave0_PRDATA(2) => 
        \CoreAPB3_0_APBmslave0_PRDATA[2]\, 
        CoreAPB3_0_APBmslave0_PRDATA(1) => 
        \CoreAPB3_0_APBmslave0_PRDATA[1]\, 
        CoreAPB3_0_APBmslave0_PRDATA(0) => 
        \CoreAPB3_0_APBmslave0_PRDATA[0]\, 
        CoreAPB3_0_APBmslave0_PADDR(7) => 
        \CoreAPB3_0_APBmslave0_PADDR[7]\, 
        CoreAPB3_0_APBmslave0_PADDR(6) => 
        \CoreAPB3_0_APBmslave0_PADDR[6]\, 
        CoreAPB3_0_APBmslave0_PADDR(5) => 
        \CoreAPB3_0_APBmslave0_PADDR[5]\, 
        CoreAPB3_0_APBmslave0_PADDR(4) => 
        \CoreAPB3_0_APBmslave0_PADDR[4]\, 
        CoreAPB3_0_APBmslave0_PADDR(3) => 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, 
        CoreAPB3_0_APBmslave0_PADDR(1) => 
        \CoreAPB3_0_APBmslave0_PADDR[1]\, 
        CoreAPB3_0_APBmslave0_PADDR(0) => 
        \CoreAPB3_0_APBmslave0_PADDR[0]\, clkdiv(3) => 
        \clkdiv[3]\, clkdiv(2) => \clkdiv[2]\, clkdiv(1) => 
        \clkdiv[1]\, clkdiv(0) => \clkdiv[0]\, 
        CoreAPB3_0_APBmslave0_PWDATA(7) => 
        \CoreAPB3_0_APBmslave0_PWDATA[7]\, 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        \CoreAPB3_0_APBmslave0_PWDATA[6]\, 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        \CoreAPB3_0_APBmslave0_PWDATA[5]\, 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        \CoreAPB3_0_APBmslave0_PWDATA[4]\, 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        \CoreAPB3_0_APBmslave0_PWDATA[3]\, 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        \CoreAPB3_0_APBmslave0_PWDATA[2]\, 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        \CoreAPB3_0_APBmslave0_PWDATA[1]\, 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        \CoreAPB3_0_APBmslave0_PWDATA[0]\, manches_in_dly(1) => 
        \manches_in_dly[1]\, manches_in_dly(0) => 
        \manches_in_dly[0]\, iRX_FIFO_Full(3) => 
        \iRX_FIFO_Full[3]\, iRX_FIFO_Full(2) => 
        \iRX_FIFO_Full[2]\, iRX_FIFO_Full(1) => 
        \iRX_FIFO_Full[1]\, iRX_FIFO_Full(0) => 
        \iRX_FIFO_Full[0]\, iRX_FIFO_Empty(3) => 
        \iRX_FIFO_Empty[3]\, iRX_FIFO_Empty(2) => 
        \iRX_FIFO_Empty[2]\, iRX_FIFO_Empty(1) => 
        \iRX_FIFO_Empty[1]\, iRX_FIFO_Empty(0) => 
        \iRX_FIFO_Empty[0]\, int_reg(7) => \int_reg[7]\, 
        int_reg(6) => \int_reg[6]\, int_reg(5) => \int_reg[5]\, 
        int_reg(4) => \int_reg[4]\, int_reg(3) => \int_reg[3]\, 
        int_reg(2) => \int_reg[2]\, int_reg(1) => \int_reg[1]\, 
        iRX_FIFO_UNDERRUN(3) => \iRX_FIFO_UNDERRUN[3]\, 
        iRX_FIFO_UNDERRUN(2) => \iRX_FIFO_UNDERRUN[2]\, 
        iRX_FIFO_UNDERRUN(1) => \iRX_FIFO_UNDERRUN[1]\, 
        iRX_FIFO_UNDERRUN(0) => \iRX_FIFO_UNDERRUN[0]\, 
        ReadFIFO_Read_Ptr(1) => \ReadFIFO_Read_Ptr[1]\, 
        ReadFIFO_Read_Ptr(0) => \ReadFIFO_Read_Ptr[0]\, 
        packet_available_clear_reg(2) => 
        \packet_available_clear_reg[2]\, 
        packet_available_clear_reg(1) => 
        \packet_available_clear_reg[1]\, 
        packet_available_clear_reg(0) => 
        \packet_available_clear_reg[0]\, p2s_data(7) => 
        \p2s_data[7]\, p2s_data(6) => \p2s_data[6]\, p2s_data(5)
         => \p2s_data[5]\, p2s_data(4) => \p2s_data[4]\, 
        p2s_data(3) => \p2s_data[3]\, p2s_data(2) => 
        \p2s_data[2]\, p2s_data(1) => \p2s_data[1]\, p2s_data(0)
         => \p2s_data[0]\, RX_FIFO_DIN_pipe(8) => 
        \RX_FIFO_DIN_pipe[8]\, RX_FIFO_DIN_pipe(7) => 
        \RX_FIFO_DIN_pipe[7]\, RX_FIFO_DIN_pipe(6) => 
        \RX_FIFO_DIN_pipe[6]\, RX_FIFO_DIN_pipe(5) => 
        \RX_FIFO_DIN_pipe[5]\, RX_FIFO_DIN_pipe(4) => 
        \RX_FIFO_DIN_pipe[4]\, RX_FIFO_DIN_pipe(3) => 
        \RX_FIFO_DIN_pipe[3]\, RX_FIFO_DIN_pipe(2) => 
        \RX_FIFO_DIN_pipe[2]\, RX_FIFO_DIN_pipe(1) => 
        \RX_FIFO_DIN_pipe[1]\, RX_FIFO_DIN_pipe(0) => 
        \RX_FIFO_DIN_pipe[0]\, ReadFIFO_Write_Ptr(1) => 
        \ReadFIFO_Write_Ptr[1]\, ReadFIFO_Write_Ptr(0) => 
        \ReadFIFO_Write_Ptr[0]\, un15(10) => \un15[10]\, un15(9)
         => \un15[9]\, un15(8) => \un15[8]\, un15(7) => \un15[7]\, 
        un15(6) => nc4, un15(5) => \un15[5]\, un15(4) => 
        \un15[4]\, un15(3) => \un15[3]\, un15(2) => \un15[2]\, 
        un15(1) => \un15[1]\, un15(0) => \un15[0]\, 
        RX_FIFO_DOUT(8) => \RX_FIFO_DOUT[8]\, RX_FIFO_DOUT(7) => 
        \RX_FIFO_DOUT[7]\, RX_FIFO_DOUT(6) => \RX_FIFO_DOUT[6]\, 
        RX_FIFO_DOUT(5) => \RX_FIFO_DOUT[5]\, RX_FIFO_DOUT(4) => 
        \RX_FIFO_DOUT[4]\, RX_FIFO_DOUT(3) => \RX_FIFO_DOUT[3]\, 
        RX_FIFO_DOUT(2) => \RX_FIFO_DOUT[2]\, RX_FIFO_DOUT(1) => 
        \RX_FIFO_DOUT[1]\, RX_FIFO_DOUT(0) => \RX_FIFO_DOUT[0]\, 
        RX_packet_depth(7) => \RX_packet_depth[7]\, 
        RX_packet_depth(6) => \RX_packet_depth[6]\, 
        RX_packet_depth(5) => \RX_packet_depth[5]\, 
        RX_packet_depth(4) => \RX_packet_depth[4]\, 
        RX_packet_depth(3) => \RX_packet_depth[3]\, 
        RX_packet_depth(2) => \RX_packet_depth[2]\, 
        RX_packet_depth(1) => \RX_packet_depth[1]\, 
        RX_packet_depth(0) => \RX_packet_depth[0]\, 
        RX_FIFO_DIN(7) => \RX_FIFO_DIN[7]\, RX_FIFO_DIN(6) => 
        \RX_FIFO_DIN[6]\, RX_FIFO_DIN(5) => \RX_FIFO_DIN[5]\, 
        RX_FIFO_DIN(4) => \RX_FIFO_DIN[4]\, RX_FIFO_DIN(3) => 
        \RX_FIFO_DIN[3]\, RX_FIFO_DIN(2) => \RX_FIFO_DIN[2]\, 
        RX_FIFO_DIN(1) => \RX_FIFO_DIN[1]\, RX_FIFO_DIN(0) => 
        \RX_FIFO_DIN[0]\, up_EOP_del(5) => \up_EOP_del[5]\, 
        up_EOP_del(4) => \up_EOP_del[4]\, up_EOP_del(3) => 
        \up_EOP_del[3]\, up_EOP_del(2) => \up_EOP_del[2]\, 
        up_EOP_del(1) => \up_EOP_del[1]\, up_EOP_del(0) => 
        \up_EOP_del[0]\, control_reg_0 => \control_reg[0]\, 
        control_reg_2 => \control_reg[2]\, control_reg_3 => 
        \control_reg[3]\, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, long_reset => long_reset, 
        CoreAPB3_0_APBmslave0_PREADY => 
        CoreAPB3_0_APBmslave0_PREADY, block_int_until_rd => 
        block_int_until_rd, m2s010_som_sb_0_POWER_ON_RESET_N => 
        m2s010_som_sb_0_POWER_ON_RESET_N, bd_reset => bd_reset, 
        CoreAPB3_0_APBmslave0_PWRITE => 
        CoreAPB3_0_APBmslave0_PWRITE, iNRZ_data => iNRZ_data, 
        external_loopback => external_loopback, internal_loopback
         => internal_loopback, start_tx_FIFO => start_tx_FIFO, 
        rx_FIFO_rst_reg => rx_FIFO_rst_reg, TX_FIFO_RST => 
        TX_FIFO_RST, irx_center_sample => irx_center_sample, 
        int_reg_clr => int_reg_clr, MANCHESTER_IN_c => 
        MANCHESTER_IN_c, MANCH_OUT_P_c => MANCH_OUT_P_c, 
        CommsFPGA_CCC_0_LOCK => CommsFPGA_CCC_0_LOCK, 
        TX_FIFO_Empty => TX_FIFO_Empty, rx_packet_avail_int => 
        rx_packet_avail_int, rx_CRC_error_int => rx_CRC_error_int, 
        RESET => RESET, rx_packet_complt => rx_packet_complt, 
        rx_FIFO_UNDERRUN_int => rx_FIFO_UNDERRUN_int, 
        RX_FIFO_rd_en => RX_FIFO_rd_en, rx_FIFO_OVERFLOW_int => 
        rx_FIFO_OVERFLOW_int, RX_FIFO_Full => RX_FIFO_Full, 
        RX_FIFO_Empty => RX_FIFO_Empty, RX_packet_depth_status
         => RX_packet_depth_status, tx_packet_complt => 
        tx_packet_complt, TX_FIFO_wr_en => TX_FIFO_wr_en, 
        TX_FIFO_Full => TX_FIFO_Full, 
        m2s010_som_sb_0_GPIO_28_SW_RESET => 
        m2s010_som_sb_0_GPIO_28_SW_RESET, iup_EOP => iup_EOP, 
        atrstb => atrstb, atms => atms, atdo => atdo, atdi => 
        atdi, atck => atck);
    
    RCVR_EN_obuf : OUTBUF
      port map(D => VCC_net_1, PAD => RCVR_EN);
    
    MANCH_OUT_N_obuf : OUTBUF
      port map(D => MANCH_OUT_P_c_i, PAD => MANCH_OUT_N);
    
    \MAC_MII_RXD_ibuf[1]\ : INBUF
      port map(PAD => MAC_MII_RXD(1), Y => \MAC_MII_RXD_c[1]\);
    
    long_reset_set : SLE
      port map(D => GND_net_1, CLK => m2s010_som_sb_0_CCC_71MHz, 
        EN => VCC_net_1, ALn => long_reset_i, ADn => GND_net_1, 
        SLn => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q
         => \long_reset_set\);
    
    MMUART_0_RXD_F2M_ibuf : INBUF
      port map(PAD => MMUART_0_RXD_F2M, Y => MMUART_0_RXD_F2M_c);
    
    MAC_MII_RX_CLK_ibuf : INBUF
      port map(PAD => MAC_MII_RX_CLK, Y => MAC_MII_RX_CLK_c);
    
    MAC_MII_CRS_ibuf : INBUF
      port map(PAD => MAC_MII_CRS, Y => MAC_MII_CRS_c);
    
    CoreAPB3_0 : CoreAPB3
      port map(m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(15) => 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[15]\, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(14) => 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[14]\, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(13) => 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[13]\, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(12) => 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[12]\, 
        CoreAPB3_0_APBmslave0_PSELx => 
        CoreAPB3_0_APBmslave0_PSELx, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx);
    
    \VCC\ : VCC
      port map(Y => VCC_net_1);
    
    CommsFPGA_CCC_0 : m2s010_som_CommsFPGA_CCC_0_FCCC
      port map(m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC => 
        m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC, 
        CommsFPGA_CCC_0_LOCK => CommsFPGA_CCC_0_LOCK, 
        CommsFPGA_CCC_0_GL1 => CommsFPGA_CCC_0_GL1, 
        CommsFPGA_CCC_0_GL0 => CommsFPGA_CCC_0_GL0);
    
    MAC_MII_TX_EN_obuf : OUTBUF
      port map(D => MAC_MII_TX_EN_c, PAD => MAC_MII_TX_EN);
    
    MAC_MII_TX_CLK_ibuf : INBUF
      port map(PAD => MAC_MII_TX_CLK, Y => MAC_MII_TX_CLK_c);
    
    I_940 : CLKINT
      port map(A => N_480_i, Y => \CommsFPGA_top_0.N_480_i_i\);
    
    \MAC_MII_TXD_obuf[1]\ : OUTBUF
      port map(D => \MAC_MII_TXD_c[1]\, PAD => MAC_MII_TXD(1));
    
    DEBOUNCE_OUT_2_obuf : OUTBUF
      port map(D => DEBOUNCE_OUT_2_c, PAD => DEBOUNCE_OUT_2);
    
    ID_RES_0 : m2s010_som_ID_RES_0_IO
      port map(ID_RES(3) => ID_RES(3), ID_RES(2) => ID_RES(2), 
        ID_RES(1) => ID_RES(1), ID_RES(0) => ID_RES(0), 
        Y_net_0(3) => \Y_net_0[3]\, Y_net_0(2) => \Y_net_0[2]\, 
        Y_net_0(1) => \Y_net_0[1]\, Y_net_0(0) => \Y_net_0[0]\);
    
    \MAC_MII_RXD_ibuf[0]\ : INBUF
      port map(PAD => MAC_MII_RXD(0), Y => \MAC_MII_RXD_c[0]\);
    
    MMUART_0_TXD_M2F_obuf : OUTBUF
      port map(D => MMUART_0_TXD_M2F_c, PAD => MMUART_0_TXD_M2F);
    
    \GND\ : GND
      port map(Y => GND_net_1);
    
    \MAC_MII_RXD_ibuf[3]\ : INBUF
      port map(PAD => MAC_MII_RXD(3), Y => \MAC_MII_RXD_c[3]\);
    
    SPI_1_DI_CAM_ibuf : INBUF
      port map(PAD => SPI_1_DI_CAM, Y => SPI_1_DI_CAM_c);
    
    \MAC_MII_TXD_obuf[0]\ : OUTBUF
      port map(D => \MAC_MII_TXD_c[0]\, PAD => MAC_MII_TXD(0));
    
    Data_FAIL_obuf : OUTBUF
      port map(D => Data_FAIL_c, PAD => Data_FAIL);
    
    MAC_MII_COL_ibuf : INBUF
      port map(PAD => MAC_MII_COL, Y => MAC_MII_COL_c);
    
    MANCH_OUT_P_obuf : OUTBUF
      port map(D => MANCH_OUT_P_c, PAD => MANCH_OUT_P);
    
    MAC_MII_MDC_obuf : OUTBUF
      port map(D => MAC_MII_MDC_c, PAD => MAC_MII_MDC);
    
    MANCHESTER_IN_ibuf : INBUF
      port map(PAD => MANCHESTER_IN, Y => MANCHESTER_IN_c);
    
    GPIO_22_M2F_obuf : OUTBUF
      port map(D => GPIO_22_M2F_c, PAD => GPIO_22_M2F);
    
    GPIO_21_M2F_obuf : OUTBUF
      port map(D => GPIO_21_M2F_c, PAD => GPIO_21_M2F);
    
    SPI_1_DO_CAM_obuf : OUTBUF
      port map(D => SPI_1_DO_CAM_c, PAD => SPI_1_DO_CAM);
    
    \MAC_MII_TXD_obuf[3]\ : OUTBUF
      port map(D => \MAC_MII_TXD_c[3]\, PAD => MAC_MII_TXD(3));
    
    \DEBOUNCE_IN_ibuf[1]\ : INBUF
      port map(PAD => DEBOUNCE_IN(1), Y => \DEBOUNCE_IN_c[1]\);
    
    MAC_MII_RX_DV_ibuf : INBUF
      port map(PAD => MAC_MII_RX_DV, Y => MAC_MII_RX_DV_c);
    
    DRVR_EN_obuf : OUTBUF
      port map(D => DRVR_EN_c, PAD => DRVR_EN);
    
    DEBOUNCE_OUT_1_obuf : OUTBUF
      port map(D => DEBOUNCE_OUT_1_c, PAD => DEBOUNCE_OUT_1);
    
    RESET_set : SLE
      port map(D => GND_net_1, CLK => \CommsFPGA_top_0.BIT_CLK\, 
        EN => VCC_net_1, ALn => RESET_i, ADn => GND_net_1, SLn
         => VCC_net_1, SD => GND_net_1, LAT => GND_net_1, Q => 
        \RESET_set\);
    
    SPI_1_DI_OTH_ibuf : INBUF
      port map(PAD => SPI_1_DI_OTH, Y => SPI_1_DI_OTH_c);
    
    m2s010_som_sb_0 : m2s010_som_sb
      port map(MDDR_DQS(1) => MDDR_DQS(1), MDDR_DQS(0) => 
        MDDR_DQS(0), MDDR_DQ(15) => MDDR_DQ(15), MDDR_DQ(14) => 
        MDDR_DQ(14), MDDR_DQ(13) => MDDR_DQ(13), MDDR_DQ(12) => 
        MDDR_DQ(12), MDDR_DQ(11) => MDDR_DQ(11), MDDR_DQ(10) => 
        MDDR_DQ(10), MDDR_DQ(9) => MDDR_DQ(9), MDDR_DQ(8) => 
        MDDR_DQ(8), MDDR_DQ(7) => MDDR_DQ(7), MDDR_DQ(6) => 
        MDDR_DQ(6), MDDR_DQ(5) => MDDR_DQ(5), MDDR_DQ(4) => 
        MDDR_DQ(4), MDDR_DQ(3) => MDDR_DQ(3), MDDR_DQ(2) => 
        MDDR_DQ(2), MDDR_DQ(1) => MDDR_DQ(1), MDDR_DQ(0) => 
        MDDR_DQ(0), MDDR_DM_RDQS(1) => MDDR_DM_RDQS(1), 
        MDDR_DM_RDQS(0) => MDDR_DM_RDQS(0), MDDR_BA(2) => 
        MDDR_BA(2), MDDR_BA(1) => MDDR_BA(1), MDDR_BA(0) => 
        MDDR_BA(0), MDDR_ADDR(15) => MDDR_ADDR(15), MDDR_ADDR(14)
         => MDDR_ADDR(14), MDDR_ADDR(13) => MDDR_ADDR(13), 
        MDDR_ADDR(12) => MDDR_ADDR(12), MDDR_ADDR(11) => 
        MDDR_ADDR(11), MDDR_ADDR(10) => MDDR_ADDR(10), 
        MDDR_ADDR(9) => MDDR_ADDR(9), MDDR_ADDR(8) => 
        MDDR_ADDR(8), MDDR_ADDR(7) => MDDR_ADDR(7), MDDR_ADDR(6)
         => MDDR_ADDR(6), MDDR_ADDR(5) => MDDR_ADDR(5), 
        MDDR_ADDR(4) => MDDR_ADDR(4), MDDR_ADDR(3) => 
        MDDR_ADDR(3), MDDR_ADDR(2) => MDDR_ADDR(2), MDDR_ADDR(1)
         => MDDR_ADDR(1), MDDR_ADDR(0) => MDDR_ADDR(0), 
        CoreAPB3_0_APBmslave0_PADDR(7) => 
        \CoreAPB3_0_APBmslave0_PADDR[7]\, 
        CoreAPB3_0_APBmslave0_PADDR(6) => 
        \CoreAPB3_0_APBmslave0_PADDR[6]\, 
        CoreAPB3_0_APBmslave0_PADDR(5) => 
        \CoreAPB3_0_APBmslave0_PADDR[5]\, 
        CoreAPB3_0_APBmslave0_PADDR(4) => 
        \CoreAPB3_0_APBmslave0_PADDR[4]\, 
        CoreAPB3_0_APBmslave0_PADDR(3) => 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, 
        CoreAPB3_0_APBmslave0_PADDR(1) => 
        \CoreAPB3_0_APBmslave0_PADDR[1]\, 
        CoreAPB3_0_APBmslave0_PADDR(0) => 
        \CoreAPB3_0_APBmslave0_PADDR[0]\, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(15) => 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[15]\, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(14) => 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[14]\, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(13) => 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[13]\, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR(12) => 
        \m2s010_som_sb_0_FIC_0_APB_MASTER_PADDR[12]\, 
        CoreAPB3_0_APBmslave0_PWDATA(7) => 
        \CoreAPB3_0_APBmslave0_PWDATA[7]\, 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        \CoreAPB3_0_APBmslave0_PWDATA[6]\, 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        \CoreAPB3_0_APBmslave0_PWDATA[5]\, 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        \CoreAPB3_0_APBmslave0_PWDATA[4]\, 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        \CoreAPB3_0_APBmslave0_PWDATA[3]\, 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        \CoreAPB3_0_APBmslave0_PWDATA[2]\, 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        \CoreAPB3_0_APBmslave0_PWDATA[1]\, 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        \CoreAPB3_0_APBmslave0_PWDATA[0]\, MAC_MII_TXD_c(3) => 
        \MAC_MII_TXD_c[3]\, MAC_MII_TXD_c(2) => 
        \MAC_MII_TXD_c[2]\, MAC_MII_TXD_c(1) => 
        \MAC_MII_TXD_c[1]\, MAC_MII_TXD_c(0) => 
        \MAC_MII_TXD_c[0]\, CoreAPB3_0_APBmslave0_PRDATA_m(7) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[7]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(6) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[6]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(5) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[5]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(4) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[4]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(3) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[3]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(2) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[2]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(1) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[1]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(0) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[0]\, Y_net_0(3) => 
        \Y_net_0[3]\, Y_net_0(2) => \Y_net_0[2]\, Y_net_0(1) => 
        \Y_net_0[1]\, Y_net_0(0) => \Y_net_0[0]\, 
        MAC_MII_RXD_c(3) => \MAC_MII_RXD_c[3]\, MAC_MII_RXD_c(2)
         => \MAC_MII_RXD_c[2]\, MAC_MII_RXD_c(1) => 
        \MAC_MII_RXD_c[1]\, MAC_MII_RXD_c(0) => 
        \MAC_MII_RXD_c[0]\, SPI_1_SS0_OTH_0 => SPI_1_SS0_OTH(0), 
        DEBOUNCE_OUT_net_0_0 => \DEBOUNCE_OUT_net_0[0]\, 
        GPIO_7_PADI_0 => GPIO_7_PADI(0), GPIO_6_PAD_0 => 
        GPIO_6_PAD(0), GPIO_1_BI_0 => GPIO_1_BI(0), 
        SPI_1_SS0_CAM_0 => SPI_1_SS0_CAM(0), SPI_1_CLK_0 => 
        SPI_1_CLK(0), SPI_0_SS1 => SPI_0_SS1, SPI_0_SS0 => 
        SPI_0_SS0, SPI_0_DO => SPI_0_DO, SPI_0_DI => SPI_0_DI, 
        SPI_0_CLK => SPI_0_CLK, MMUART_1_TXD => MMUART_1_TXD, 
        MMUART_1_RXD => MMUART_1_RXD, MDDR_WE_N => MDDR_WE_N, 
        MDDR_RESET_N => MDDR_RESET_N, MDDR_RAS_N => MDDR_RAS_N, 
        MDDR_ODT => MDDR_ODT, MDDR_DQS_TMATCH_0_OUT => 
        MDDR_DQS_TMATCH_0_OUT, MDDR_DQS_TMATCH_0_IN => 
        MDDR_DQS_TMATCH_0_IN, MDDR_CS_N => MDDR_CS_N, MDDR_CKE
         => MDDR_CKE, MDDR_CAS_N => MDDR_CAS_N, I2C_1_SDA => 
        I2C_1_SDA, I2C_1_SCL => I2C_1_SCL, GPIO_31_BI => 
        GPIO_31_BI, GPIO_26_BI => GPIO_26_BI, GPIO_25_BI => 
        GPIO_25_BI, GPIO_20_OUT => GPIO_20_OUT, GPIO_18_BI => 
        GPIO_18_BI, GPIO_17_BI => GPIO_17_BI, GPIO_16_BI => 
        GPIO_16_BI, GPIO_15_BI => GPIO_15_BI, GPIO_14_BI => 
        GPIO_14_BI, GPIO_12_BI => GPIO_12_BI, GPIO_4_BI => 
        GPIO_4_BI, GPIO_3_BI => GPIO_3_BI, GPIO_0_BI => GPIO_0_BI, 
        CoreAPB3_0_APBmslave0_PENABLE => 
        CoreAPB3_0_APBmslave0_PENABLE, 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx => 
        m2s010_som_sb_0_FIC_0_APB_MASTER_PSELx, 
        CoreAPB3_0_APBmslave0_PWRITE => 
        CoreAPB3_0_APBmslave0_PWRITE, MAC_MII_MDC_c => 
        MAC_MII_MDC_c, GPIO_22_M2F_c => GPIO_22_M2F_c, 
        GPIO_21_M2F_c => GPIO_21_M2F_c, 
        m2s010_som_sb_0_GPIO_28_SW_RESET => 
        m2s010_som_sb_0_GPIO_28_SW_RESET, MMUART_0_TXD_M2F_c => 
        MMUART_0_TXD_M2F_c, GPIO_24_M2F_c => GPIO_24_M2F_c, 
        GPIO_5_M2F_c => GPIO_5_M2F_c, GPIO_8_M2F_c => 
        GPIO_8_M2F_c, GPIO_11_M2F_c => GPIO_11_M2F_c, 
        MAC_MII_TX_EN_c => MAC_MII_TX_EN_c, MAC_MII_COL_c => 
        MAC_MII_COL_c, MAC_MII_CRS_c => MAC_MII_CRS_c, 
        CommsFPGA_top_0_INT => CommsFPGA_top_0_INT, 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i => 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i, DEBOUNCE_OUT_1_c => 
        DEBOUNCE_OUT_1_c, DEBOUNCE_OUT_2_c => DEBOUNCE_OUT_2_c, 
        MMUART_0_RXD_F2M_c => MMUART_0_RXD_F2M_c, 
        MAC_MII_RX_CLK_c => MAC_MII_RX_CLK_c, MAC_MII_RX_DV_c => 
        MAC_MII_RX_DV_c, MAC_MII_RX_ER_c => MAC_MII_RX_ER_c, 
        MAC_MII_TX_CLK_c => MAC_MII_TX_CLK_c, MDDR_CLK_N => 
        MDDR_CLK_N, MDDR_CLK => MDDR_CLK, XTL => XTL, 
        m2s010_som_sb_0_CCC_71MHz => m2s010_som_sb_0_CCC_71MHz, 
        m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC => 
        m2s010_som_sb_0_XTLOSC_CCC_OUT_XTLOSC_CCC, SPI_1_DI_CAM_c
         => SPI_1_DI_CAM_c, SPI_1_DI_OTH_c => SPI_1_DI_OTH_c, 
        CommsFPGA_top_0_CAMERA_NODE => 
        CommsFPGA_top_0_CAMERA_NODE, DEVRST_N => DEVRST_N, 
        m2s010_som_sb_0_POWER_ON_RESET_N => 
        m2s010_som_sb_0_POWER_ON_RESET_N, MAC_MII_MDIO => 
        MAC_MII_MDIO, SPI_1_DO_CAM_c => SPI_1_DO_CAM_c, 
        SPI_1_DO_OTH => SPI_1_DO_OTH);
    
    GPIO_24_M2F_obuf : OUTBUF
      port map(D => GPIO_24_M2F_c, PAD => GPIO_24_M2F);
    
    \DEBOUNCE_IN_ibuf[2]\ : INBUF
      port map(PAD => DEBOUNCE_IN(2), Y => \DEBOUNCE_IN_c[2]\);
    
    \MAC_MII_RXD_ibuf[2]\ : INBUF
      port map(PAD => MAC_MII_RXD(2), Y => \MAC_MII_RXD_c[2]\);
    
    PULLDOWN_R9_ibuf : INBUF
      port map(PAD => PULLDOWN_R9, Y => Data_FAIL_c);
    
    GPIO_11_M2F_obuf : OUTBUF
      port map(D => GPIO_11_M2F_c, PAD => GPIO_11_M2F);
    
    GPIO_8_M2F_obuf : OUTBUF
      port map(D => GPIO_8_M2F_c, PAD => GPIO_8_M2F);
    
    \MAC_MII_TXD_obuf[2]\ : OUTBUF
      port map(D => \MAC_MII_TXD_c[2]\, PAD => MAC_MII_TXD(2));
    
    MAC_MII_RX_ER_ibuf : INBUF
      port map(PAD => MAC_MII_RX_ER, Y => MAC_MII_RX_ER_c);
    
    \DEBOUNCE_IN_ibuf[0]\ : INBUF
      port map(PAD => DEBOUNCE_IN(0), Y => \DEBOUNCE_IN_c[0]\);
    
    GPIO_5_M2F_obuf : OUTBUF
      port map(D => GPIO_5_M2F_c, PAD => GPIO_5_M2F);
    
    CommsFPGA_top_0 : CommsFPGA_top
      port map(packet_available_clear_reg(2) => 
        \packet_available_clear_reg[2]\, 
        packet_available_clear_reg(1) => 
        \packet_available_clear_reg[1]\, 
        packet_available_clear_reg(0) => 
        \packet_available_clear_reg[0]\, ReadFIFO_Read_Ptr(1) => 
        \ReadFIFO_Read_Ptr[1]\, ReadFIFO_Read_Ptr(0) => 
        \ReadFIFO_Read_Ptr[0]\, ReadFIFO_Write_Ptr(1) => 
        \ReadFIFO_Write_Ptr[1]\, ReadFIFO_Write_Ptr(0) => 
        \ReadFIFO_Write_Ptr[0]\, iRX_FIFO_Empty(3) => 
        \iRX_FIFO_Empty[3]\, iRX_FIFO_Empty(2) => 
        \iRX_FIFO_Empty[2]\, iRX_FIFO_Empty(1) => 
        \iRX_FIFO_Empty[1]\, iRX_FIFO_Empty(0) => 
        \iRX_FIFO_Empty[0]\, iRX_FIFO_UNDERRUN(3) => 
        \iRX_FIFO_UNDERRUN[3]\, iRX_FIFO_UNDERRUN(2) => 
        \iRX_FIFO_UNDERRUN[2]\, iRX_FIFO_UNDERRUN(1) => 
        \iRX_FIFO_UNDERRUN[1]\, iRX_FIFO_UNDERRUN(0) => 
        \iRX_FIFO_UNDERRUN[0]\, iRX_FIFO_Full(3) => 
        \iRX_FIFO_Full[3]\, iRX_FIFO_Full(2) => 
        \iRX_FIFO_Full[2]\, iRX_FIFO_Full(1) => 
        \iRX_FIFO_Full[1]\, iRX_FIFO_Full(0) => 
        \iRX_FIFO_Full[0]\, CoreAPB3_0_APBmslave0_PRDATA_m(7) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[7]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(6) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[6]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(5) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[5]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(4) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[4]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(3) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[3]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(2) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[2]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(1) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[1]\, 
        CoreAPB3_0_APBmslave0_PRDATA_m(0) => 
        \CoreAPB3_0_APBmslave0_PRDATA_m[0]\, un15(10) => 
        \un15[10]\, un15(9) => \un15[9]\, un15(8) => \un15[8]\, 
        un15(7) => \un15[7]\, un15(6) => nc3, un15(5) => 
        \un15[5]\, un15(4) => \un15[4]\, un15(3) => \un15[3]\, 
        un15(2) => \un15[2]\, un15(1) => \un15[1]\, un15(0) => 
        \un15[0]\, RX_FIFO_DIN(7) => \RX_FIFO_DIN[7]\, 
        RX_FIFO_DIN(6) => \RX_FIFO_DIN[6]\, RX_FIFO_DIN(5) => 
        \RX_FIFO_DIN[5]\, RX_FIFO_DIN(4) => \RX_FIFO_DIN[4]\, 
        RX_FIFO_DIN(3) => \RX_FIFO_DIN[3]\, RX_FIFO_DIN(2) => 
        \RX_FIFO_DIN[2]\, RX_FIFO_DIN(1) => \RX_FIFO_DIN[1]\, 
        RX_FIFO_DIN(0) => \RX_FIFO_DIN[0]\, RX_FIFO_DIN_pipe(8)
         => \RX_FIFO_DIN_pipe[8]\, RX_FIFO_DIN_pipe(7) => 
        \RX_FIFO_DIN_pipe[7]\, RX_FIFO_DIN_pipe(6) => 
        \RX_FIFO_DIN_pipe[6]\, RX_FIFO_DIN_pipe(5) => 
        \RX_FIFO_DIN_pipe[5]\, RX_FIFO_DIN_pipe(4) => 
        \RX_FIFO_DIN_pipe[4]\, RX_FIFO_DIN_pipe(3) => 
        \RX_FIFO_DIN_pipe[3]\, RX_FIFO_DIN_pipe(2) => 
        \RX_FIFO_DIN_pipe[2]\, RX_FIFO_DIN_pipe(1) => 
        \RX_FIFO_DIN_pipe[1]\, RX_FIFO_DIN_pipe(0) => 
        \RX_FIFO_DIN_pipe[0]\, clkdiv(3) => \clkdiv[3]\, 
        clkdiv(2) => \clkdiv[2]\, clkdiv(1) => \clkdiv[1]\, 
        clkdiv(0) => \clkdiv[0]\, un6(5) => \un6[5]\, un6(4) => 
        \un6[4]\, un6(3) => \un6[3]\, un6(2) => \un6[2]\, un6(1)
         => nc1, un6(0) => \un6[0]\, p2s_data(7) => \p2s_data[7]\, 
        p2s_data(6) => \p2s_data[6]\, p2s_data(5) => 
        \p2s_data[5]\, p2s_data(4) => \p2s_data[4]\, p2s_data(3)
         => \p2s_data[3]\, p2s_data(2) => \p2s_data[2]\, 
        p2s_data(1) => \p2s_data[1]\, p2s_data(0) => 
        \p2s_data[0]\, manches_in_dly(1) => \manches_in_dly[1]\, 
        manches_in_dly(0) => \manches_in_dly[0]\, 
        CoreAPB3_0_APBmslave0_PWDATA(7) => 
        \CoreAPB3_0_APBmslave0_PWDATA[7]\, 
        CoreAPB3_0_APBmslave0_PWDATA(6) => 
        \CoreAPB3_0_APBmslave0_PWDATA[6]\, 
        CoreAPB3_0_APBmslave0_PWDATA(5) => 
        \CoreAPB3_0_APBmslave0_PWDATA[5]\, 
        CoreAPB3_0_APBmslave0_PWDATA(4) => 
        \CoreAPB3_0_APBmslave0_PWDATA[4]\, 
        CoreAPB3_0_APBmslave0_PWDATA(3) => 
        \CoreAPB3_0_APBmslave0_PWDATA[3]\, 
        CoreAPB3_0_APBmslave0_PWDATA(2) => 
        \CoreAPB3_0_APBmslave0_PWDATA[2]\, 
        CoreAPB3_0_APBmslave0_PWDATA(1) => 
        \CoreAPB3_0_APBmslave0_PWDATA[1]\, 
        CoreAPB3_0_APBmslave0_PWDATA(0) => 
        \CoreAPB3_0_APBmslave0_PWDATA[0]\, 
        CoreAPB3_0_APBmslave0_PRDATA(7) => 
        \CoreAPB3_0_APBmslave0_PRDATA[7]\, 
        CoreAPB3_0_APBmslave0_PRDATA(6) => 
        \CoreAPB3_0_APBmslave0_PRDATA[6]\, 
        CoreAPB3_0_APBmslave0_PRDATA(5) => 
        \CoreAPB3_0_APBmslave0_PRDATA[5]\, 
        CoreAPB3_0_APBmslave0_PRDATA(4) => 
        \CoreAPB3_0_APBmslave0_PRDATA[4]\, 
        CoreAPB3_0_APBmslave0_PRDATA(3) => 
        \CoreAPB3_0_APBmslave0_PRDATA[3]\, 
        CoreAPB3_0_APBmslave0_PRDATA(2) => 
        \CoreAPB3_0_APBmslave0_PRDATA[2]\, 
        CoreAPB3_0_APBmslave0_PRDATA(1) => 
        \CoreAPB3_0_APBmslave0_PRDATA[1]\, 
        CoreAPB3_0_APBmslave0_PRDATA(0) => 
        \CoreAPB3_0_APBmslave0_PRDATA[0]\, RX_packet_depth(7) => 
        \RX_packet_depth[7]\, RX_packet_depth(6) => 
        \RX_packet_depth[6]\, RX_packet_depth(5) => 
        \RX_packet_depth[5]\, RX_packet_depth(4) => 
        \RX_packet_depth[4]\, RX_packet_depth(3) => 
        \RX_packet_depth[3]\, RX_packet_depth(2) => 
        \RX_packet_depth[2]\, RX_packet_depth(1) => 
        \RX_packet_depth[1]\, RX_packet_depth(0) => 
        \RX_packet_depth[0]\, CoreAPB3_0_APBmslave0_PADDR(7) => 
        \CoreAPB3_0_APBmslave0_PADDR[7]\, 
        CoreAPB3_0_APBmslave0_PADDR(6) => 
        \CoreAPB3_0_APBmslave0_PADDR[6]\, 
        CoreAPB3_0_APBmslave0_PADDR(5) => 
        \CoreAPB3_0_APBmslave0_PADDR[5]\, 
        CoreAPB3_0_APBmslave0_PADDR(4) => 
        \CoreAPB3_0_APBmslave0_PADDR[4]\, 
        CoreAPB3_0_APBmslave0_PADDR(3) => 
        \CoreAPB3_0_APBmslave0_PADDR[3]\, 
        CoreAPB3_0_APBmslave0_PADDR(2) => 
        \CoreAPB3_0_APBmslave0_PADDR[2]\, 
        CoreAPB3_0_APBmslave0_PADDR(1) => 
        \CoreAPB3_0_APBmslave0_PADDR[1]\, 
        CoreAPB3_0_APBmslave0_PADDR(0) => 
        \CoreAPB3_0_APBmslave0_PADDR[0]\, RX_FIFO_DOUT(8) => 
        \RX_FIFO_DOUT[8]\, RX_FIFO_DOUT(7) => \RX_FIFO_DOUT[7]\, 
        RX_FIFO_DOUT(6) => \RX_FIFO_DOUT[6]\, RX_FIFO_DOUT(5) => 
        \RX_FIFO_DOUT[5]\, RX_FIFO_DOUT(4) => \RX_FIFO_DOUT[4]\, 
        RX_FIFO_DOUT(3) => \RX_FIFO_DOUT[3]\, RX_FIFO_DOUT(2) => 
        \RX_FIFO_DOUT[2]\, RX_FIFO_DOUT(1) => \RX_FIFO_DOUT[1]\, 
        RX_FIFO_DOUT(0) => \RX_FIFO_DOUT[0]\, int_reg(7) => 
        \int_reg[7]\, int_reg(6) => \int_reg[6]\, int_reg(5) => 
        \int_reg[5]\, int_reg(4) => \int_reg[4]\, int_reg(3) => 
        \int_reg[3]\, int_reg(2) => \int_reg[2]\, int_reg(1) => 
        \int_reg[1]\, up_EOP_del(5) => \up_EOP_del[5]\, 
        up_EOP_del(4) => \up_EOP_del[4]\, up_EOP_del(3) => 
        \up_EOP_del[3]\, up_EOP_del(2) => \up_EOP_del[2]\, 
        up_EOP_del(1) => \up_EOP_del[1]\, up_EOP_del(0) => 
        \up_EOP_del[0]\, DEBOUNCE_IN_c(2) => \DEBOUNCE_IN_c[2]\, 
        DEBOUNCE_IN_c(1) => \DEBOUNCE_IN_c[1]\, DEBOUNCE_IN_c(0)
         => \DEBOUNCE_IN_c[0]\, Y_net_0(3) => \Y_net_0[3]\, 
        Y_net_0(2) => \Y_net_0[2]\, Y_net_0(1) => \Y_net_0[1]\, 
        control_reg_0 => \control_reg[0]\, control_reg_2 => 
        \control_reg[2]\, control_reg_3 => \control_reg[3]\, 
        DEBOUNCE_OUT_net_0_0 => \DEBOUNCE_OUT_net_0[0]\, 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i => 
        CoreAPB3_0_APBmslave0_PREADY_i_m_i, MANCHESTER_IN_c => 
        MANCHESTER_IN_c, irx_center_sample => irx_center_sample, 
        iNRZ_data => iNRZ_data, MANCH_OUT_P_c => MANCH_OUT_P_c, 
        MANCH_OUT_P_c_i => MANCH_OUT_P_c_i, DRVR_EN_c => 
        DRVR_EN_c, iup_EOP => iup_EOP, long_reset_set => 
        \long_reset_set\, CoreAPB3_0_APBmslave0_PREADY => 
        CoreAPB3_0_APBmslave0_PREADY, external_loopback => 
        external_loopback, internal_loopback => internal_loopback, 
        start_tx_FIFO => start_tx_FIFO, TX_FIFO_RST => 
        TX_FIFO_RST, N_480_i_i => \CommsFPGA_top_0.N_480_i_i\, 
        RX_FIFO_rd_en => RX_FIFO_rd_en, TX_FIFO_wr_en => 
        TX_FIFO_wr_en, RX_packet_depth_status => 
        RX_packet_depth_status, rx_packet_complt => 
        rx_packet_complt, rx_packet_avail_int => 
        rx_packet_avail_int, TX_FIFO_Full => TX_FIFO_Full, 
        TX_FIFO_Empty => TX_FIFO_Empty, 
        CoreAPB3_0_APBmslave0_PSELx => 
        CoreAPB3_0_APBmslave0_PSELx, 
        CoreAPB3_0_APBmslave0_PENABLE => 
        CoreAPB3_0_APBmslave0_PENABLE, RX_FIFO_Full => 
        RX_FIFO_Full, RX_FIFO_Empty => RX_FIFO_Empty, 
        CoreAPB3_0_APBmslave0_PWRITE => 
        CoreAPB3_0_APBmslave0_PWRITE, N_480_i => N_480_i, 
        CommsFPGA_top_0_INT => CommsFPGA_top_0_INT, int_reg_clr
         => int_reg_clr, rx_FIFO_UNDERRUN_int => 
        rx_FIFO_UNDERRUN_int, rx_FIFO_OVERFLOW_int => 
        rx_FIFO_OVERFLOW_int, rx_CRC_error_int => 
        rx_CRC_error_int, tx_packet_complt => tx_packet_complt, 
        block_int_until_rd => block_int_until_rd, RESET_set => 
        \RESET_set\, DEBOUNCE_OUT_1_c => DEBOUNCE_OUT_1_c, 
        DEBOUNCE_OUT_2_c => DEBOUNCE_OUT_2_c, 
        CommsFPGA_top_0_CAMERA_NODE => 
        CommsFPGA_top_0_CAMERA_NODE, CommsFPGA_CCC_0_LOCK => 
        CommsFPGA_CCC_0_LOCK, m2s010_som_sb_0_POWER_ON_RESET_N
         => m2s010_som_sb_0_POWER_ON_RESET_N, 
        m2s010_som_sb_0_GPIO_28_SW_RESET => 
        m2s010_som_sb_0_GPIO_28_SW_RESET, rx_FIFO_rst_reg => 
        rx_FIFO_rst_reg, CommsFPGA_CCC_0_GL1 => 
        CommsFPGA_CCC_0_GL1, CommsFPGA_CCC_0_GL0 => 
        CommsFPGA_CCC_0_GL0, m2s010_som_sb_0_CCC_71MHz => 
        m2s010_som_sb_0_CCC_71MHz, long_reset_i => long_reset_i, 
        RESET_i => RESET_i, RESET => RESET, BIT_CLK => 
        \CommsFPGA_top_0.BIT_CLK\, long_reset => long_reset, 
        bd_reset => bd_reset);
    

end DEF_ARCH; 
